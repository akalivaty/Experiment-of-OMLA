//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n829, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1031, new_n1032,
    new_n1033;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(KEYINPUT16), .A3(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT97), .ZN(new_n205));
  OAI221_X1 g004(.A(new_n204), .B1(new_n205), .B2(G8gat), .C1(new_n203), .C2(new_n202), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(G8gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT98), .ZN(new_n209));
  INV_X1    g008(.A(new_n207), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n206), .B(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT98), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n209), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G29gat), .ZN(new_n215));
  INV_X1    g014(.A(G36gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n217), .B(KEYINPUT14), .ZN(new_n218));
  NAND2_X1  g017(.A1(G29gat), .A2(G36gat), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT15), .ZN(new_n221));
  INV_X1    g020(.A(G50gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G43gat), .ZN(new_n223));
  INV_X1    g022(.A(G43gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G50gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n221), .B1(new_n226), .B2(KEYINPUT94), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(KEYINPUT94), .B2(new_n226), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n220), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT95), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n225), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(new_n223), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n225), .A2(new_n230), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n221), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  XOR2_X1   g033(.A(new_n219), .B(KEYINPUT96), .Z(new_n235));
  NAND4_X1  g034(.A1(new_n228), .A2(new_n218), .A3(new_n234), .A4(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n229), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n214), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n237), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT17), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT17), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n240), .A2(new_n211), .A3(new_n242), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G229gat), .A2(G233gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n244), .A2(KEYINPUT18), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT99), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n247), .B1(new_n214), .B2(new_n237), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n213), .A2(new_n209), .A3(KEYINPUT99), .A4(new_n239), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(new_n238), .A3(new_n249), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n245), .B(KEYINPUT13), .Z(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n238), .A2(new_n243), .A3(new_n245), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT18), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n246), .A2(new_n252), .A3(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G113gat), .B(G141gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(KEYINPUT11), .ZN(new_n258));
  INV_X1    g057(.A(G169gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(G197gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT12), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n256), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT100), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n246), .A2(new_n252), .A3(new_n262), .A4(new_n255), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n265), .B1(new_n264), .B2(new_n266), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G78gat), .B(G106gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT31), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(new_n222), .ZN(new_n272));
  INV_X1    g071(.A(G22gat), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT3), .ZN(new_n274));
  INV_X1    g073(.A(G162gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(G155gat), .ZN(new_n276));
  INV_X1    g075(.A(G155gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(G162gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G141gat), .B(G148gat), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n279), .B1(new_n280), .B2(KEYINPUT2), .ZN(new_n281));
  INV_X1    g080(.A(G148gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n282), .A2(G141gat), .ZN(new_n283));
  AND2_X1   g082(.A1(KEYINPUT82), .A2(G148gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(KEYINPUT82), .A2(G148gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n283), .B1(new_n286), .B2(G141gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(KEYINPUT83), .A2(G162gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT2), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n289), .A2(new_n276), .A3(new_n278), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n274), .B(new_n281), .C1(new_n287), .C2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT29), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G211gat), .B(G218gat), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT77), .ZN(new_n297));
  AND2_X1   g096(.A1(G197gat), .A2(G204gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(G197gat), .A2(G204gat), .ZN(new_n299));
  OAI22_X1  g098(.A1(new_n296), .A2(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AND2_X1   g099(.A1(new_n296), .A2(new_n297), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n295), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AND2_X1   g101(.A1(G211gat), .A2(G218gat), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT77), .B1(new_n303), .B2(KEYINPUT22), .ZN(new_n304));
  XNOR2_X1  g103(.A(G197gat), .B(G204gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n296), .A2(new_n297), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n304), .A2(new_n294), .A3(new_n305), .A4(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n281), .B1(new_n287), .B2(new_n290), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT29), .B1(new_n302), .B2(new_n307), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n311), .B1(new_n312), .B2(KEYINPUT3), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G228gat), .ZN(new_n315));
  INV_X1    g114(.A(G233gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT82), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(new_n282), .ZN(new_n320));
  NAND2_X1  g119(.A1(KEYINPUT82), .A2(G148gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(G141gat), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n283), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AND3_X1   g123(.A1(new_n289), .A2(new_n276), .A3(new_n278), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT2), .ZN(new_n326));
  INV_X1    g125(.A(G141gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n327), .A2(G148gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n283), .B2(new_n328), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n324), .A2(new_n325), .B1(new_n329), .B2(new_n279), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT29), .B1(new_n330), .B2(new_n274), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT87), .B1(new_n331), .B2(new_n308), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n314), .A2(new_n318), .A3(new_n332), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n310), .B(new_n313), .C1(KEYINPUT87), .C2(new_n317), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n273), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT88), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n272), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n308), .B1(new_n292), .B2(new_n291), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n308), .A2(new_n292), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n274), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n338), .B1(new_n340), .B2(new_n311), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT87), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n318), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n334), .ZN(new_n345));
  OAI21_X1  g144(.A(G22gat), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n333), .A2(new_n273), .A3(new_n334), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n337), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n346), .A2(new_n336), .A3(new_n347), .A4(new_n272), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT85), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT4), .ZN(new_n354));
  INV_X1    g153(.A(G113gat), .ZN(new_n355));
  INV_X1    g154(.A(G120gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT1), .ZN(new_n358));
  NAND2_X1  g157(.A1(G113gat), .A2(G120gat), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(G127gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(G134gat), .ZN(new_n362));
  INV_X1    g161(.A(G134gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(G127gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT72), .B1(new_n360), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G127gat), .B(G134gat), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT72), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT1), .B1(new_n355), .B2(new_n356), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n367), .A2(new_n368), .A3(new_n359), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n363), .A2(G127gat), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT71), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n369), .A2(new_n359), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n367), .A2(KEYINPUT71), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AND4_X1   g175(.A1(new_n354), .A2(new_n330), .A3(new_n371), .A4(new_n376), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n366), .A2(new_n370), .B1(new_n375), .B2(new_n374), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n354), .B1(new_n378), .B2(new_n330), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n353), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n330), .A2(new_n371), .A3(new_n376), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT4), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n378), .A2(new_n354), .A3(new_n330), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(KEYINPUT85), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(G225gat), .A2(G233gat), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  AOI22_X1  g185(.A1(KEYINPUT3), .A2(new_n311), .B1(new_n371), .B2(new_n376), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n386), .B1(new_n387), .B2(new_n291), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT5), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n380), .A2(new_n384), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT86), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI211_X1 g191(.A(KEYINPUT5), .B(new_n386), .C1(new_n387), .C2(new_n291), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n393), .A2(KEYINPUT86), .A3(new_n384), .A4(new_n380), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  AND3_X1   g194(.A1(new_n330), .A2(new_n371), .A3(new_n376), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n324), .A2(new_n325), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n371), .A2(new_n376), .B1(new_n397), .B2(new_n281), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n386), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT5), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n382), .A2(new_n383), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n388), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n400), .B1(KEYINPUT84), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT84), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n395), .A2(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G1gat), .B(G29gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(KEYINPUT0), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(G57gat), .ZN(new_n410));
  INV_X1    g209(.A(G85gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n407), .A2(KEYINPUT6), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n415));
  AOI22_X1  g214(.A1(new_n392), .A2(new_n394), .B1(new_n403), .B2(new_n405), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n415), .B1(new_n416), .B2(new_n412), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n395), .A2(new_n406), .A3(new_n412), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n414), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT25), .ZN(new_n421));
  NAND2_X1  g220(.A1(G169gat), .A2(G176gat), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT65), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(G176gat), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n259), .A2(new_n427), .A3(KEYINPUT23), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT66), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  AND3_X1   g228(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n428), .B(KEYINPUT66), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(G183gat), .A2(G190gat), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT67), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT24), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n437), .B1(new_n436), .B2(new_n435), .ZN(new_n438));
  INV_X1    g237(.A(G183gat), .ZN(new_n439));
  INV_X1    g238(.A(G190gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT23), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n259), .A2(new_n427), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n438), .A2(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n421), .B1(new_n434), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT24), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n435), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n450), .A2(new_n441), .A3(new_n442), .ZN(new_n451));
  OR2_X1    g250(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n452));
  NAND2_X1  g251(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n452), .A2(KEYINPUT23), .A3(new_n259), .A4(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT25), .B1(new_n446), .B2(new_n445), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n451), .A2(new_n454), .A3(new_n455), .A4(new_n426), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n446), .A2(KEYINPUT69), .A3(KEYINPUT26), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT69), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n457), .A2(new_n426), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT26), .ZN(new_n462));
  AND4_X1   g261(.A1(KEYINPUT70), .A2(new_n462), .A3(new_n259), .A4(new_n427), .ZN(new_n463));
  NOR2_X1   g262(.A1(G169gat), .A2(G176gat), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT70), .B1(new_n464), .B2(new_n462), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT27), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(G183gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n439), .A2(KEYINPUT27), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(new_n470), .A3(new_n440), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT28), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n468), .A2(KEYINPUT68), .A3(G183gat), .ZN(new_n473));
  NOR2_X1   g272(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n474));
  AND2_X1   g273(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n473), .B(new_n474), .C1(new_n475), .C2(new_n468), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n472), .A2(new_n435), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n456), .B1(new_n467), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n292), .B1(new_n448), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(G226gat), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n480), .A2(new_n316), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  AND4_X1   g282(.A1(new_n426), .A2(new_n451), .A3(new_n454), .A4(new_n455), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n472), .A2(new_n435), .A3(new_n476), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n424), .A2(new_n425), .B1(new_n458), .B2(new_n459), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n486), .B(new_n457), .C1(new_n465), .C2(new_n463), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n484), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n435), .A2(new_n436), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT67), .B1(G183gat), .B2(G190gat), .ZN(new_n490));
  NOR3_X1   g289(.A1(new_n489), .A2(new_n490), .A3(KEYINPUT24), .ZN(new_n491));
  OAI22_X1  g290(.A1(new_n491), .A2(new_n443), .B1(KEYINPUT23), .B2(new_n464), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n428), .B1(new_n430), .B2(new_n431), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT66), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n432), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT25), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n482), .B1(new_n488), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n308), .A3(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G8gat), .B(G36gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(G92gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(KEYINPUT79), .B(G64gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT29), .B1(new_n488), .B2(new_n497), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT78), .B1(new_n505), .B2(new_n481), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT78), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n479), .A2(new_n507), .A3(new_n482), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n498), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n500), .B(new_n504), .C1(new_n509), .C2(new_n308), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT30), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT81), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n510), .A2(KEYINPUT81), .A3(new_n511), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n420), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n504), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n518), .A2(new_n511), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n500), .B(new_n519), .C1(new_n509), .C2(new_n308), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n483), .A2(new_n308), .A3(new_n499), .ZN(new_n521));
  NOR3_X1   g320(.A1(new_n505), .A2(KEYINPUT78), .A3(new_n481), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n507), .B1(new_n479), .B2(new_n482), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n499), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n521), .B1(new_n524), .B2(new_n309), .ZN(new_n525));
  OAI211_X1 g324(.A(KEYINPUT80), .B(new_n520), .C1(new_n525), .C2(new_n504), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n500), .B1(new_n509), .B2(new_n308), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(new_n518), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT80), .B1(new_n529), .B2(new_n520), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n352), .B1(new_n517), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT36), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n378), .B1(new_n448), .B2(new_n478), .ZN(new_n534));
  INV_X1    g333(.A(new_n378), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n488), .A2(new_n535), .A3(new_n497), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(G227gat), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n538), .A2(new_n316), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT34), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT34), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n537), .A2(new_n543), .A3(new_n540), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(G15gat), .B(G43gat), .Z(new_n547));
  XNOR2_X1  g346(.A(G71gat), .B(G99gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n534), .A2(new_n539), .A3(new_n536), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT33), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(KEYINPUT32), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT75), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n554), .A2(KEYINPUT75), .A3(new_n555), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n551), .A2(new_n553), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n552), .A2(new_n561), .A3(KEYINPUT32), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT76), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n552), .A2(new_n561), .A3(KEYINPUT76), .A4(KEYINPUT32), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n546), .B1(new_n560), .B2(new_n566), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n554), .A2(KEYINPUT75), .A3(new_n555), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT75), .B1(new_n554), .B2(new_n555), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n546), .B(new_n566), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n533), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(new_n545), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n574), .A2(KEYINPUT36), .A3(new_n570), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n532), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT89), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n520), .B1(new_n525), .B2(new_n504), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT80), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(new_n526), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n582), .A2(new_n420), .A3(new_n516), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n583), .A2(new_n352), .B1(new_n572), .B2(new_n575), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT89), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT38), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT37), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n504), .B1(new_n525), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n528), .A2(KEYINPUT37), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n587), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n518), .B1(new_n528), .B2(KEYINPUT37), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n509), .A2(new_n309), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n483), .A2(new_n309), .A3(new_n499), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT37), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n587), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n510), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n591), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n420), .A2(KEYINPUT91), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT91), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n414), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n311), .A2(KEYINPUT3), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n535), .A2(new_n603), .A3(new_n291), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n380), .A2(new_n384), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT39), .ZN(new_n606));
  AND3_X1   g405(.A1(new_n605), .A2(new_n606), .A3(new_n386), .ZN(new_n607));
  INV_X1    g406(.A(new_n398), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n608), .A2(new_n381), .A3(new_n385), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT39), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n610), .B1(new_n605), .B2(new_n386), .ZN(new_n611));
  NOR3_X1   g410(.A1(new_n607), .A2(new_n611), .A3(new_n413), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT90), .ZN(new_n613));
  OAI21_X1  g412(.A(KEYINPUT40), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n407), .A2(new_n413), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT40), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n605), .A2(new_n386), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n412), .B1(new_n617), .B2(new_n610), .ZN(new_n618));
  OAI211_X1 g417(.A(KEYINPUT90), .B(new_n616), .C1(new_n618), .C2(new_n607), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n614), .A2(new_n615), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n515), .ZN(new_n621));
  AOI21_X1  g420(.A(KEYINPUT81), .B1(new_n510), .B2(new_n511), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n529), .B(new_n520), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n352), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n602), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n578), .A2(new_n586), .A3(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n601), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n627), .B1(KEYINPUT91), .B2(new_n420), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT92), .B(KEYINPUT35), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n623), .A2(new_n630), .ZN(new_n631));
  AND3_X1   g430(.A1(new_n574), .A2(new_n351), .A3(new_n570), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n629), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n574), .A2(new_n351), .A3(new_n570), .ZN(new_n634));
  OAI211_X1 g433(.A(KEYINPUT93), .B(KEYINPUT35), .C1(new_n583), .C2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n615), .A2(new_n415), .A3(new_n418), .ZN(new_n637));
  AOI22_X1  g436(.A1(new_n637), .A2(new_n414), .B1(new_n514), .B2(new_n515), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n632), .A2(new_n638), .A3(new_n582), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT93), .B1(new_n639), .B2(KEYINPUT35), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n633), .B1(new_n636), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n269), .B1(new_n626), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G120gat), .B(G148gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(G176gat), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n645), .B(G204gat), .Z(new_n646));
  NAND2_X1  g445(.A1(G85gat), .A2(G92gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT7), .ZN(new_n648));
  NAND2_X1  g447(.A1(G99gat), .A2(G106gat), .ZN(new_n649));
  INV_X1    g448(.A(G92gat), .ZN(new_n650));
  AOI22_X1  g449(.A1(KEYINPUT8), .A2(new_n649), .B1(new_n411), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G99gat), .B(G106gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(G64gat), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n655), .A2(G57gat), .ZN(new_n656));
  INV_X1    g455(.A(G57gat), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n657), .A2(G64gat), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n656), .B1(KEYINPUT101), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n659), .B1(KEYINPUT101), .B2(new_n658), .ZN(new_n660));
  NAND2_X1  g459(.A1(G71gat), .A2(G78gat), .ZN(new_n661));
  OR2_X1    g460(.A1(G71gat), .A2(G78gat), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT9), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(KEYINPUT9), .B1(new_n658), .B2(new_n656), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n666), .A2(new_n661), .A3(new_n662), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n654), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(G230gat), .A2(G233gat), .ZN(new_n670));
  OR3_X1    g469(.A1(new_n669), .A2(KEYINPUT104), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT104), .B1(new_n669), .B2(new_n670), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT10), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n654), .A2(KEYINPUT10), .A3(new_n667), .A4(new_n665), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n670), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n646), .B1(new_n673), .B2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT106), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n675), .A2(new_n683), .A3(new_n676), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n683), .B1(new_n675), .B2(new_n676), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n670), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT103), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI211_X1 g487(.A(KEYINPUT103), .B(new_n670), .C1(new_n684), .C2(new_n685), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n646), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n682), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  AOI211_X1 g492(.A(KEYINPUT105), .B(new_n691), .C1(new_n688), .C2(new_n689), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n681), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT21), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n209), .B(new_n213), .C1(new_n697), .C2(new_n668), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(G183gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n700));
  NAND2_X1  g499(.A1(G231gat), .A2(G233gat), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n700), .B(new_n701), .Z(new_n702));
  XNOR2_X1  g501(.A(new_n699), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n668), .A2(new_n697), .ZN(new_n704));
  XOR2_X1   g503(.A(G127gat), .B(G155gat), .Z(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(G211gat), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n703), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n703), .A2(new_n708), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n654), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n240), .A2(new_n242), .A3(new_n712), .ZN(new_n713));
  AND2_X1   g512(.A1(G232gat), .A2(G233gat), .ZN(new_n714));
  AOI22_X1  g513(.A1(new_n237), .A2(new_n654), .B1(KEYINPUT41), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(G134gat), .B(G162gat), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n716), .B(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n714), .A2(KEYINPUT41), .ZN(new_n720));
  XNOR2_X1  g519(.A(G190gat), .B(G218gat), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n719), .B(new_n722), .Z(new_n723));
  NAND3_X1  g522(.A1(new_n696), .A2(new_n711), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(KEYINPUT107), .B1(new_n643), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n726));
  INV_X1    g525(.A(new_n724), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n642), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n420), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g531(.A(KEYINPUT16), .B(G8gat), .Z(new_n733));
  NAND3_X1  g532(.A1(new_n729), .A2(new_n623), .A3(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT42), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n725), .A2(new_n728), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n579), .B1(new_n514), .B2(new_n515), .ZN(new_n738));
  OAI21_X1  g537(.A(G8gat), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n729), .A2(KEYINPUT42), .A3(new_n623), .A4(new_n733), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n736), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT108), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n736), .A2(new_n739), .A3(KEYINPUT108), .A4(new_n740), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(G1325gat));
  NOR2_X1   g544(.A1(new_n567), .A2(new_n571), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  OR3_X1    g546(.A1(new_n737), .A2(G15gat), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(G15gat), .B1(new_n737), .B2(new_n576), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(G1326gat));
  NAND2_X1  g549(.A1(new_n729), .A2(new_n352), .ZN(new_n751));
  XNOR2_X1  g550(.A(KEYINPUT43), .B(G22gat), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(G1327gat));
  NOR3_X1   g552(.A1(new_n711), .A2(new_n695), .A3(new_n723), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n642), .A2(new_n215), .A3(new_n730), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT45), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n626), .A2(new_n641), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n723), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n711), .B(KEYINPUT109), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n264), .A2(new_n266), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n761), .A2(new_n763), .A3(new_n695), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n614), .A2(new_n619), .A3(new_n615), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n351), .B1(new_n738), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n766), .B1(new_n628), .B2(new_n598), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT110), .B1(new_n767), .B2(new_n577), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT110), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n625), .A2(new_n584), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n723), .B1(new_n771), .B2(new_n641), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n760), .B(new_n764), .C1(new_n772), .C2(KEYINPUT44), .ZN(new_n773));
  OAI21_X1  g572(.A(G29gat), .B1(new_n773), .B2(new_n420), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n756), .A2(new_n774), .ZN(G1328gat));
  NAND4_X1  g574(.A1(new_n642), .A2(new_n216), .A3(new_n623), .A4(new_n754), .ZN(new_n776));
  XOR2_X1   g575(.A(new_n776), .B(KEYINPUT46), .Z(new_n777));
  OAI21_X1  g576(.A(KEYINPUT111), .B1(new_n773), .B2(new_n738), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(G36gat), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n773), .A2(KEYINPUT111), .A3(new_n738), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n777), .B1(new_n779), .B2(new_n780), .ZN(G1329gat));
  OAI21_X1  g580(.A(G43gat), .B1(new_n773), .B2(new_n576), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT47), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n754), .A2(new_n224), .A3(new_n746), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n782), .B1(new_n643), .B2(new_n785), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n784), .B(new_n786), .ZN(G1330gat));
  NOR2_X1   g586(.A1(new_n222), .A2(KEYINPUT113), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n788), .B1(new_n773), .B2(new_n351), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n351), .A2(KEYINPUT113), .A3(G50gat), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n642), .A2(new_n754), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  XOR2_X1   g591(.A(new_n792), .B(KEYINPUT48), .Z(G1331gat));
  AOI21_X1  g592(.A(new_n769), .B1(new_n625), .B2(new_n584), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n625), .A2(new_n584), .A3(new_n769), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n641), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n711), .A2(new_n695), .A3(new_n763), .A4(new_n723), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n730), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(G57gat), .ZN(G1332gat));
  INV_X1    g600(.A(new_n799), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n799), .A2(KEYINPUT114), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n738), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT115), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n799), .B(new_n803), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n809), .A2(new_n810), .A3(new_n806), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(KEYINPUT116), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n808), .A2(new_n811), .A3(new_n814), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(G1333gat));
  INV_X1    g617(.A(G71gat), .ZN(new_n819));
  INV_X1    g618(.A(new_n576), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n809), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n802), .A2(G71gat), .A3(new_n747), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n822), .A2(KEYINPUT50), .A3(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT50), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n826), .B1(new_n821), .B2(new_n823), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(G1334gat));
  NAND2_X1  g627(.A1(new_n809), .A2(new_n352), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g629(.A1(new_n696), .A2(new_n762), .A3(new_n711), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n760), .B(new_n831), .C1(new_n772), .C2(KEYINPUT44), .ZN(new_n832));
  OAI21_X1  g631(.A(G85gat), .B1(new_n832), .B2(new_n420), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n711), .A2(new_n762), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT51), .B1(new_n772), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n723), .ZN(new_n836));
  AND4_X1   g635(.A1(KEYINPUT51), .A2(new_n796), .A3(new_n836), .A4(new_n834), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n695), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n730), .A2(new_n411), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n833), .B1(new_n839), .B2(new_n840), .ZN(G1336gat));
  NOR2_X1   g640(.A1(new_n738), .A2(G92gat), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n838), .A2(new_n695), .A3(new_n842), .ZN(new_n843));
  OAI211_X1 g642(.A(KEYINPUT52), .B(G92gat), .C1(new_n832), .C2(new_n738), .ZN(new_n844));
  OR2_X1    g643(.A1(KEYINPUT117), .A2(KEYINPUT52), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(KEYINPUT118), .B1(new_n832), .B2(new_n738), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(G92gat), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n832), .A2(KEYINPUT118), .A3(new_n738), .ZN(new_n849));
  OAI22_X1  g648(.A1(new_n843), .A2(KEYINPUT117), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n846), .B1(new_n850), .B2(new_n851), .ZN(G1337gat));
  INV_X1    g651(.A(G99gat), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n832), .A2(new_n853), .A3(new_n576), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n838), .A2(new_n746), .A3(new_n695), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n854), .B1(new_n855), .B2(new_n853), .ZN(G1338gat));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n351), .A2(G106gat), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n695), .B(new_n858), .C1(new_n835), .C2(new_n837), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n860));
  OAI21_X1  g659(.A(G106gat), .B1(new_n832), .B2(new_n351), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n860), .B1(new_n859), .B2(new_n861), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n857), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n859), .A2(new_n861), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(KEYINPUT119), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(KEYINPUT53), .A3(new_n867), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n864), .A2(new_n868), .ZN(G1339gat));
  INV_X1    g668(.A(KEYINPUT109), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n711), .B(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n677), .A2(KEYINPUT102), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n675), .A2(new_n683), .A3(new_n676), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(KEYINPUT103), .B1(new_n874), .B2(new_n670), .ZN(new_n875));
  INV_X1    g674(.A(new_n689), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n692), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT105), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n690), .A2(new_n682), .A3(new_n692), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT54), .B1(new_n677), .B2(new_n670), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n882), .B1(new_n875), .B2(new_n876), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n678), .A2(KEYINPUT54), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(new_n646), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n883), .A2(KEYINPUT55), .A3(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT55), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n881), .B1(new_n688), .B2(new_n689), .ZN(new_n888));
  INV_X1    g687(.A(new_n885), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n880), .A2(new_n762), .A3(new_n886), .A4(new_n890), .ZN(new_n891));
  OAI22_X1  g690(.A1(new_n250), .A2(new_n251), .B1(new_n244), .B2(new_n245), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n261), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n266), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n695), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n836), .B1(new_n891), .B2(new_n896), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n886), .B(new_n890), .C1(new_n693), .C2(new_n694), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n898), .A2(new_n723), .A3(new_n894), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n871), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n724), .A2(new_n762), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n352), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n747), .A2(new_n420), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n903), .A2(new_n738), .A3(new_n904), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n905), .A2(new_n355), .A3(new_n269), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n903), .A2(new_n904), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n907), .A2(KEYINPUT120), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(KEYINPUT120), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n908), .A2(new_n738), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n762), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n906), .B1(new_n911), .B2(new_n355), .ZN(G1340gat));
  NOR2_X1   g711(.A1(new_n696), .A2(G120gat), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n908), .A2(new_n738), .A3(new_n909), .A4(new_n913), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n903), .A2(new_n738), .A3(new_n695), .A4(new_n904), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n915), .A2(KEYINPUT121), .A3(G120gat), .ZN(new_n916));
  AOI21_X1  g715(.A(KEYINPUT121), .B1(new_n915), .B2(G120gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n914), .B(KEYINPUT122), .C1(new_n916), .C2(new_n917), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1341gat));
  NAND3_X1  g721(.A1(new_n910), .A2(new_n361), .A3(new_n711), .ZN(new_n923));
  OAI21_X1  g722(.A(G127gat), .B1(new_n905), .B2(new_n871), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(G1342gat));
  NOR2_X1   g724(.A1(new_n723), .A2(G134gat), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n908), .A2(new_n738), .A3(new_n909), .A4(new_n926), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n927), .A2(KEYINPUT56), .ZN(new_n928));
  OAI21_X1  g727(.A(G134gat), .B1(new_n905), .B2(new_n723), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(KEYINPUT56), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(G1343gat));
  OAI21_X1  g730(.A(new_n896), .B1(new_n269), .B2(new_n898), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n723), .ZN(new_n933));
  INV_X1    g732(.A(new_n899), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n711), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n352), .B1(new_n935), .B2(new_n901), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(KEYINPUT57), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n820), .A2(new_n420), .A3(new_n623), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n351), .B1(new_n900), .B2(new_n902), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT57), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n269), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n937), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT124), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n937), .A2(new_n942), .A3(KEYINPUT124), .A4(new_n943), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n946), .A2(G141gat), .A3(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT58), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n940), .A2(new_n938), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n943), .A2(new_n327), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n948), .A2(new_n949), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n937), .A2(new_n942), .A3(new_n762), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(G141gat), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(new_n953), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT123), .B1(new_n957), .B2(KEYINPUT58), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n952), .B1(new_n955), .B2(G141gat), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT123), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n959), .A2(new_n960), .A3(new_n949), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n954), .B1(new_n958), .B2(new_n961), .ZN(G1344gat));
  INV_X1    g761(.A(new_n950), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n963), .A2(new_n286), .A3(new_n695), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n937), .A2(new_n942), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n965), .A2(new_n696), .ZN(new_n966));
  NOR3_X1   g765(.A1(new_n966), .A2(KEYINPUT59), .A3(new_n286), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT59), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n727), .A2(new_n269), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(KEYINPUT125), .ZN(new_n970));
  OAI211_X1 g769(.A(new_n941), .B(new_n352), .C1(new_n970), .C2(new_n935), .ZN(new_n971));
  OR2_X1    g770(.A1(new_n940), .A2(new_n941), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n971), .A2(new_n695), .A3(new_n938), .A4(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n968), .B1(new_n973), .B2(G148gat), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n964), .B1(new_n967), .B2(new_n974), .ZN(G1345gat));
  OAI21_X1  g774(.A(G155gat), .B1(new_n965), .B2(new_n871), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n963), .A2(new_n277), .A3(new_n711), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(G1346gat));
  XOR2_X1   g777(.A(KEYINPUT83), .B(G162gat), .Z(new_n979));
  NAND3_X1  g778(.A1(new_n963), .A2(new_n836), .A3(new_n979), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n965), .A2(new_n723), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n980), .B1(new_n981), .B2(new_n979), .ZN(G1347gat));
  NAND2_X1  g781(.A1(new_n623), .A2(new_n420), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n983), .A2(new_n747), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n903), .A2(new_n984), .ZN(new_n985));
  NOR3_X1   g784(.A1(new_n985), .A2(new_n259), .A3(new_n269), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n900), .A2(new_n902), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n987), .A2(new_n420), .ZN(new_n988));
  OR2_X1    g787(.A1(new_n988), .A2(KEYINPUT126), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n738), .B1(new_n988), .B2(KEYINPUT126), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n989), .A2(new_n632), .A3(new_n990), .ZN(new_n991));
  OR2_X1    g790(.A1(new_n991), .A2(new_n763), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n986), .B1(new_n992), .B2(new_n259), .ZN(G1348gat));
  OR2_X1    g792(.A1(new_n991), .A2(new_n696), .ZN(new_n994));
  INV_X1    g793(.A(new_n985), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n696), .B1(new_n452), .B2(new_n453), .ZN(new_n996));
  AOI22_X1  g795(.A1(new_n994), .A2(new_n427), .B1(new_n995), .B2(new_n996), .ZN(G1349gat));
  OAI21_X1  g796(.A(G183gat), .B1(new_n985), .B2(new_n871), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n711), .A2(new_n469), .A3(new_n470), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n998), .B1(new_n991), .B2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g799(.A(new_n1000), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g800(.A(G190gat), .B1(new_n985), .B2(new_n723), .ZN(new_n1002));
  AND2_X1   g801(.A1(new_n1002), .A2(KEYINPUT61), .ZN(new_n1003));
  NOR2_X1   g802(.A1(new_n1002), .A2(KEYINPUT61), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n836), .A2(new_n440), .ZN(new_n1005));
  OAI22_X1  g804(.A1(new_n1003), .A2(new_n1004), .B1(new_n991), .B2(new_n1005), .ZN(G1351gat));
  NOR2_X1   g805(.A1(new_n820), .A2(new_n351), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n989), .A2(new_n990), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT127), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g809(.A1(new_n989), .A2(new_n990), .A3(KEYINPUT127), .A4(new_n1007), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n1010), .A2(new_n762), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g811(.A(G197gat), .ZN(new_n1013));
  AND2_X1   g812(.A1(new_n971), .A2(new_n972), .ZN(new_n1014));
  NOR2_X1   g813(.A1(new_n820), .A2(new_n983), .ZN(new_n1015));
  AND2_X1   g814(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g815(.A1(new_n269), .A2(new_n1013), .ZN(new_n1017));
  AOI22_X1  g816(.A1(new_n1012), .A2(new_n1013), .B1(new_n1016), .B2(new_n1017), .ZN(G1352gat));
  NAND3_X1  g817(.A1(new_n1014), .A2(new_n695), .A3(new_n1015), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1019), .A2(G204gat), .ZN(new_n1020));
  OR2_X1    g819(.A1(new_n696), .A2(G204gat), .ZN(new_n1021));
  OAI21_X1  g820(.A(KEYINPUT62), .B1(new_n1008), .B2(new_n1021), .ZN(new_n1022));
  OR3_X1    g821(.A1(new_n1008), .A2(KEYINPUT62), .A3(new_n1021), .ZN(new_n1023));
  NAND3_X1  g822(.A1(new_n1020), .A2(new_n1022), .A3(new_n1023), .ZN(G1353gat));
  INV_X1    g823(.A(G211gat), .ZN(new_n1025));
  NAND4_X1  g824(.A1(new_n1010), .A2(new_n1025), .A3(new_n711), .A4(new_n1011), .ZN(new_n1026));
  NAND4_X1  g825(.A1(new_n971), .A2(new_n711), .A3(new_n972), .A4(new_n1015), .ZN(new_n1027));
  AND3_X1   g826(.A1(new_n1027), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1028));
  AOI21_X1  g827(.A(KEYINPUT63), .B1(new_n1027), .B2(G211gat), .ZN(new_n1029));
  OAI21_X1  g828(.A(new_n1026), .B1(new_n1028), .B2(new_n1029), .ZN(G1354gat));
  NAND3_X1  g829(.A1(new_n1010), .A2(new_n836), .A3(new_n1011), .ZN(new_n1031));
  INV_X1    g830(.A(G218gat), .ZN(new_n1032));
  NOR2_X1   g831(.A1(new_n723), .A2(new_n1032), .ZN(new_n1033));
  AOI22_X1  g832(.A1(new_n1031), .A2(new_n1032), .B1(new_n1016), .B2(new_n1033), .ZN(G1355gat));
endmodule


