//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n449, new_n452, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n567, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1163, new_n1164;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT67), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT68), .Z(G217));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT69), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(new_n455), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2106), .ZN(new_n461));
  INV_X1    g036(.A(new_n456), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G567), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n466), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT70), .B(G2105), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n467), .A2(G2105), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n473), .A2(new_n475), .B1(G101), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n474), .A2(G137), .ZN(new_n478));
  OR3_X1    g053(.A1(new_n478), .A2(KEYINPUT71), .A3(new_n471), .ZN(new_n479));
  OAI21_X1  g054(.A(KEYINPUT71), .B1(new_n478), .B2(new_n471), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n477), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  NOR2_X1   g057(.A1(new_n471), .A2(new_n474), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n471), .A2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  OAI221_X1 g061(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n474), .C2(G112), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n484), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  AND2_X1   g064(.A1(new_n468), .A2(new_n470), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n490), .A2(G126), .A3(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT72), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n493), .B(G2104), .C1(G114), .C2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT72), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n490), .A2(new_n496), .A3(G126), .A4(G2105), .ZN(new_n497));
  AND3_X1   g072(.A1(new_n492), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n499), .B1(KEYINPUT73), .B2(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n490), .A2(new_n474), .A3(new_n500), .ZN(new_n501));
  OR2_X1    g076(.A1(KEYINPUT73), .A2(KEYINPUT4), .ZN(new_n502));
  XNOR2_X1  g077(.A(new_n501), .B(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(G88), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT74), .B1(new_n509), .B2(G651), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT74), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n511), .A2(new_n507), .A3(KEYINPUT6), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n508), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n517), .B2(KEYINPUT5), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n514), .A2(KEYINPUT75), .A3(G543), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n513), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n513), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G50), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n506), .A2(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n520), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n507), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n524), .A2(new_n526), .ZN(G166));
  NAND3_X1  g102(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n528));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n522), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT76), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT76), .ZN(new_n532));
  OAI211_X1 g107(.A(new_n528), .B(new_n532), .C1(new_n522), .C2(new_n529), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n513), .A2(new_n520), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n531), .A2(new_n533), .B1(G89), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n535), .A2(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(new_n515), .ZN(new_n541));
  AND3_X1   g116(.A1(new_n514), .A2(KEYINPUT75), .A3(G543), .ZN(new_n542));
  AOI21_X1  g117(.A(KEYINPUT75), .B1(new_n514), .B2(G543), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G64), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n540), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G651), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n513), .A2(new_n520), .A3(G90), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n513), .A2(G52), .A3(G543), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT77), .ZN(new_n550));
  AND3_X1   g125(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n550), .B1(new_n548), .B2(new_n549), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n547), .B1(new_n551), .B2(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  NAND3_X1  g129(.A1(new_n513), .A2(new_n520), .A3(G81), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n510), .A2(new_n512), .ZN(new_n556));
  INV_X1    g131(.A(new_n508), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n556), .A2(G43), .A3(G543), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT78), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT78), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n555), .A2(new_n561), .A3(new_n558), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n564), .A2(new_n507), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(G860), .A3(new_n565), .ZN(G153));
  AND3_X1   g141(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G36), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n567), .A2(new_n570), .ZN(G188));
  AND2_X1   g146(.A1(new_n534), .A2(G91), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT80), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n544), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n520), .A2(KEYINPUT80), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n574), .A2(G65), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(G78), .A2(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n572), .B1(new_n578), .B2(G651), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n556), .A2(G53), .A3(G543), .A4(new_n557), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT79), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n513), .A2(new_n582), .A3(G53), .A4(G543), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(KEYINPUT9), .A3(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT9), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n580), .A2(KEYINPUT79), .A3(new_n585), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n579), .A2(new_n587), .ZN(G299));
  OR2_X1    g163(.A1(new_n524), .A2(new_n526), .ZN(G303));
  INV_X1    g164(.A(new_n522), .ZN(new_n590));
  AOI22_X1  g165(.A1(G49), .A2(new_n590), .B1(new_n534), .B2(G87), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n592), .A2(new_n593), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n591), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT82), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(G288));
  NAND2_X1  g173(.A1(new_n534), .A2(G86), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT83), .ZN(new_n600));
  NAND2_X1  g175(.A1(G73), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G61), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n544), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(new_n590), .B2(G48), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(G305));
  INV_X1    g180(.A(G85), .ZN(new_n606));
  INV_X1    g181(.A(G47), .ZN(new_n607));
  OAI22_X1  g182(.A1(new_n606), .A2(new_n521), .B1(new_n522), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n609), .A2(new_n507), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n608), .A2(new_n610), .ZN(G290));
  NAND2_X1  g186(.A1(G301), .A2(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n590), .A2(G54), .ZN(new_n613));
  AND3_X1   g188(.A1(new_n574), .A2(G66), .A3(new_n575), .ZN(new_n614));
  AND2_X1   g189(.A1(G79), .A2(G543), .ZN(new_n615));
  OAI21_X1  g190(.A(G651), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G92), .ZN(new_n617));
  OAI21_X1  g192(.A(KEYINPUT84), .B1(new_n521), .B2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n619));
  NAND4_X1  g194(.A1(new_n513), .A2(new_n520), .A3(new_n619), .A4(G92), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT10), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n618), .A2(KEYINPUT10), .A3(new_n620), .ZN(new_n624));
  AND4_X1   g199(.A1(new_n613), .A2(new_n616), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n612), .B1(new_n625), .B2(G868), .ZN(G284));
  OAI21_X1  g201(.A(new_n612), .B1(new_n625), .B2(G868), .ZN(G321));
  MUX2_X1   g202(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g203(.A(G299), .B(G286), .S(G868), .Z(G280));
  XNOR2_X1  g204(.A(KEYINPUT85), .B(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n625), .B1(G860), .B2(new_n630), .ZN(G148));
  AND3_X1   g206(.A1(new_n555), .A2(new_n561), .A3(new_n558), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n561), .B1(new_n555), .B2(new_n558), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n565), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n625), .A2(new_n630), .ZN(new_n635));
  MUX2_X1   g210(.A(new_n634), .B(new_n635), .S(G868), .Z(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g212(.A1(new_n490), .A2(new_n476), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT12), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2100), .ZN(new_n641));
  INV_X1    g216(.A(new_n485), .ZN(new_n642));
  INV_X1    g217(.A(G135), .ZN(new_n643));
  OR3_X1    g218(.A1(new_n642), .A2(KEYINPUT86), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n483), .A2(G123), .ZN(new_n645));
  OAI21_X1  g220(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n646));
  INV_X1    g221(.A(KEYINPUT87), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n648), .B(new_n649), .C1(G111), .C2(new_n474), .ZN(new_n650));
  OAI21_X1  g225(.A(KEYINPUT86), .B1(new_n642), .B2(new_n643), .ZN(new_n651));
  NAND4_X1  g226(.A1(new_n644), .A2(new_n645), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(G2096), .Z(new_n653));
  NAND2_X1  g228(.A1(new_n641), .A2(new_n653), .ZN(G156));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT88), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2438), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2427), .B(G2430), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(KEYINPUT14), .ZN(new_n660));
  XOR2_X1   g235(.A(G2451), .B(G2454), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n660), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1341), .B(G1348), .ZN(new_n664));
  AND2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2443), .B(G2446), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  OR3_X1    g243(.A1(new_n665), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n668), .B1(new_n665), .B2(new_n666), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n669), .A2(G14), .A3(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(G401));
  XOR2_X1   g247(.A(G2072), .B(G2078), .Z(new_n673));
  XOR2_X1   g248(.A(G2067), .B(G2678), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2084), .B(G2090), .Z(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n673), .B1(new_n677), .B2(KEYINPUT18), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G2096), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G2100), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n677), .A2(KEYINPUT17), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n675), .A2(new_n676), .ZN(new_n682));
  AOI21_X1  g257(.A(KEYINPUT18), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n680), .B(new_n683), .Z(G227));
  XNOR2_X1  g259(.A(G1971), .B(G1976), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT89), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT19), .Z(new_n687));
  XOR2_X1   g262(.A(G1956), .B(G2474), .Z(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  AND2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT20), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n688), .A2(new_n689), .ZN(new_n693));
  AOI22_X1  g268(.A1(new_n691), .A2(new_n692), .B1(new_n687), .B2(new_n693), .ZN(new_n694));
  OR3_X1    g269(.A1(new_n687), .A2(new_n690), .A3(new_n693), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n694), .B(new_n695), .C1(new_n692), .C2(new_n691), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT21), .B(G1986), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1991), .B(G1996), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT22), .B(G1981), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n700), .B(new_n701), .Z(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(G229));
  INV_X1    g278(.A(G25), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n704), .A2(G29), .ZN(new_n705));
  AOI22_X1  g280(.A1(G119), .A2(new_n483), .B1(new_n485), .B2(G131), .ZN(new_n706));
  OAI221_X1 g281(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n474), .C2(G107), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n705), .B1(new_n708), .B2(G29), .ZN(new_n709));
  MUX2_X1   g284(.A(new_n705), .B(new_n709), .S(KEYINPUT90), .Z(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT35), .B(G1991), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G24), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n608), .A2(new_n610), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n713), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G1986), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n716), .A2(G1986), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n712), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(G16), .A2(G23), .ZN(new_n720));
  INV_X1    g295(.A(new_n596), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(G16), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT33), .B(G1976), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n713), .A2(G22), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G166), .B2(new_n713), .ZN(new_n726));
  INV_X1    g301(.A(G1971), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n713), .A2(G6), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G305), .B2(G16), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT32), .B(G1981), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT34), .ZN(new_n734));
  OR3_X1    g309(.A1(new_n729), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n729), .B2(new_n733), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n719), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT91), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  AOI211_X1 g315(.A(KEYINPUT91), .B(new_n719), .C1(new_n735), .C2(new_n736), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n740), .A2(KEYINPUT92), .A3(KEYINPUT36), .A4(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT36), .ZN(new_n744));
  NOR3_X1   g319(.A1(new_n739), .A2(new_n741), .A3(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT92), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n737), .B2(new_n744), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n743), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  MUX2_X1   g323(.A(G19), .B(new_n634), .S(G16), .Z(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(G1341), .Z(new_n750));
  NOR2_X1   g325(.A1(G16), .A2(G21), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G168), .B2(G16), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n752), .A2(G1966), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT98), .Z(new_n754));
  INV_X1    g329(.A(G29), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n755), .A2(G35), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n488), .B2(G29), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT29), .ZN(new_n758));
  INV_X1    g333(.A(G2090), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT99), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT100), .B(KEYINPUT23), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n713), .A2(G20), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G299), .B2(G16), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G1956), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n761), .A2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT101), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n761), .A2(KEYINPUT101), .A3(new_n766), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n769), .A2(new_n770), .B1(G1966), .B2(new_n752), .ZN(new_n771));
  NOR2_X1   g346(.A1(G27), .A2(G29), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G164), .B2(G29), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G2078), .ZN(new_n774));
  INV_X1    g349(.A(G2084), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT24), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n755), .B1(new_n776), .B2(G34), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT95), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n776), .A2(G34), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n777), .A2(new_n778), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n481), .B2(new_n755), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n774), .B1(new_n775), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n713), .A2(G5), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G171), .B2(new_n713), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G1961), .ZN(new_n787));
  NOR2_X1   g362(.A1(G29), .A2(G33), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n490), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n789), .A2(new_n474), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT25), .ZN(new_n792));
  AOI211_X1 g367(.A(new_n790), .B(new_n792), .C1(G139), .C2(new_n485), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n788), .B1(new_n793), .B2(G29), .ZN(new_n794));
  AOI211_X1 g369(.A(new_n784), .B(new_n787), .C1(G2072), .C2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT30), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n796), .A2(G28), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(G28), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n797), .A2(new_n798), .A3(new_n755), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n652), .B2(new_n755), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n758), .B2(new_n759), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n713), .A2(G4), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n625), .B2(new_n713), .ZN(new_n803));
  INV_X1    g378(.A(G1348), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n771), .A2(new_n795), .A3(new_n801), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(G29), .A2(G32), .ZN(new_n807));
  AOI22_X1  g382(.A1(G129), .A2(new_n483), .B1(new_n485), .B2(G141), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n476), .A2(G105), .ZN(new_n809));
  NAND3_X1  g384(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT26), .Z(new_n811));
  NAND3_X1  g386(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT96), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n807), .B1(new_n813), .B2(G29), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT27), .B(G1996), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n783), .A2(new_n775), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT93), .B(KEYINPUT28), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT94), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n755), .A2(G26), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n820), .B(new_n821), .Z(new_n822));
  AOI22_X1  g397(.A1(G128), .A2(new_n483), .B1(new_n485), .B2(G140), .ZN(new_n823));
  OAI221_X1 g398(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n474), .C2(G116), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(G29), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G2067), .ZN(new_n828));
  XOR2_X1   g403(.A(KEYINPUT97), .B(KEYINPUT31), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(G11), .ZN(new_n830));
  OAI221_X1 g405(.A(new_n830), .B1(new_n773), .B2(G2078), .C1(new_n794), .C2(G2072), .ZN(new_n831));
  NOR4_X1   g406(.A1(new_n806), .A2(new_n818), .A3(new_n828), .A4(new_n831), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n748), .A2(new_n750), .A3(new_n754), .A4(new_n832), .ZN(G150));
  INV_X1    g408(.A(G150), .ZN(G311));
  NAND3_X1  g409(.A1(new_n513), .A2(G55), .A3(G543), .ZN(new_n835));
  INV_X1    g410(.A(G93), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n521), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n520), .A2(G67), .ZN(new_n838));
  NAND2_X1  g413(.A1(G80), .A2(G543), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n507), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(G860), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT37), .Z(new_n842));
  NAND2_X1  g417(.A1(new_n625), .A2(G559), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT38), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT39), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT102), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(new_n837), .B2(new_n840), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n838), .A2(new_n839), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G651), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n534), .A2(G93), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n849), .A2(KEYINPUT102), .A3(new_n850), .A4(new_n835), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n634), .A2(new_n847), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n837), .A2(new_n840), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n563), .A2(KEYINPUT102), .A3(new_n565), .A4(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n845), .B(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n842), .B1(new_n857), .B2(G860), .ZN(G145));
  XNOR2_X1  g433(.A(new_n481), .B(new_n488), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n652), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(new_n793), .Z(new_n861));
  XOR2_X1   g436(.A(new_n708), .B(new_n825), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n813), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT103), .ZN(new_n864));
  INV_X1    g439(.A(G142), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n864), .B1(new_n642), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n483), .A2(G130), .ZN(new_n867));
  OAI221_X1 g442(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n474), .C2(G118), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n485), .A2(KEYINPUT103), .A3(G142), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n866), .A2(new_n867), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n863), .B(new_n871), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n861), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n861), .A2(new_n872), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n504), .B(new_n639), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(G37), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n873), .A2(new_n876), .A3(new_n874), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g457(.A(KEYINPUT104), .ZN(new_n883));
  NAND2_X1  g458(.A1(G299), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n579), .A2(new_n587), .A3(KEYINPUT104), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n625), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT41), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n616), .A2(new_n623), .A3(new_n613), .A4(new_n624), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n888), .A2(G299), .A3(new_n883), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n892), .B1(new_n886), .B2(new_n889), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n635), .B(new_n856), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n886), .A2(new_n889), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n895), .A2(new_n900), .ZN(new_n901));
  OR3_X1    g476(.A1(new_n897), .A2(new_n898), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(G290), .A2(G166), .ZN(new_n903));
  NAND2_X1  g478(.A1(G303), .A2(new_n715), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n903), .A2(new_n904), .A3(new_n596), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n596), .B1(new_n903), .B2(new_n904), .ZN(new_n906));
  OR3_X1    g481(.A1(new_n905), .A2(new_n906), .A3(G305), .ZN(new_n907));
  OAI21_X1  g482(.A(G305), .B1(new_n905), .B2(new_n906), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n898), .B1(new_n897), .B2(new_n901), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n902), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n910), .B1(new_n902), .B2(new_n911), .ZN(new_n913));
  OAI21_X1  g488(.A(G868), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n914), .B1(G868), .B2(new_n853), .ZN(G295));
  OAI21_X1  g490(.A(new_n914), .B1(G868), .B2(new_n853), .ZN(G331));
  OAI211_X1 g491(.A(KEYINPUT107), .B(new_n547), .C1(new_n551), .C2(new_n552), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n852), .A2(new_n854), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n920));
  AOI22_X1  g495(.A1(new_n535), .A2(new_n537), .B1(G301), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n917), .B1(new_n852), .B2(new_n854), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n919), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n917), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n855), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n921), .B1(new_n926), .B2(new_n918), .ZN(new_n927));
  OAI22_X1  g502(.A1(new_n890), .A2(new_n893), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(new_n921), .A3(new_n918), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n922), .B1(new_n919), .B2(new_n923), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n900), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n909), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n879), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n579), .A2(KEYINPUT104), .A3(new_n587), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT104), .B1(new_n579), .B2(new_n587), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n934), .A2(new_n935), .A3(new_n888), .ZN(new_n936));
  INV_X1    g511(.A(new_n889), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n887), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n886), .A2(new_n889), .A3(new_n891), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n938), .B(new_n939), .C1(new_n924), .C2(new_n927), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n909), .B1(new_n940), .B2(new_n931), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT109), .B1(new_n933), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n931), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n910), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT109), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n944), .A2(new_n945), .A3(new_n879), .A4(new_n932), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n942), .A2(KEYINPUT43), .A3(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n891), .B1(new_n936), .B2(new_n937), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n948), .A2(new_n949), .B1(new_n930), .B2(new_n929), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n924), .A2(new_n927), .A3(new_n899), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n910), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n952), .A2(new_n879), .A3(new_n932), .ZN(new_n953));
  OR2_X1    g528(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n947), .A2(KEYINPUT44), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n944), .A2(new_n958), .A3(new_n879), .A4(new_n932), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n956), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AOI211_X1 g537(.A(KEYINPUT108), .B(KEYINPUT44), .C1(new_n957), .C2(new_n959), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n955), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT110), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n966), .B(new_n955), .C1(new_n962), .C2(new_n963), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(G397));
  INV_X1    g543(.A(G1384), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n504), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT45), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(G160), .A2(G40), .ZN(new_n973));
  OR3_X1    g548(.A1(new_n972), .A2(KEYINPUT111), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT111), .B1(new_n972), .B2(new_n973), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OR3_X1    g551(.A1(new_n976), .A2(KEYINPUT112), .A3(G1996), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT112), .B1(new_n976), .B2(G1996), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G2067), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n825), .B(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G1996), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n981), .B1(new_n813), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT113), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n976), .B(new_n984), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n979), .A2(new_n813), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n708), .A2(new_n711), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n708), .A2(new_n711), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n976), .ZN(new_n990));
  NOR2_X1   g565(.A1(G290), .A2(G1986), .ZN(new_n991));
  AND2_X1   g566(.A1(G290), .A2(G1986), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n986), .A2(new_n989), .A3(new_n993), .ZN(new_n994));
  XOR2_X1   g569(.A(new_n994), .B(KEYINPUT114), .Z(new_n995));
  INV_X1    g570(.A(G8), .ZN(new_n996));
  AND2_X1   g571(.A1(G160), .A2(G40), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n969), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n972), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G1966), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT50), .B1(new_n504), .B2(new_n969), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n1003));
  AOI211_X1 g578(.A(new_n1003), .B(G1384), .C1(new_n498), .C2(new_n503), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n775), .B(new_n997), .C1(new_n1002), .C2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n996), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(KEYINPUT116), .B(G8), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(G168), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(KEYINPUT51), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1008), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1009), .A2(KEYINPUT51), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT122), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT122), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n970), .A2(new_n1003), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n504), .A2(KEYINPUT50), .A3(new_n969), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n973), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n775), .A2(new_n1018), .B1(new_n999), .B2(new_n1000), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1015), .B(new_n1012), .C1(new_n1019), .C2(new_n1008), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1010), .A2(new_n1014), .A3(new_n1020), .ZN(new_n1021));
  OR3_X1    g596(.A1(new_n1019), .A2(G168), .A3(new_n1008), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT62), .ZN(new_n1024));
  XOR2_X1   g599(.A(KEYINPUT115), .B(G2090), .Z(new_n1025));
  AOI22_X1  g600(.A1(new_n1018), .A2(new_n1025), .B1(new_n999), .B2(new_n727), .ZN(new_n1026));
  NAND2_X1  g601(.A1(G303), .A2(G8), .ZN(new_n1027));
  XOR2_X1   g602(.A(new_n1027), .B(KEYINPUT55), .Z(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n1026), .A2(new_n1029), .A3(new_n996), .ZN(new_n1030));
  XOR2_X1   g605(.A(KEYINPUT117), .B(G1976), .Z(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT52), .B1(G288), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n970), .A2(new_n973), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1033), .A2(new_n1008), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n721), .A2(G1976), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1032), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT52), .ZN(new_n1038));
  INV_X1    g613(.A(G1981), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n600), .A2(new_n1039), .A3(new_n604), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT49), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n604), .A2(new_n599), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(G1981), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1041), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1034), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1036), .A2(new_n1038), .A3(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1030), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1029), .B1(new_n1026), .B2(new_n1008), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT62), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1021), .A2(new_n1052), .A3(new_n1022), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n972), .A2(new_n998), .ZN(new_n1054));
  INV_X1    g629(.A(G2078), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1054), .A2(KEYINPUT53), .A3(new_n1055), .A4(new_n997), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n997), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1057));
  INV_X1    g632(.A(G1961), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(new_n999), .B2(G2078), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1056), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1062), .A2(KEYINPUT123), .A3(G171), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT123), .B1(new_n1062), .B2(G171), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1024), .A2(new_n1051), .A3(new_n1053), .A4(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT124), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT124), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1068), .A2(new_n1069), .A3(new_n1065), .A4(new_n1024), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n1072));
  XNOR2_X1  g647(.A(G299), .B(new_n1072), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT56), .B(G2072), .Z(new_n1074));
  OAI221_X1 g649(.A(new_n1073), .B1(new_n999), .B2(new_n1074), .C1(G1956), .C2(new_n1018), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1057), .A2(new_n804), .B1(new_n980), .B2(new_n1033), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1076), .A2(new_n888), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  OAI22_X1  g653(.A1(new_n1018), .A2(G1956), .B1(new_n999), .B2(new_n1074), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1073), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n1075), .A2(KEYINPUT61), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n997), .A2(new_n504), .A3(new_n969), .ZN(new_n1083));
  OAI22_X1  g658(.A1(new_n1018), .A2(G1348), .B1(G2067), .B2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1084), .A2(new_n625), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT60), .B1(new_n1085), .B2(new_n1077), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n563), .A2(KEYINPUT120), .A3(new_n565), .ZN(new_n1087));
  XOR2_X1   g662(.A(KEYINPUT58), .B(G1341), .Z(new_n1088));
  NAND2_X1  g663(.A1(new_n1083), .A2(new_n1088), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT119), .B(G1996), .Z(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n972), .A2(new_n997), .A3(new_n998), .A4(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1087), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n1093), .B(new_n1094), .ZN(new_n1095));
  OR3_X1    g670(.A1(new_n1084), .A2(KEYINPUT60), .A3(new_n888), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1082), .A2(new_n1086), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1075), .A2(KEYINPUT121), .A3(KEYINPUT61), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT121), .B1(new_n1075), .B2(KEYINPUT61), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1078), .B(new_n1081), .C1(new_n1097), .C2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1056), .A2(G301), .A3(new_n1061), .A4(new_n1059), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1062), .A2(G171), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n1103), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT54), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1050), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1102), .A2(new_n1110), .A3(new_n1023), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1036), .A2(new_n1038), .A3(new_n1046), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n1030), .ZN(new_n1113));
  NOR4_X1   g688(.A1(new_n1044), .A2(new_n1045), .A3(G288), .A4(G1976), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1040), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1034), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1018), .A2(new_n1025), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n999), .A2(new_n727), .ZN(new_n1118));
  OAI211_X1 g693(.A(G8), .B(new_n1028), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1019), .A2(G286), .A3(new_n1008), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1112), .A2(new_n1119), .A3(new_n1120), .A4(new_n1049), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT63), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT118), .ZN(new_n1124));
  OAI21_X1  g699(.A(G8), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1122), .B1(new_n1125), .B2(new_n1029), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1048), .A2(new_n1120), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT118), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1121), .A2(new_n1128), .A3(new_n1122), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1124), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1111), .A2(new_n1113), .A3(new_n1116), .A4(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n995), .B1(new_n1071), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n990), .A2(new_n991), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT48), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n986), .A2(new_n989), .A3(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n825), .A2(G2067), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1136), .B1(new_n986), .B2(new_n987), .ZN(new_n1137));
  INV_X1    g712(.A(new_n985), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1135), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT46), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1140), .A2(KEYINPUT125), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n813), .A2(new_n981), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1141), .B1(new_n985), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1140), .A2(KEYINPUT125), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n977), .A2(new_n978), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1144), .B1(new_n977), .B2(new_n978), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1143), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT126), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT126), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1143), .B(new_n1149), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(KEYINPUT47), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT47), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1148), .A2(new_n1153), .A3(new_n1150), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1139), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1132), .A2(new_n1155), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g731(.A1(G401), .A2(G227), .ZN(new_n1158));
  AND2_X1   g732(.A1(new_n1158), .A2(new_n881), .ZN(new_n1159));
  AOI21_X1  g733(.A(new_n464), .B1(new_n957), .B2(new_n959), .ZN(new_n1160));
  NAND4_X1  g734(.A1(new_n1159), .A2(KEYINPUT127), .A3(new_n702), .A4(new_n1160), .ZN(new_n1161));
  NAND4_X1  g735(.A1(new_n702), .A2(new_n1158), .A3(new_n881), .A4(new_n1160), .ZN(G225));
  INV_X1    g736(.A(KEYINPUT127), .ZN(new_n1163));
  NAND2_X1  g737(.A1(G225), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g738(.A1(new_n1161), .A2(new_n1164), .ZN(G308));
endmodule


