

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U556 ( .A(KEYINPUT101), .B(n692), .Z(n521) );
  NAND2_X1 U557 ( .A1(n624), .A2(G2072), .ZN(n594) );
  XNOR2_X1 U558 ( .A(n594), .B(KEYINPUT95), .ZN(n596) );
  INV_X1 U559 ( .A(KEYINPUT97), .ZN(n644) );
  NOR2_X1 U560 ( .A1(n971), .A2(n601), .ZN(n600) );
  INV_X1 U561 ( .A(KEYINPUT29), .ZN(n636) );
  XNOR2_X1 U562 ( .A(n637), .B(n636), .ZN(n641) );
  NAND2_X1 U563 ( .A1(n700), .A2(n702), .ZN(n655) );
  INV_X1 U564 ( .A(KEYINPUT102), .ZN(n694) );
  NOR2_X1 U565 ( .A1(G651), .A2(n546), .ZN(n791) );
  XOR2_X1 U566 ( .A(KEYINPUT17), .B(n528), .Z(n873) );
  NOR2_X1 U567 ( .A1(n532), .A2(n531), .ZN(G164) );
  AND2_X1 U568 ( .A1(G2105), .A2(G2104), .ZN(n877) );
  NAND2_X1 U569 ( .A1(G114), .A2(n877), .ZN(n522) );
  XNOR2_X1 U570 ( .A(n522), .B(KEYINPUT88), .ZN(n526) );
  INV_X1 U571 ( .A(G2105), .ZN(n527) );
  AND2_X1 U572 ( .A1(n527), .A2(G2104), .ZN(n523) );
  XNOR2_X2 U573 ( .A(n523), .B(KEYINPUT64), .ZN(n874) );
  NAND2_X1 U574 ( .A1(n874), .A2(G102), .ZN(n524) );
  XOR2_X1 U575 ( .A(KEYINPUT89), .B(n524), .Z(n525) );
  NAND2_X1 U576 ( .A1(n526), .A2(n525), .ZN(n532) );
  NOR2_X1 U577 ( .A1(G2104), .A2(n527), .ZN(n878) );
  NAND2_X1 U578 ( .A1(G126), .A2(n878), .ZN(n530) );
  NOR2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n528) );
  NAND2_X1 U580 ( .A1(G138), .A2(n873), .ZN(n529) );
  NAND2_X1 U581 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U582 ( .A(KEYINPUT0), .B(G543), .Z(n546) );
  INV_X1 U583 ( .A(G651), .ZN(n536) );
  NOR2_X1 U584 ( .A1(n546), .A2(n536), .ZN(n795) );
  NAND2_X1 U585 ( .A1(G73), .A2(n795), .ZN(n533) );
  XNOR2_X1 U586 ( .A(n533), .B(KEYINPUT2), .ZN(n542) );
  NOR2_X1 U587 ( .A1(G651), .A2(G543), .ZN(n796) );
  NAND2_X1 U588 ( .A1(G86), .A2(n796), .ZN(n535) );
  NAND2_X1 U589 ( .A1(G48), .A2(n791), .ZN(n534) );
  NAND2_X1 U590 ( .A1(n535), .A2(n534), .ZN(n540) );
  NOR2_X1 U591 ( .A1(G543), .A2(n536), .ZN(n537) );
  XOR2_X1 U592 ( .A(KEYINPUT1), .B(n537), .Z(n790) );
  NAND2_X1 U593 ( .A1(G61), .A2(n790), .ZN(n538) );
  XNOR2_X1 U594 ( .A(KEYINPUT83), .B(n538), .ZN(n539) );
  NOR2_X1 U595 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U596 ( .A1(n542), .A2(n541), .ZN(G305) );
  NAND2_X1 U597 ( .A1(G49), .A2(n791), .ZN(n544) );
  NAND2_X1 U598 ( .A1(G74), .A2(G651), .ZN(n543) );
  NAND2_X1 U599 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U600 ( .A1(n790), .A2(n545), .ZN(n548) );
  NAND2_X1 U601 ( .A1(n546), .A2(G87), .ZN(n547) );
  NAND2_X1 U602 ( .A1(n548), .A2(n547), .ZN(G288) );
  NAND2_X1 U603 ( .A1(G75), .A2(n795), .ZN(n550) );
  NAND2_X1 U604 ( .A1(G88), .A2(n796), .ZN(n549) );
  NAND2_X1 U605 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U606 ( .A1(G62), .A2(n790), .ZN(n552) );
  NAND2_X1 U607 ( .A1(G50), .A2(n791), .ZN(n551) );
  NAND2_X1 U608 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U609 ( .A1(n554), .A2(n553), .ZN(G166) );
  INV_X1 U610 ( .A(G166), .ZN(G303) );
  NAND2_X1 U611 ( .A1(G77), .A2(n795), .ZN(n556) );
  NAND2_X1 U612 ( .A1(G90), .A2(n796), .ZN(n555) );
  NAND2_X1 U613 ( .A1(n556), .A2(n555), .ZN(n558) );
  XOR2_X1 U614 ( .A(KEYINPUT9), .B(KEYINPUT68), .Z(n557) );
  XNOR2_X1 U615 ( .A(n558), .B(n557), .ZN(n563) );
  NAND2_X1 U616 ( .A1(G64), .A2(n790), .ZN(n560) );
  NAND2_X1 U617 ( .A1(G52), .A2(n791), .ZN(n559) );
  NAND2_X1 U618 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U619 ( .A(KEYINPUT67), .B(n561), .Z(n562) );
  NOR2_X1 U620 ( .A1(n563), .A2(n562), .ZN(G171) );
  NAND2_X1 U621 ( .A1(n796), .A2(G89), .ZN(n564) );
  XNOR2_X1 U622 ( .A(n564), .B(KEYINPUT4), .ZN(n566) );
  NAND2_X1 U623 ( .A1(G76), .A2(n795), .ZN(n565) );
  NAND2_X1 U624 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U625 ( .A(n567), .B(KEYINPUT5), .ZN(n572) );
  NAND2_X1 U626 ( .A1(G63), .A2(n790), .ZN(n569) );
  NAND2_X1 U627 ( .A1(G51), .A2(n791), .ZN(n568) );
  NAND2_X1 U628 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U629 ( .A(KEYINPUT6), .B(n570), .Z(n571) );
  NAND2_X1 U630 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U631 ( .A(n573), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U632 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U633 ( .A1(G72), .A2(n795), .ZN(n575) );
  NAND2_X1 U634 ( .A1(G85), .A2(n796), .ZN(n574) );
  NAND2_X1 U635 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U636 ( .A1(G47), .A2(n791), .ZN(n576) );
  XOR2_X1 U637 ( .A(KEYINPUT66), .B(n576), .Z(n577) );
  NOR2_X1 U638 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U639 ( .A1(n790), .A2(G60), .ZN(n579) );
  NAND2_X1 U640 ( .A1(n580), .A2(n579), .ZN(G290) );
  XOR2_X1 U641 ( .A(G1981), .B(G305), .Z(n987) );
  NOR2_X1 U642 ( .A1(G1976), .A2(G288), .ZN(n973) );
  OR2_X1 U643 ( .A1(G1971), .A2(G303), .ZN(n970) );
  XOR2_X1 U644 ( .A(KEYINPUT99), .B(n970), .Z(n672) );
  NAND2_X1 U645 ( .A1(G65), .A2(n790), .ZN(n582) );
  NAND2_X1 U646 ( .A1(G53), .A2(n791), .ZN(n581) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U648 ( .A1(G78), .A2(n795), .ZN(n584) );
  NAND2_X1 U649 ( .A1(G91), .A2(n796), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n971) );
  NAND2_X1 U652 ( .A1(G113), .A2(n877), .ZN(n588) );
  NAND2_X1 U653 ( .A1(G125), .A2(n878), .ZN(n587) );
  AND2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n755) );
  AND2_X1 U655 ( .A1(n755), .A2(G40), .ZN(n593) );
  NAND2_X1 U656 ( .A1(n874), .A2(G101), .ZN(n589) );
  XNOR2_X1 U657 ( .A(n589), .B(KEYINPUT23), .ZN(n590) );
  XNOR2_X1 U658 ( .A(n590), .B(KEYINPUT65), .ZN(n592) );
  NAND2_X1 U659 ( .A1(G137), .A2(n873), .ZN(n591) );
  AND2_X1 U660 ( .A1(n592), .A2(n591), .ZN(n754) );
  AND2_X1 U661 ( .A1(n593), .A2(n754), .ZN(n700) );
  NOR2_X1 U662 ( .A1(G164), .A2(G1384), .ZN(n702) );
  INV_X1 U663 ( .A(n655), .ZN(n624) );
  INV_X1 U664 ( .A(KEYINPUT27), .ZN(n595) );
  XNOR2_X1 U665 ( .A(n596), .B(n595), .ZN(n599) );
  NAND2_X1 U666 ( .A1(G1956), .A2(n655), .ZN(n597) );
  XOR2_X1 U667 ( .A(KEYINPUT96), .B(n597), .Z(n598) );
  NOR2_X1 U668 ( .A1(n599), .A2(n598), .ZN(n601) );
  XOR2_X1 U669 ( .A(n600), .B(KEYINPUT28), .Z(n635) );
  NAND2_X1 U670 ( .A1(n971), .A2(n601), .ZN(n633) );
  NAND2_X1 U671 ( .A1(G56), .A2(n790), .ZN(n602) );
  XOR2_X1 U672 ( .A(KEYINPUT14), .B(n602), .Z(n609) );
  NAND2_X1 U673 ( .A1(n796), .A2(G81), .ZN(n603) );
  XOR2_X1 U674 ( .A(KEYINPUT12), .B(n603), .Z(n606) );
  NAND2_X1 U675 ( .A1(n795), .A2(G68), .ZN(n604) );
  XOR2_X1 U676 ( .A(KEYINPUT72), .B(n604), .Z(n605) );
  NOR2_X1 U677 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U678 ( .A(n607), .B(KEYINPUT13), .ZN(n608) );
  NOR2_X1 U679 ( .A1(n609), .A2(n608), .ZN(n611) );
  NAND2_X1 U680 ( .A1(n791), .A2(G43), .ZN(n610) );
  NAND2_X1 U681 ( .A1(n611), .A2(n610), .ZN(n982) );
  AND2_X1 U682 ( .A1(n624), .A2(G1996), .ZN(n612) );
  XOR2_X1 U683 ( .A(n612), .B(KEYINPUT26), .Z(n614) );
  NAND2_X1 U684 ( .A1(n655), .A2(G1341), .ZN(n613) );
  NAND2_X1 U685 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U686 ( .A1(n982), .A2(n615), .ZN(n628) );
  NAND2_X1 U687 ( .A1(G92), .A2(n796), .ZN(n617) );
  NAND2_X1 U688 ( .A1(G66), .A2(n790), .ZN(n616) );
  NAND2_X1 U689 ( .A1(n617), .A2(n616), .ZN(n622) );
  NAND2_X1 U690 ( .A1(G79), .A2(n795), .ZN(n619) );
  NAND2_X1 U691 ( .A1(G54), .A2(n791), .ZN(n618) );
  NAND2_X1 U692 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U693 ( .A(KEYINPUT74), .B(n620), .ZN(n621) );
  NOR2_X1 U694 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U695 ( .A(n623), .B(KEYINPUT15), .ZN(n986) );
  NAND2_X1 U696 ( .A1(G1348), .A2(n655), .ZN(n626) );
  NAND2_X1 U697 ( .A1(G2067), .A2(n624), .ZN(n625) );
  NAND2_X1 U698 ( .A1(n626), .A2(n625), .ZN(n629) );
  NOR2_X1 U699 ( .A1(n986), .A2(n629), .ZN(n627) );
  OR2_X1 U700 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U701 ( .A1(n986), .A2(n629), .ZN(n630) );
  NAND2_X1 U702 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U703 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U704 ( .A1(n635), .A2(n634), .ZN(n637) );
  XNOR2_X1 U705 ( .A(G2078), .B(KEYINPUT25), .ZN(n955) );
  NOR2_X1 U706 ( .A1(n655), .A2(n955), .ZN(n639) );
  AND2_X1 U707 ( .A1(n655), .A2(G1961), .ZN(n638) );
  NOR2_X1 U708 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U709 ( .A1(G171), .A2(n642), .ZN(n640) );
  NAND2_X1 U710 ( .A1(n641), .A2(n640), .ZN(n654) );
  INV_X1 U711 ( .A(KEYINPUT31), .ZN(n652) );
  NOR2_X1 U712 ( .A1(G171), .A2(n642), .ZN(n650) );
  NAND2_X1 U713 ( .A1(G8), .A2(n655), .ZN(n693) );
  NOR2_X1 U714 ( .A1(G1966), .A2(n693), .ZN(n667) );
  NOR2_X1 U715 ( .A1(n655), .A2(G2084), .ZN(n643) );
  XNOR2_X1 U716 ( .A(n643), .B(KEYINPUT94), .ZN(n664) );
  NOR2_X1 U717 ( .A1(n667), .A2(n664), .ZN(n645) );
  XNOR2_X1 U718 ( .A(n645), .B(n644), .ZN(n646) );
  NAND2_X1 U719 ( .A1(n646), .A2(G8), .ZN(n647) );
  XNOR2_X1 U720 ( .A(KEYINPUT30), .B(n647), .ZN(n648) );
  NOR2_X1 U721 ( .A1(G168), .A2(n648), .ZN(n649) );
  NOR2_X1 U722 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U723 ( .A(n652), .B(n651), .ZN(n653) );
  NAND2_X1 U724 ( .A1(n654), .A2(n653), .ZN(n665) );
  NAND2_X1 U725 ( .A1(n665), .A2(G286), .ZN(n661) );
  NOR2_X1 U726 ( .A1(G1971), .A2(n693), .ZN(n657) );
  NOR2_X1 U727 ( .A1(G2090), .A2(n655), .ZN(n656) );
  NOR2_X1 U728 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U729 ( .A(n658), .B(KEYINPUT98), .ZN(n659) );
  NAND2_X1 U730 ( .A1(n659), .A2(G303), .ZN(n660) );
  NAND2_X1 U731 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U732 ( .A1(n662), .A2(G8), .ZN(n663) );
  XNOR2_X1 U733 ( .A(n663), .B(KEYINPUT32), .ZN(n671) );
  NAND2_X1 U734 ( .A1(n664), .A2(G8), .ZN(n669) );
  INV_X1 U735 ( .A(n665), .ZN(n666) );
  NOR2_X1 U736 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U737 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U738 ( .A1(n671), .A2(n670), .ZN(n691) );
  NAND2_X1 U739 ( .A1(n672), .A2(n691), .ZN(n673) );
  NOR2_X1 U740 ( .A1(KEYINPUT33), .A2(n673), .ZN(n675) );
  NOR2_X1 U741 ( .A1(n693), .A2(KEYINPUT100), .ZN(n674) );
  NOR2_X1 U742 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U743 ( .A1(n973), .A2(n676), .ZN(n685) );
  NAND2_X1 U744 ( .A1(G1976), .A2(G288), .ZN(n969) );
  INV_X1 U745 ( .A(KEYINPUT100), .ZN(n677) );
  NOR2_X1 U746 ( .A1(n693), .A2(n677), .ZN(n680) );
  NAND2_X1 U747 ( .A1(n969), .A2(n680), .ZN(n679) );
  INV_X1 U748 ( .A(KEYINPUT33), .ZN(n678) );
  NAND2_X1 U749 ( .A1(n679), .A2(n678), .ZN(n683) );
  AND2_X1 U750 ( .A1(n973), .A2(KEYINPUT33), .ZN(n681) );
  NAND2_X1 U751 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U752 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U753 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U754 ( .A1(n987), .A2(n686), .ZN(n699) );
  NOR2_X1 U755 ( .A1(G1981), .A2(G305), .ZN(n687) );
  XOR2_X1 U756 ( .A(n687), .B(KEYINPUT24), .Z(n688) );
  NOR2_X1 U757 ( .A1(n693), .A2(n688), .ZN(n697) );
  NOR2_X1 U758 ( .A1(G2090), .A2(G303), .ZN(n689) );
  NAND2_X1 U759 ( .A1(G8), .A2(n689), .ZN(n690) );
  NAND2_X1 U760 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U761 ( .A1(n521), .A2(n693), .ZN(n695) );
  XNOR2_X1 U762 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X1 U763 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U764 ( .A1(n699), .A2(n698), .ZN(n735) );
  INV_X1 U765 ( .A(n700), .ZN(n701) );
  NOR2_X1 U766 ( .A1(n702), .A2(n701), .ZN(n749) );
  NAND2_X1 U767 ( .A1(n873), .A2(G140), .ZN(n704) );
  NAND2_X1 U768 ( .A1(G104), .A2(n874), .ZN(n703) );
  NAND2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U770 ( .A(KEYINPUT34), .B(n705), .ZN(n710) );
  NAND2_X1 U771 ( .A1(G116), .A2(n877), .ZN(n707) );
  NAND2_X1 U772 ( .A1(G128), .A2(n878), .ZN(n706) );
  NAND2_X1 U773 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U774 ( .A(n708), .B(KEYINPUT35), .Z(n709) );
  NOR2_X1 U775 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U776 ( .A(KEYINPUT36), .B(n711), .Z(n712) );
  XOR2_X1 U777 ( .A(KEYINPUT90), .B(n712), .Z(n895) );
  XNOR2_X1 U778 ( .A(KEYINPUT37), .B(G2067), .ZN(n736) );
  NOR2_X1 U779 ( .A1(n895), .A2(n736), .ZN(n932) );
  NAND2_X1 U780 ( .A1(n749), .A2(n932), .ZN(n747) );
  NAND2_X1 U781 ( .A1(n874), .A2(G105), .ZN(n713) );
  XNOR2_X1 U782 ( .A(n713), .B(KEYINPUT38), .ZN(n720) );
  NAND2_X1 U783 ( .A1(G117), .A2(n877), .ZN(n715) );
  NAND2_X1 U784 ( .A1(G129), .A2(n878), .ZN(n714) );
  NAND2_X1 U785 ( .A1(n715), .A2(n714), .ZN(n718) );
  NAND2_X1 U786 ( .A1(n873), .A2(G141), .ZN(n716) );
  XOR2_X1 U787 ( .A(KEYINPUT92), .B(n716), .Z(n717) );
  NOR2_X1 U788 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U789 ( .A1(n720), .A2(n719), .ZN(n891) );
  NAND2_X1 U790 ( .A1(G1996), .A2(n891), .ZN(n729) );
  NAND2_X1 U791 ( .A1(G107), .A2(n877), .ZN(n722) );
  NAND2_X1 U792 ( .A1(G131), .A2(n873), .ZN(n721) );
  NAND2_X1 U793 ( .A1(n722), .A2(n721), .ZN(n725) );
  NAND2_X1 U794 ( .A1(G119), .A2(n878), .ZN(n723) );
  XNOR2_X1 U795 ( .A(KEYINPUT91), .B(n723), .ZN(n724) );
  NOR2_X1 U796 ( .A1(n725), .A2(n724), .ZN(n727) );
  NAND2_X1 U797 ( .A1(G95), .A2(n874), .ZN(n726) );
  NAND2_X1 U798 ( .A1(n727), .A2(n726), .ZN(n886) );
  NAND2_X1 U799 ( .A1(G1991), .A2(n886), .ZN(n728) );
  NAND2_X1 U800 ( .A1(n729), .A2(n728), .ZN(n936) );
  NAND2_X1 U801 ( .A1(n936), .A2(n749), .ZN(n730) );
  XNOR2_X1 U802 ( .A(n730), .B(KEYINPUT93), .ZN(n742) );
  INV_X1 U803 ( .A(n742), .ZN(n731) );
  NAND2_X1 U804 ( .A1(n747), .A2(n731), .ZN(n733) );
  XNOR2_X1 U805 ( .A(G1986), .B(G290), .ZN(n979) );
  AND2_X1 U806 ( .A1(n979), .A2(n749), .ZN(n732) );
  NOR2_X1 U807 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U808 ( .A1(n735), .A2(n734), .ZN(n752) );
  NAND2_X1 U809 ( .A1(n895), .A2(n736), .ZN(n737) );
  XNOR2_X1 U810 ( .A(n737), .B(KEYINPUT106), .ZN(n939) );
  XNOR2_X1 U811 ( .A(KEYINPUT105), .B(KEYINPUT39), .ZN(n745) );
  NOR2_X1 U812 ( .A1(G1991), .A2(n886), .ZN(n930) );
  NOR2_X1 U813 ( .A1(G1986), .A2(G290), .ZN(n738) );
  XOR2_X1 U814 ( .A(n738), .B(KEYINPUT103), .Z(n739) );
  NOR2_X1 U815 ( .A1(n930), .A2(n739), .ZN(n740) );
  XNOR2_X1 U816 ( .A(n740), .B(KEYINPUT104), .ZN(n741) );
  NOR2_X1 U817 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U818 ( .A1(G1996), .A2(n891), .ZN(n925) );
  NOR2_X1 U819 ( .A1(n743), .A2(n925), .ZN(n744) );
  XOR2_X1 U820 ( .A(n745), .B(n744), .Z(n746) );
  NAND2_X1 U821 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U822 ( .A1(n939), .A2(n748), .ZN(n750) );
  NAND2_X1 U823 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U824 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U825 ( .A(n753), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U826 ( .A1(n755), .A2(n754), .ZN(G160) );
  INV_X1 U827 ( .A(G132), .ZN(G219) );
  INV_X1 U828 ( .A(G82), .ZN(G220) );
  INV_X1 U829 ( .A(G120), .ZN(G236) );
  INV_X1 U830 ( .A(G69), .ZN(G235) );
  INV_X1 U831 ( .A(G108), .ZN(G238) );
  NAND2_X1 U832 ( .A1(G94), .A2(G452), .ZN(n756) );
  XNOR2_X1 U833 ( .A(n756), .B(KEYINPUT69), .ZN(G173) );
  NAND2_X1 U834 ( .A1(G7), .A2(G661), .ZN(n757) );
  XNOR2_X1 U835 ( .A(n757), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U836 ( .A(G223), .ZN(n829) );
  NAND2_X1 U837 ( .A1(n829), .A2(G567), .ZN(n758) );
  XNOR2_X1 U838 ( .A(n758), .B(KEYINPUT71), .ZN(n759) );
  XNOR2_X1 U839 ( .A(KEYINPUT11), .B(n759), .ZN(G234) );
  INV_X1 U840 ( .A(n982), .ZN(n760) );
  NAND2_X1 U841 ( .A1(n760), .A2(G860), .ZN(G153) );
  INV_X1 U842 ( .A(G868), .ZN(n764) );
  NOR2_X1 U843 ( .A1(n764), .A2(G171), .ZN(n761) );
  XNOR2_X1 U844 ( .A(n761), .B(KEYINPUT73), .ZN(n763) );
  NAND2_X1 U845 ( .A1(n764), .A2(n986), .ZN(n762) );
  NAND2_X1 U846 ( .A1(n763), .A2(n762), .ZN(G284) );
  XOR2_X1 U847 ( .A(n971), .B(KEYINPUT70), .Z(G299) );
  NOR2_X1 U848 ( .A1(G286), .A2(n764), .ZN(n766) );
  NOR2_X1 U849 ( .A1(G299), .A2(G868), .ZN(n765) );
  NOR2_X1 U850 ( .A1(n766), .A2(n765), .ZN(G297) );
  INV_X1 U851 ( .A(G559), .ZN(n767) );
  NOR2_X1 U852 ( .A1(G860), .A2(n767), .ZN(n768) );
  XNOR2_X1 U853 ( .A(KEYINPUT75), .B(n768), .ZN(n769) );
  INV_X1 U854 ( .A(n986), .ZN(n788) );
  NAND2_X1 U855 ( .A1(n769), .A2(n788), .ZN(n770) );
  XNOR2_X1 U856 ( .A(n770), .B(KEYINPUT16), .ZN(n771) );
  XNOR2_X1 U857 ( .A(KEYINPUT76), .B(n771), .ZN(G148) );
  NAND2_X1 U858 ( .A1(n788), .A2(G868), .ZN(n772) );
  XOR2_X1 U859 ( .A(KEYINPUT77), .B(n772), .Z(n773) );
  NOR2_X1 U860 ( .A1(G559), .A2(n773), .ZN(n775) );
  NOR2_X1 U861 ( .A1(G868), .A2(n982), .ZN(n774) );
  NOR2_X1 U862 ( .A1(n775), .A2(n774), .ZN(G282) );
  NAND2_X1 U863 ( .A1(n878), .A2(G123), .ZN(n776) );
  XNOR2_X1 U864 ( .A(n776), .B(KEYINPUT18), .ZN(n778) );
  NAND2_X1 U865 ( .A1(G135), .A2(n873), .ZN(n777) );
  NAND2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U867 ( .A(KEYINPUT78), .B(n779), .Z(n781) );
  NAND2_X1 U868 ( .A1(n877), .A2(G111), .ZN(n780) );
  NAND2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n784) );
  NAND2_X1 U870 ( .A1(G99), .A2(n874), .ZN(n782) );
  XNOR2_X1 U871 ( .A(KEYINPUT79), .B(n782), .ZN(n783) );
  NOR2_X1 U872 ( .A1(n784), .A2(n783), .ZN(n929) );
  XNOR2_X1 U873 ( .A(n929), .B(G2096), .ZN(n785) );
  XNOR2_X1 U874 ( .A(n785), .B(KEYINPUT80), .ZN(n787) );
  INV_X1 U875 ( .A(G2100), .ZN(n786) );
  NAND2_X1 U876 ( .A1(n787), .A2(n786), .ZN(G156) );
  NAND2_X1 U877 ( .A1(G559), .A2(n788), .ZN(n789) );
  XNOR2_X1 U878 ( .A(n789), .B(n982), .ZN(n811) );
  NOR2_X1 U879 ( .A1(n811), .A2(G860), .ZN(n802) );
  NAND2_X1 U880 ( .A1(G67), .A2(n790), .ZN(n793) );
  NAND2_X1 U881 ( .A1(G55), .A2(n791), .ZN(n792) );
  NAND2_X1 U882 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U883 ( .A(KEYINPUT82), .B(n794), .ZN(n801) );
  NAND2_X1 U884 ( .A1(G80), .A2(n795), .ZN(n798) );
  NAND2_X1 U885 ( .A1(G93), .A2(n796), .ZN(n797) );
  NAND2_X1 U886 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U887 ( .A(KEYINPUT81), .B(n799), .Z(n800) );
  NOR2_X1 U888 ( .A1(n801), .A2(n800), .ZN(n806) );
  XNOR2_X1 U889 ( .A(n802), .B(n806), .ZN(G145) );
  NOR2_X1 U890 ( .A1(G868), .A2(n806), .ZN(n803) );
  XNOR2_X1 U891 ( .A(n803), .B(KEYINPUT85), .ZN(n814) );
  XOR2_X1 U892 ( .A(KEYINPUT84), .B(KEYINPUT19), .Z(n804) );
  XNOR2_X1 U893 ( .A(G288), .B(n804), .ZN(n805) );
  XNOR2_X1 U894 ( .A(G299), .B(n805), .ZN(n808) );
  XNOR2_X1 U895 ( .A(G305), .B(n806), .ZN(n807) );
  XNOR2_X1 U896 ( .A(n808), .B(n807), .ZN(n809) );
  XNOR2_X1 U897 ( .A(G166), .B(n809), .ZN(n810) );
  XNOR2_X1 U898 ( .A(n810), .B(G290), .ZN(n899) );
  XNOR2_X1 U899 ( .A(n899), .B(n811), .ZN(n812) );
  NAND2_X1 U900 ( .A1(G868), .A2(n812), .ZN(n813) );
  NAND2_X1 U901 ( .A1(n814), .A2(n813), .ZN(G295) );
  NAND2_X1 U902 ( .A1(G2078), .A2(G2084), .ZN(n815) );
  XOR2_X1 U903 ( .A(KEYINPUT20), .B(n815), .Z(n816) );
  NAND2_X1 U904 ( .A1(G2090), .A2(n816), .ZN(n817) );
  XNOR2_X1 U905 ( .A(KEYINPUT21), .B(n817), .ZN(n818) );
  NAND2_X1 U906 ( .A1(n818), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U907 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U908 ( .A1(G235), .A2(G236), .ZN(n819) );
  XOR2_X1 U909 ( .A(KEYINPUT86), .B(n819), .Z(n820) );
  NOR2_X1 U910 ( .A1(G238), .A2(n820), .ZN(n821) );
  NAND2_X1 U911 ( .A1(G57), .A2(n821), .ZN(n834) );
  NAND2_X1 U912 ( .A1(n834), .A2(G567), .ZN(n826) );
  NOR2_X1 U913 ( .A1(G220), .A2(G219), .ZN(n822) );
  XOR2_X1 U914 ( .A(KEYINPUT22), .B(n822), .Z(n823) );
  NOR2_X1 U915 ( .A1(G218), .A2(n823), .ZN(n824) );
  NAND2_X1 U916 ( .A1(G96), .A2(n824), .ZN(n835) );
  NAND2_X1 U917 ( .A1(n835), .A2(G2106), .ZN(n825) );
  NAND2_X1 U918 ( .A1(n826), .A2(n825), .ZN(n836) );
  NAND2_X1 U919 ( .A1(G661), .A2(G483), .ZN(n827) );
  NOR2_X1 U920 ( .A1(n836), .A2(n827), .ZN(n828) );
  XOR2_X1 U921 ( .A(KEYINPUT87), .B(n828), .Z(n833) );
  NAND2_X1 U922 ( .A1(n833), .A2(G36), .ZN(G176) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n829), .ZN(G217) );
  NAND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n830) );
  XOR2_X1 U925 ( .A(KEYINPUT108), .B(n830), .Z(n831) );
  NAND2_X1 U926 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U928 ( .A1(n833), .A2(n832), .ZN(G188) );
  XNOR2_X1 U929 ( .A(G96), .B(KEYINPUT109), .ZN(G221) );
  NOR2_X1 U931 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  INV_X1 U933 ( .A(n836), .ZN(G319) );
  XOR2_X1 U934 ( .A(KEYINPUT110), .B(KEYINPUT112), .Z(n838) );
  XNOR2_X1 U935 ( .A(G2678), .B(G2100), .ZN(n837) );
  XNOR2_X1 U936 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U937 ( .A(n839), .B(KEYINPUT111), .Z(n841) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2072), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U940 ( .A(G2096), .B(G2090), .Z(n843) );
  XNOR2_X1 U941 ( .A(G2078), .B(G2084), .ZN(n842) );
  XNOR2_X1 U942 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U943 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U944 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n846) );
  XNOR2_X1 U945 ( .A(n847), .B(n846), .ZN(G227) );
  XOR2_X1 U946 ( .A(G1971), .B(G1961), .Z(n849) );
  XNOR2_X1 U947 ( .A(G1986), .B(G1976), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U949 ( .A(G1966), .B(G1981), .Z(n851) );
  XNOR2_X1 U950 ( .A(G1996), .B(G1991), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U952 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U953 ( .A(KEYINPUT113), .B(KEYINPUT41), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n857) );
  XOR2_X1 U955 ( .A(G1956), .B(G2474), .Z(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(G229) );
  NAND2_X1 U957 ( .A1(G124), .A2(n878), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n858), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U959 ( .A1(n877), .A2(G112), .ZN(n859) );
  NAND2_X1 U960 ( .A1(n860), .A2(n859), .ZN(n864) );
  NAND2_X1 U961 ( .A1(n873), .A2(G136), .ZN(n862) );
  NAND2_X1 U962 ( .A1(G100), .A2(n874), .ZN(n861) );
  NAND2_X1 U963 ( .A1(n862), .A2(n861), .ZN(n863) );
  NOR2_X1 U964 ( .A1(n864), .A2(n863), .ZN(G162) );
  NAND2_X1 U965 ( .A1(G118), .A2(n877), .ZN(n866) );
  NAND2_X1 U966 ( .A1(G130), .A2(n878), .ZN(n865) );
  NAND2_X1 U967 ( .A1(n866), .A2(n865), .ZN(n871) );
  NAND2_X1 U968 ( .A1(n873), .A2(G142), .ZN(n868) );
  NAND2_X1 U969 ( .A1(G106), .A2(n874), .ZN(n867) );
  NAND2_X1 U970 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U971 ( .A(KEYINPUT45), .B(n869), .Z(n870) );
  NOR2_X1 U972 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U973 ( .A(n929), .B(n872), .ZN(n890) );
  NAND2_X1 U974 ( .A1(n873), .A2(G139), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G103), .A2(n874), .ZN(n875) );
  NAND2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n884) );
  NAND2_X1 U977 ( .A1(G115), .A2(n877), .ZN(n880) );
  NAND2_X1 U978 ( .A1(G127), .A2(n878), .ZN(n879) );
  NAND2_X1 U979 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U980 ( .A(KEYINPUT114), .B(n881), .Z(n882) );
  XNOR2_X1 U981 ( .A(KEYINPUT47), .B(n882), .ZN(n883) );
  NOR2_X1 U982 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U983 ( .A(KEYINPUT115), .B(n885), .Z(n920) );
  XNOR2_X1 U984 ( .A(n886), .B(n920), .ZN(n888) );
  XNOR2_X1 U985 ( .A(G164), .B(G160), .ZN(n887) );
  XNOR2_X1 U986 ( .A(n888), .B(n887), .ZN(n889) );
  XNOR2_X1 U987 ( .A(n890), .B(n889), .ZN(n897) );
  XNOR2_X1 U988 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n893) );
  XNOR2_X1 U989 ( .A(n891), .B(G162), .ZN(n892) );
  XNOR2_X1 U990 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U991 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U992 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U993 ( .A1(G37), .A2(n898), .ZN(G395) );
  XNOR2_X1 U994 ( .A(G286), .B(n982), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n902) );
  XNOR2_X1 U996 ( .A(n986), .B(G171), .ZN(n901) );
  XNOR2_X1 U997 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U998 ( .A1(G37), .A2(n903), .ZN(G397) );
  XOR2_X1 U999 ( .A(G2430), .B(G2451), .Z(n905) );
  XNOR2_X1 U1000 ( .A(G2446), .B(G2427), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n912) );
  XOR2_X1 U1002 ( .A(G2438), .B(G2435), .Z(n907) );
  XNOR2_X1 U1003 ( .A(G2443), .B(KEYINPUT107), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1005 ( .A(n908), .B(G2454), .Z(n910) );
  XNOR2_X1 U1006 ( .A(G1341), .B(G1348), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(n912), .B(n911), .ZN(n913) );
  NAND2_X1 U1009 ( .A1(n913), .A2(G14), .ZN(n919) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n919), .ZN(n916) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n914), .ZN(n915) );
  NOR2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G171), .ZN(G301) );
  INV_X1 U1018 ( .A(G57), .ZN(G237) );
  INV_X1 U1019 ( .A(n919), .ZN(G401) );
  XOR2_X1 U1020 ( .A(G2072), .B(n920), .Z(n922) );
  XOR2_X1 U1021 ( .A(G164), .B(G2078), .Z(n921) );
  NOR2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1023 ( .A(KEYINPUT50), .B(n923), .ZN(n928) );
  XOR2_X1 U1024 ( .A(G2090), .B(G162), .Z(n924) );
  NOR2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1026 ( .A(KEYINPUT51), .B(n926), .Z(n927) );
  NAND2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n941) );
  NOR2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n934) );
  XOR2_X1 U1029 ( .A(G160), .B(G2084), .Z(n931) );
  NOR2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1033 ( .A(n937), .B(KEYINPUT116), .ZN(n938) );
  NAND2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1036 ( .A(KEYINPUT52), .B(n942), .ZN(n944) );
  INV_X1 U1037 ( .A(KEYINPUT55), .ZN(n943) );
  NAND2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1039 ( .A1(n945), .A2(G29), .ZN(n946) );
  XOR2_X1 U1040 ( .A(KEYINPUT117), .B(n946), .Z(n1028) );
  XNOR2_X1 U1041 ( .A(G1996), .B(G32), .ZN(n948) );
  XNOR2_X1 U1042 ( .A(G33), .B(G2072), .ZN(n947) );
  NOR2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n954) );
  XOR2_X1 U1044 ( .A(G2067), .B(G26), .Z(n949) );
  NAND2_X1 U1045 ( .A1(n949), .A2(G28), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(G25), .B(G1991), .ZN(n950) );
  XNOR2_X1 U1047 ( .A(KEYINPUT118), .B(n950), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n957) );
  XOR2_X1 U1050 ( .A(G27), .B(n955), .Z(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(n958), .B(KEYINPUT119), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(n959), .B(KEYINPUT53), .ZN(n962) );
  XOR2_X1 U1054 ( .A(G2084), .B(G34), .Z(n960) );
  XNOR2_X1 U1055 ( .A(KEYINPUT54), .B(n960), .ZN(n961) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(G35), .B(G2090), .ZN(n963) );
  NOR2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1059 ( .A(KEYINPUT55), .B(n965), .Z(n966) );
  NOR2_X1 U1060 ( .A1(G29), .A2(n966), .ZN(n967) );
  XOR2_X1 U1061 ( .A(KEYINPUT120), .B(n967), .Z(n968) );
  NAND2_X1 U1062 ( .A1(G11), .A2(n968), .ZN(n1026) );
  XNOR2_X1 U1063 ( .A(G16), .B(KEYINPUT56), .ZN(n996) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n977) );
  XOR2_X1 U1065 ( .A(n971), .B(G1956), .Z(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n975) );
  NAND2_X1 U1067 ( .A1(G1971), .A2(G303), .ZN(n974) );
  NAND2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n981) );
  XNOR2_X1 U1070 ( .A(G1961), .B(G301), .ZN(n978) );
  NOR2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n985) );
  XNOR2_X1 U1073 ( .A(G1341), .B(n982), .ZN(n983) );
  XNOR2_X1 U1074 ( .A(KEYINPUT122), .B(n983), .ZN(n984) );
  NOR2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n994) );
  XNOR2_X1 U1076 ( .A(n986), .B(G1348), .ZN(n992) );
  XNOR2_X1 U1077 ( .A(G1966), .B(G168), .ZN(n988) );
  NAND2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(n989), .B(KEYINPUT57), .ZN(n990) );
  XNOR2_X1 U1080 ( .A(KEYINPUT121), .B(n990), .ZN(n991) );
  NOR2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n1024) );
  INV_X1 U1084 ( .A(G16), .ZN(n1022) );
  XOR2_X1 U1085 ( .A(G1971), .B(G22), .Z(n999) );
  XOR2_X1 U1086 ( .A(G24), .B(KEYINPUT126), .Z(n997) );
  XNOR2_X1 U1087 ( .A(n997), .B(G1986), .ZN(n998) );
  NAND2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1002) );
  XOR2_X1 U1089 ( .A(KEYINPUT125), .B(G1976), .Z(n1000) );
  XNOR2_X1 U1090 ( .A(G23), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1092 ( .A(KEYINPUT58), .B(n1003), .Z(n1019) );
  XNOR2_X1 U1093 ( .A(G1961), .B(G5), .ZN(n1016) );
  XNOR2_X1 U1094 ( .A(G1348), .B(KEYINPUT59), .ZN(n1004) );
  XNOR2_X1 U1095 ( .A(n1004), .B(G4), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(G1981), .B(G6), .ZN(n1006) );
  XNOR2_X1 U1097 ( .A(G1341), .B(G19), .ZN(n1005) );
  NOR2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(G20), .B(G1956), .ZN(n1009) );
  NOR2_X1 U1101 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1102 ( .A(KEYINPUT60), .B(n1011), .Z(n1013) );
  XNOR2_X1 U1103 ( .A(G1966), .B(G21), .ZN(n1012) );
  NOR2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1105 ( .A(KEYINPUT123), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1106 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1107 ( .A(KEYINPUT124), .B(n1017), .Z(n1018) );
  NOR2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1109 ( .A(KEYINPUT61), .B(n1020), .ZN(n1021) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1114 ( .A(n1029), .B(KEYINPUT127), .ZN(n1030) );
  XNOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1030), .ZN(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

