//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 1 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1223, new_n1224,
    new_n1225, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(new_n205));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  AND2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n210), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n202), .A2(new_n203), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(new_n214), .A2(new_n215), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  INV_X1    g0023(.A(G107), .ZN(new_n224));
  INV_X1    g0024(.A(G264), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n222), .B1(new_n202), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n212), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n221), .B1(new_n215), .B2(new_n214), .C1(new_n230), .C2(KEYINPUT1), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT65), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G169), .ZN(new_n249));
  AOI21_X1  g0049(.A(new_n249), .B1(KEYINPUT70), .B2(KEYINPUT14), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G33), .ZN(new_n254));
  AND2_X1   g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(G226), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(G232), .A3(G1698), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G97), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  OAI211_X1 g0061(.A(G1), .B(G13), .C1(new_n251), .C2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT13), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n266));
  INV_X1    g0066(.A(G274), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n262), .A2(new_n266), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n268), .B1(new_n270), .B2(G238), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n264), .A2(new_n265), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n265), .B1(new_n264), .B2(new_n271), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n250), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(KEYINPUT70), .A2(KEYINPUT14), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n274), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n272), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(new_n250), .A3(new_n276), .ZN(new_n281));
  INV_X1    g0081(.A(G179), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n278), .B(new_n281), .C1(new_n282), .C2(new_n280), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n209), .A2(G13), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G20), .A3(new_n203), .ZN(new_n286));
  XNOR2_X1  g0086(.A(new_n286), .B(KEYINPUT12), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n216), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n290), .B1(G1), .B2(new_n210), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n287), .B1(new_n203), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G20), .A2(G33), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n293), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n210), .A2(G33), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n294), .B1(new_n206), .B2(new_n295), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n296), .A2(KEYINPUT11), .A3(new_n289), .ZN(new_n297));
  AOI21_X1  g0097(.A(KEYINPUT11), .B1(new_n296), .B2(new_n289), .ZN(new_n298));
  OR3_X1    g0098(.A1(new_n292), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n283), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G200), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n280), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G190), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n279), .A2(new_n303), .A3(new_n272), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n299), .ZN(new_n306));
  AOI21_X1  g0106(.A(KEYINPUT69), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT69), .ZN(new_n308));
  AOI211_X1 g0108(.A(new_n308), .B(new_n299), .C1(new_n302), .C2(new_n304), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n300), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n293), .A2(G150), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT66), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G58), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT8), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n313), .B(new_n314), .ZN(new_n315));
  OAI221_X1 g0115(.A(new_n311), .B1(new_n315), .B2(new_n295), .C1(new_n205), .C2(new_n210), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n289), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n291), .A2(G50), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n318), .B1(G50), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n322), .B(KEYINPUT9), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n255), .A2(G222), .A3(new_n256), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n255), .A2(G1698), .ZN(new_n325));
  INV_X1    g0125(.A(G223), .ZN(new_n326));
  OAI221_X1 g0126(.A(new_n324), .B1(new_n206), .B2(new_n255), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n263), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n268), .B1(new_n270), .B2(G226), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n301), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(G190), .B2(new_n330), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n323), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT68), .ZN(new_n334));
  AOI21_X1  g0134(.A(KEYINPUT10), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n323), .B(new_n332), .C1(new_n334), .C2(KEYINPUT10), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n330), .A2(G169), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(new_n282), .B2(new_n330), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n322), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n336), .A2(new_n337), .A3(new_n340), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT15), .B(G87), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n342), .A2(new_n295), .B1(new_n210), .B2(new_n206), .ZN(new_n343));
  XOR2_X1   g0143(.A(KEYINPUT8), .B(G58), .Z(new_n344));
  XNOR2_X1  g0144(.A(new_n344), .B(KEYINPUT67), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n343), .B1(new_n345), .B2(new_n293), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n346), .A2(new_n290), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n320), .A2(G77), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(new_n291), .B2(G77), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n255), .A2(G232), .A3(new_n256), .ZN(new_n352));
  INV_X1    g0152(.A(G238), .ZN(new_n353));
  OAI221_X1 g0153(.A(new_n352), .B1(new_n224), .B2(new_n255), .C1(new_n325), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n263), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n268), .B1(new_n270), .B2(G244), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n303), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(new_n301), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n351), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n358), .A2(G179), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n357), .A2(G169), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n350), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NOR4_X1   g0164(.A1(new_n310), .A2(new_n341), .A3(new_n361), .A4(new_n364), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n313), .B(KEYINPUT8), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n291), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n315), .A2(new_n319), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g0169(.A(new_n369), .B(KEYINPUT74), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G58), .A2(G68), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n371), .B(KEYINPUT72), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n218), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n373), .A2(G20), .B1(G159), .B2(new_n293), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT71), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n253), .ZN(new_n376));
  NAND2_X1  g0176(.A1(KEYINPUT71), .A2(KEYINPUT3), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n376), .A2(G33), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(G20), .B1(new_n378), .B2(new_n252), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT7), .ZN(new_n380));
  OAI21_X1  g0180(.A(G68), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AOI211_X1 g0181(.A(KEYINPUT7), .B(G20), .C1(new_n378), .C2(new_n252), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n374), .B(KEYINPUT16), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n289), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n210), .A2(KEYINPUT7), .ZN(new_n385));
  AND2_X1   g0185(.A1(KEYINPUT71), .A2(KEYINPUT3), .ZN(new_n386));
  NOR2_X1   g0186(.A1(KEYINPUT71), .A2(KEYINPUT3), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n251), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n254), .A2(KEYINPUT73), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI211_X1 g0190(.A(KEYINPUT73), .B(new_n251), .C1(new_n386), .C2(new_n387), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n385), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n252), .A2(new_n254), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT7), .B1(new_n393), .B2(new_n210), .ZN(new_n394));
  OAI21_X1  g0194(.A(G68), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT16), .B1(new_n395), .B2(new_n374), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n370), .B1(new_n384), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G226), .A2(G1698), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(new_n326), .B2(G1698), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n378), .A2(new_n252), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G33), .A2(G87), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n262), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI22_X1  g0202(.A1(new_n269), .A2(new_n223), .B1(new_n267), .B2(new_n266), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT75), .ZN(new_n404));
  NOR4_X1   g0204(.A1(new_n402), .A2(new_n403), .A3(new_n404), .A4(G179), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n402), .A2(new_n403), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT75), .B1(new_n406), .B2(G169), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n282), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n397), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT18), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT18), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n397), .A2(new_n412), .A3(new_n409), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n406), .A2(new_n303), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(G200), .B2(new_n406), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n416), .B(new_n370), .C1(new_n396), .C2(new_n384), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT17), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n395), .A2(new_n374), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n289), .B(new_n383), .C1(new_n420), .C2(KEYINPUT16), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n421), .A2(KEYINPUT17), .A3(new_n370), .A4(new_n416), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n419), .A2(new_n422), .A3(KEYINPUT76), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT76), .B1(new_n419), .B2(new_n422), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n414), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n365), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n285), .A2(G20), .A3(new_n224), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n429), .A2(KEYINPUT25), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(KEYINPUT25), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n209), .A2(G33), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n319), .A2(new_n432), .A3(new_n216), .A4(new_n288), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n430), .B(new_n431), .C1(new_n224), .C2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT22), .ZN(new_n435));
  INV_X1    g0235(.A(G87), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n378), .A2(new_n210), .A3(new_n252), .A4(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G116), .ZN(new_n439));
  NOR3_X1   g0239(.A1(new_n251), .A2(new_n439), .A3(G20), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT23), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n210), .B2(G107), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n224), .A2(KEYINPUT23), .A3(G20), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n440), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n210), .A2(G87), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n435), .B1(new_n393), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n438), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT24), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n438), .A2(new_n444), .A3(new_n446), .A4(KEYINPUT24), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n449), .A2(new_n289), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT84), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n449), .A2(KEYINPUT84), .A3(new_n289), .A4(new_n450), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n434), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(G257), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(new_n256), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n378), .A2(new_n252), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT85), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G294), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n378), .A2(G250), .A3(new_n256), .A4(new_n252), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n378), .A2(KEYINPUT85), .A3(new_n252), .A4(new_n457), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n460), .A2(new_n461), .A3(new_n462), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n263), .ZN(new_n465));
  INV_X1    g0265(.A(G45), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(G1), .ZN(new_n467));
  AND2_X1   g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  NOR2_X1   g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n262), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(new_n225), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n467), .B(G274), .C1(new_n469), .C2(new_n468), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n465), .A2(new_n303), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n465), .A2(new_n473), .A3(new_n474), .ZN(new_n476));
  AOI22_X1  g0276(.A1(KEYINPUT86), .A2(new_n475), .B1(new_n476), .B2(new_n301), .ZN(new_n477));
  INV_X1    g0277(.A(new_n474), .ZN(new_n478));
  AOI211_X1 g0278(.A(new_n472), .B(new_n478), .C1(new_n464), .C2(new_n263), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT86), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n479), .A2(new_n480), .A3(G200), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n455), .B1(new_n477), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT87), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI211_X1 g0284(.A(KEYINPUT87), .B(new_n455), .C1(new_n477), .C2(new_n481), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G264), .A2(G1698), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n456), .B2(G1698), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n378), .A2(new_n252), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n393), .A2(G303), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT80), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n490), .A2(KEYINPUT80), .A3(new_n491), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n494), .A2(new_n263), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n470), .A2(G270), .A3(new_n262), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n474), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT79), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT79), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n497), .A2(new_n500), .A3(new_n474), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n249), .B1(new_n496), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n433), .A2(new_n439), .ZN(new_n504));
  XNOR2_X1  g0304(.A(new_n504), .B(KEYINPUT81), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n439), .A2(G20), .ZN(new_n506));
  OR2_X1    g0306(.A1(new_n284), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G283), .ZN(new_n508));
  INV_X1    g0308(.A(G97), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n508), .B(new_n210), .C1(G33), .C2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(new_n289), .A3(new_n506), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT20), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT82), .ZN(new_n514));
  OR2_X1    g0314(.A1(new_n511), .A2(new_n512), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n513), .A2(KEYINPUT82), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n505), .B(new_n507), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n503), .A2(KEYINPUT21), .A3(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT83), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n503), .A2(new_n518), .A3(KEYINPUT83), .A4(KEYINPUT21), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n503), .A2(new_n518), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT21), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n496), .A2(new_n502), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n526), .A2(new_n282), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n524), .A2(new_n525), .B1(new_n527), .B2(new_n518), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n474), .B1(new_n471), .B2(new_n456), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n378), .A2(G244), .A3(new_n256), .A4(new_n252), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT4), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n252), .A2(new_n254), .A3(G250), .A4(G1698), .ZN(new_n534));
  AND2_X1   g0334(.A1(KEYINPUT4), .A2(G244), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n252), .A2(new_n254), .A3(new_n535), .A4(new_n256), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n534), .A2(new_n536), .A3(new_n508), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n530), .B1(new_n538), .B2(new_n263), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G179), .ZN(new_n540));
  INV_X1    g0340(.A(new_n530), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n534), .A2(new_n536), .A3(new_n508), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n542), .B1(new_n532), .B2(new_n531), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n541), .B1(new_n543), .B2(new_n262), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G169), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n293), .A2(G77), .ZN(new_n547));
  XOR2_X1   g0347(.A(new_n547), .B(KEYINPUT77), .Z(new_n548));
  NAND3_X1  g0348(.A1(new_n224), .A2(KEYINPUT6), .A3(G97), .ZN(new_n549));
  XOR2_X1   g0349(.A(G97), .B(G107), .Z(new_n550));
  OAI21_X1  g0350(.A(new_n549), .B1(new_n550), .B2(KEYINPUT6), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n548), .B1(G20), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(G107), .B1(new_n392), .B2(new_n394), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n290), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n320), .A2(new_n509), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n433), .B2(new_n509), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT78), .ZN(new_n557));
  XNOR2_X1  g0357(.A(new_n556), .B(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n546), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n552), .A2(new_n553), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n558), .B1(new_n560), .B2(new_n289), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n539), .A2(G200), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n544), .A2(G190), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(G250), .B1(new_n466), .B2(G1), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n467), .A2(G274), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n263), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n378), .A2(G238), .A3(new_n256), .A4(new_n252), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n378), .A2(G244), .A3(G1698), .A4(new_n252), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n568), .B(new_n569), .C1(new_n251), .C2(new_n439), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n567), .B1(new_n570), .B2(new_n263), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n378), .A2(new_n210), .A3(G68), .A4(new_n252), .ZN(new_n572));
  NOR2_X1   g0372(.A1(G87), .A2(G97), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n573), .A2(new_n224), .B1(new_n259), .B2(new_n210), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT19), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n259), .A2(KEYINPUT19), .A3(G20), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n572), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n578), .A2(new_n289), .B1(new_n320), .B2(new_n342), .ZN(new_n579));
  INV_X1    g0379(.A(new_n433), .ZN(new_n580));
  INV_X1    g0380(.A(new_n342), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n571), .A2(new_n282), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n570), .A2(new_n263), .ZN(new_n584));
  INV_X1    g0384(.A(new_n567), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n249), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(G200), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n571), .A2(G190), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n580), .A2(G87), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n589), .A2(new_n579), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n559), .A2(new_n564), .A3(new_n588), .A4(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n518), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n526), .A2(G190), .ZN(new_n596));
  AOI21_X1  g0396(.A(G200), .B1(new_n496), .B2(new_n502), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n479), .A2(G179), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n476), .A2(G169), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n453), .A2(new_n454), .ZN(new_n602));
  INV_X1    g0402(.A(new_n434), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n529), .A2(new_n594), .A3(new_n598), .A4(new_n605), .ZN(new_n606));
  NOR3_X1   g0406(.A1(new_n428), .A2(new_n487), .A3(new_n606), .ZN(G372));
  NAND2_X1  g0407(.A1(new_n362), .A2(new_n363), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n351), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n609), .B1(new_n306), .B2(new_n305), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(new_n299), .B2(new_n283), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n423), .A2(new_n424), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n414), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n336), .A2(new_n337), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n613), .A2(new_n614), .B1(new_n322), .B2(new_n339), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n523), .A2(new_n605), .A3(new_n528), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n476), .A2(KEYINPUT86), .A3(new_n301), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n480), .B1(new_n479), .B2(new_n303), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n479), .A2(G200), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT87), .B1(new_n620), .B2(new_n455), .ZN(new_n621));
  INV_X1    g0421(.A(new_n485), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n594), .B(new_n616), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n592), .A2(new_n588), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT26), .B1(new_n624), .B2(new_n559), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n561), .B1(new_n540), .B2(new_n545), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT26), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n626), .A2(new_n627), .A3(new_n588), .A4(new_n592), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n625), .A2(new_n588), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n615), .B1(new_n428), .B2(new_n631), .ZN(G369));
  INV_X1    g0432(.A(new_n605), .ZN(new_n633));
  OR3_X1    g0433(.A1(new_n284), .A2(KEYINPUT27), .A3(G20), .ZN(new_n634));
  OAI21_X1  g0434(.A(KEYINPUT27), .B1(new_n284), .B2(G20), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(G213), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(G343), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n633), .A2(new_n639), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n484), .A2(new_n485), .B1(new_n604), .B2(new_n638), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n640), .B1(new_n641), .B2(new_n633), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n523), .A2(new_n528), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n639), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n523), .A2(new_n528), .A3(new_n598), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n518), .A2(new_n638), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n648), .B1(new_n643), .B2(new_n647), .ZN(new_n649));
  INV_X1    g0449(.A(G330), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n645), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n641), .A2(new_n643), .A3(new_n605), .A4(new_n639), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n640), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n652), .A2(new_n654), .ZN(G399));
  INV_X1    g0455(.A(new_n213), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n656), .A2(G41), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(new_n209), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n573), .A2(new_n224), .A3(new_n439), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n658), .A2(new_n660), .B1(new_n220), .B2(new_n657), .ZN(new_n661));
  XOR2_X1   g0461(.A(new_n661), .B(KEYINPUT28), .Z(new_n662));
  INV_X1    g0462(.A(KEYINPUT88), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n472), .B1(new_n464), .B2(new_n263), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n663), .B1(new_n664), .B2(new_n571), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n539), .A2(new_n502), .A3(G179), .A4(new_n496), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n664), .A2(new_n663), .A3(new_n571), .ZN(new_n668));
  AOI21_X1  g0468(.A(KEYINPUT30), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n526), .A2(new_n544), .A3(new_n586), .A4(new_n282), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(new_n479), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT89), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n668), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n673), .A2(new_n665), .A3(new_n666), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(KEYINPUT30), .ZN(new_n675));
  INV_X1    g0475(.A(new_n671), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT89), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n676), .B(new_n677), .C1(new_n674), .C2(KEYINPUT30), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n672), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT31), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n639), .A2(new_n680), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n679), .A2(KEYINPUT90), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(KEYINPUT90), .B1(new_n679), .B2(new_n681), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(KEYINPUT31), .B1(new_n606), .B2(new_n487), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n664), .A2(new_n571), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT88), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n687), .A2(new_n527), .A3(new_n539), .A4(new_n668), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT30), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n671), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n675), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n638), .B1(new_n691), .B2(KEYINPUT31), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n685), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n650), .B1(new_n684), .B2(new_n693), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n559), .A2(new_n564), .A3(new_n592), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n616), .B(new_n695), .C1(new_n621), .C2(new_n622), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n638), .B1(new_n696), .B2(new_n629), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT29), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n631), .A2(new_n638), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  XNOR2_X1  g0500(.A(KEYINPUT91), .B(KEYINPUT29), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n694), .B1(new_n698), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n662), .B1(new_n703), .B2(G1), .ZN(G364));
  AND2_X1   g0504(.A1(new_n210), .A2(G13), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G45), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT92), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n658), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n210), .A2(new_n303), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n282), .A2(new_n301), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(G326), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n301), .A2(G179), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(G303), .ZN(new_n715));
  OAI22_X1  g0515(.A1(new_n711), .A2(new_n712), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n210), .A2(G190), .ZN(new_n717));
  NOR2_X1   g0517(.A1(G179), .A2(G200), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI211_X1 g0520(.A(new_n255), .B(new_n716), .C1(G329), .C2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n717), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n722), .A2(new_n282), .A3(G200), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n710), .A2(new_n717), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  XNOR2_X1  g0525(.A(KEYINPUT33), .B(G317), .ZN(new_n726));
  AOI22_X1  g0526(.A1(new_n723), .A2(G311), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n709), .A2(G179), .A3(new_n301), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n717), .A2(new_n713), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n729), .A2(G322), .B1(new_n731), .B2(G283), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n718), .A2(G190), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G20), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G294), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n721), .A2(new_n727), .A3(new_n732), .A4(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n723), .ZN(new_n737));
  OAI22_X1  g0537(.A1(new_n737), .A2(new_n206), .B1(new_n202), .B2(new_n728), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n738), .A2(KEYINPUT96), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(KEYINPUT96), .ZN(new_n740));
  INV_X1    g0540(.A(G159), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n719), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT32), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n739), .A2(new_n740), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n730), .A2(new_n224), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n745), .B1(G68), .B2(new_n725), .ZN(new_n746));
  INV_X1    g0546(.A(new_n711), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G50), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n734), .A2(G97), .ZN(new_n749));
  INV_X1    g0549(.A(new_n714), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n393), .B1(new_n750), .B2(G87), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n746), .A2(new_n748), .A3(new_n749), .A4(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n736), .B1(new_n744), .B2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n216), .B1(G20), .B2(new_n249), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n708), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n656), .A2(new_n393), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G355), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(G116), .B2(new_n213), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n244), .A2(G45), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n759), .B1(G45), .B2(new_n220), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n378), .A2(new_n252), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n213), .A2(new_n761), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n762), .B(KEYINPUT93), .Z(new_n763));
  AOI21_X1  g0563(.A(new_n758), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT94), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G13), .A2(G33), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n210), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT95), .Z(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n754), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(new_n764), .B2(new_n765), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n755), .B1(new_n766), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n769), .B(KEYINPUT97), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n772), .B1(new_n649), .B2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n708), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n651), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n649), .A2(new_n650), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(G396));
  INV_X1    g0580(.A(KEYINPUT98), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n350), .A2(new_n639), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n609), .B1(new_n361), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n364), .A2(new_n639), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n699), .A2(new_n781), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(KEYINPUT98), .B1(new_n700), .B2(new_n785), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n630), .A2(new_n639), .A3(new_n786), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n694), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n792), .A2(new_n708), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n754), .A2(new_n767), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n708), .B1(new_n206), .B2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n754), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n729), .A2(G143), .B1(new_n725), .B2(G150), .ZN(new_n798));
  INV_X1    g0598(.A(G137), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n798), .B1(new_n799), .B2(new_n711), .C1(new_n741), .C2(new_n737), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT34), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  INV_X1    g0603(.A(G132), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n714), .A2(new_n201), .B1(new_n719), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n761), .ZN(new_n806));
  INV_X1    g0606(.A(new_n734), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n806), .B1(new_n202), .B2(new_n807), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n805), .B(new_n808), .C1(G68), .C2(new_n731), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n802), .A2(new_n803), .A3(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(G311), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n714), .A2(new_n224), .B1(new_n719), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n730), .A2(new_n436), .ZN(new_n813));
  NOR3_X1   g0613(.A1(new_n812), .A2(new_n255), .A3(new_n813), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n723), .A2(G116), .B1(new_n729), .B2(G294), .ZN(new_n815));
  AOI22_X1  g0615(.A1(G303), .A2(new_n747), .B1(new_n725), .B2(G283), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n814), .A2(new_n749), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n810), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n767), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n796), .B1(new_n797), .B2(new_n818), .C1(new_n786), .C2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n794), .A2(new_n820), .ZN(G384));
  OAI211_X1 g0621(.A(G116), .B(new_n217), .C1(new_n551), .C2(KEYINPUT35), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(KEYINPUT35), .B2(new_n551), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT36), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n372), .A2(new_n220), .A3(G77), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n201), .A2(G68), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n209), .B(G13), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n636), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n397), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n410), .A2(new_n830), .A3(new_n417), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(KEYINPUT37), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(KEYINPUT100), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n831), .A2(KEYINPUT37), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT100), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n831), .A2(new_n835), .A3(KEYINPUT37), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n830), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n411), .A2(new_n413), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n419), .A2(new_n422), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT101), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI211_X1 g0643(.A(KEYINPUT101), .B(new_n838), .C1(new_n839), .C2(new_n840), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n837), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT38), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT39), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n381), .A2(new_n382), .ZN(new_n849));
  AOI21_X1  g0649(.A(KEYINPUT16), .B1(new_n849), .B2(new_n374), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n370), .B1(new_n850), .B2(new_n384), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n829), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n425), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n851), .A2(new_n409), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n855), .A2(new_n852), .A3(new_n417), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(KEYINPUT37), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n834), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n854), .A2(KEYINPUT38), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n847), .A2(new_n848), .A3(new_n859), .ZN(new_n860));
  AOI221_X4 g0660(.A(new_n846), .B1(new_n834), .B2(new_n857), .C1(new_n425), .C2(new_n853), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT38), .B1(new_n854), .B2(new_n858), .ZN(new_n862));
  OAI21_X1  g0662(.A(KEYINPUT39), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT99), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n283), .B2(new_n299), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n275), .A2(new_n277), .B1(new_n280), .B2(new_n282), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n276), .B1(new_n280), .B2(new_n250), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n865), .B(new_n299), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n871), .A2(new_n638), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n864), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n306), .A2(new_n639), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(new_n305), .B2(new_n306), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n310), .A2(new_n874), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n638), .B(new_n785), .C1(new_n623), .C2(new_n629), .ZN(new_n879));
  INV_X1    g0679(.A(new_n784), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n861), .A2(new_n862), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n414), .A2(new_n829), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n873), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n702), .A2(new_n427), .A3(new_n698), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n615), .ZN(new_n889));
  XOR2_X1   g0689(.A(new_n887), .B(new_n889), .Z(new_n890));
  INV_X1    g0690(.A(KEYINPUT40), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n691), .A2(new_n681), .ZN(new_n892));
  NOR3_X1   g0692(.A1(new_n646), .A2(new_n593), .A3(new_n633), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n680), .B1(new_n893), .B2(new_n486), .ZN(new_n894));
  INV_X1    g0694(.A(new_n692), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(new_n786), .A3(new_n878), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n891), .B1(new_n897), .B2(new_n882), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n785), .B1(new_n693), .B2(new_n892), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n847), .A2(new_n859), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n899), .A2(new_n900), .A3(KEYINPUT40), .A4(new_n878), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n427), .A2(new_n896), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n902), .B(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n904), .A2(new_n650), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n890), .A2(new_n905), .B1(new_n209), .B2(new_n705), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n890), .A2(new_n905), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n828), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n908), .B(KEYINPUT102), .Z(G367));
  INV_X1    g0709(.A(new_n652), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n559), .B(new_n564), .C1(new_n561), .C2(new_n639), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n559), .B2(new_n639), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  OR3_X1    g0714(.A1(new_n653), .A2(KEYINPUT42), .A3(new_n913), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT42), .B1(new_n653), .B2(new_n913), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n559), .B1(new_n911), .B2(new_n605), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n639), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n579), .A2(new_n591), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n638), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(new_n587), .B2(new_n583), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n624), .B2(new_n920), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT103), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n923), .A2(KEYINPUT43), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n915), .A2(new_n916), .A3(new_n918), .A4(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT105), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n924), .B1(KEYINPUT43), .B2(new_n922), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n927), .B1(new_n926), .B2(new_n928), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n925), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n931), .A2(KEYINPUT104), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(KEYINPUT104), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n914), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n932), .A2(new_n914), .A3(new_n933), .ZN(new_n936));
  XNOR2_X1  g0736(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n657), .B(new_n937), .Z(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n654), .A2(new_n913), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n940), .B(KEYINPUT45), .Z(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n654), .A2(new_n913), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT44), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n942), .A2(new_n910), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n652), .B1(new_n941), .B2(new_n944), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n645), .A2(new_n651), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n652), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n653), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n950), .A2(KEYINPUT107), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n949), .B(new_n951), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n946), .A2(new_n703), .A3(new_n947), .A4(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n939), .B1(new_n953), .B2(new_n703), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n707), .A2(G1), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n935), .B(new_n936), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n763), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n957), .A2(new_n240), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n770), .B1(new_n213), .B2(new_n342), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n776), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n730), .A2(new_n509), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(G317), .B2(new_n720), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n962), .B(new_n761), .C1(new_n224), .C2(new_n807), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n714), .A2(new_n439), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT46), .ZN(new_n965));
  INV_X1    g0765(.A(G283), .ZN(new_n966));
  INV_X1    g0766(.A(G294), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n737), .A2(new_n966), .B1(new_n967), .B2(new_n724), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n728), .A2(new_n715), .B1(new_n711), .B2(new_n811), .ZN(new_n969));
  NOR4_X1   g0769(.A1(new_n963), .A2(new_n965), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n734), .A2(G68), .ZN(new_n971));
  INV_X1    g0771(.A(G143), .ZN(new_n972));
  INV_X1    g0772(.A(G150), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n971), .B1(new_n972), .B2(new_n711), .C1(new_n973), .C2(new_n728), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT108), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n730), .A2(new_n206), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n714), .A2(new_n202), .B1(new_n719), .B2(new_n799), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n977), .B(new_n978), .C1(G50), .C2(new_n723), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n974), .A2(new_n975), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n393), .B1(new_n725), .B2(G159), .ZN(new_n981));
  AND3_X1   g0781(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n970), .B1(new_n976), .B2(new_n982), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n983), .A2(KEYINPUT47), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n797), .B1(new_n983), .B2(KEYINPUT47), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n960), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n773), .B2(new_n922), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n956), .A2(new_n987), .ZN(G387));
  NOR2_X1   g0788(.A1(new_n714), .A2(new_n206), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n728), .A2(new_n201), .B1(new_n719), .B2(new_n973), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n989), .B(new_n990), .C1(G68), .C2(new_n723), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n761), .B(new_n961), .C1(G159), .C2(new_n747), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n366), .A2(new_n725), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n581), .A2(new_n734), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n991), .A2(new_n992), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  AOI22_X1  g0795(.A1(G322), .A2(new_n747), .B1(new_n725), .B2(G311), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT110), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n723), .A2(G303), .B1(new_n729), .B2(G317), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n1000), .A2(KEYINPUT48), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n750), .A2(G294), .B1(new_n734), .B2(G283), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n1000), .B2(KEYINPUT48), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1001), .A2(KEYINPUT49), .A3(new_n1004), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(G116), .A2(new_n731), .B1(new_n720), .B2(G326), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1005), .A2(new_n761), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(KEYINPUT49), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n995), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n754), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n345), .A2(new_n201), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT50), .Z(new_n1012));
  AOI21_X1  g0812(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1012), .A2(new_n660), .A3(new_n1013), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1014), .B(new_n763), .C1(new_n466), .C2(new_n236), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n756), .A2(new_n659), .B1(new_n224), .B2(new_n656), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1017), .A2(KEYINPUT109), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(KEYINPUT109), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n770), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1010), .B(new_n776), .C1(new_n1018), .C2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n642), .B2(new_n774), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n952), .B2(new_n955), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n952), .A2(new_n703), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n657), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n952), .A2(new_n703), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1023), .B1(new_n1025), .B2(new_n1026), .ZN(G393));
  INV_X1    g0827(.A(new_n947), .ZN(new_n1028));
  NOR3_X1   g0828(.A1(new_n941), .A2(new_n652), .A3(new_n944), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1024), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1030), .A2(new_n953), .A3(new_n657), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT111), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1030), .A2(new_n953), .A3(KEYINPUT111), .A4(new_n657), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n729), .A2(G311), .B1(new_n747), .B2(G317), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT52), .Z(new_n1036));
  AOI22_X1  g0836(.A1(G303), .A2(new_n725), .B1(new_n720), .B2(G322), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n723), .A2(G294), .B1(new_n750), .B2(G283), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n255), .B(new_n745), .C1(G116), .C2(new_n734), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n714), .A2(new_n203), .B1(new_n719), .B2(new_n972), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n813), .B(new_n1041), .C1(G50), .C2(new_n725), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n728), .A2(new_n741), .B1(new_n711), .B2(new_n973), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT51), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n345), .A2(new_n723), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n761), .B1(G77), .B2(new_n734), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1042), .A2(new_n1044), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n797), .B1(new_n1040), .B2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n957), .A2(new_n247), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n770), .B1(new_n509), .B2(new_n213), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n776), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n1048), .B(new_n1051), .C1(new_n913), .C2(new_n769), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1052), .B1(new_n1053), .B2(new_n955), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1033), .A2(new_n1034), .A3(new_n1054), .ZN(G390));
  AOI22_X1  g0855(.A1(new_n871), .A2(new_n875), .B1(new_n310), .B2(new_n874), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n791), .B2(new_n785), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n896), .A2(G330), .A3(new_n786), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1058), .A2(new_n1056), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n880), .B2(new_n879), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n679), .A2(new_n681), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT90), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n679), .A2(KEYINPUT90), .A3(new_n681), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(new_n895), .C2(new_n894), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1067), .A2(G330), .A3(new_n786), .A4(new_n878), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(KEYINPUT114), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT114), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n694), .A2(new_n1070), .A3(new_n786), .A4(new_n878), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n696), .A2(new_n629), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1073), .A2(new_n639), .A3(new_n783), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n784), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT112), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1074), .A2(KEYINPUT112), .A3(new_n784), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1077), .A2(new_n1078), .B1(new_n1058), .B2(new_n1056), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n1072), .A2(KEYINPUT115), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(KEYINPUT115), .B1(new_n1072), .B2(new_n1079), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1062), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n888), .B(new_n615), .C1(new_n903), .C2(new_n650), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT113), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1056), .B1(new_n789), .B2(new_n784), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1086), .B1(new_n1087), .B2(new_n872), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n872), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n881), .A2(KEYINPUT113), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n864), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n900), .A2(new_n1089), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1076), .B(new_n880), .C1(new_n697), .C2(new_n783), .ZN(new_n1093));
  AOI21_X1  g0893(.A(KEYINPUT112), .B1(new_n1074), .B2(new_n784), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1092), .B1(new_n1095), .B2(new_n878), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1059), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n860), .A2(new_n863), .ZN(new_n1098));
  NOR3_X1   g0898(.A1(new_n1087), .A2(new_n1086), .A3(new_n872), .ZN(new_n1099));
  AOI21_X1  g0899(.A(KEYINPUT113), .B1(new_n881), .B2(new_n1089), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1077), .A2(new_n878), .A3(new_n1078), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1102), .A2(new_n1089), .A3(new_n900), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1101), .A2(new_n1072), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1097), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1085), .A2(new_n1105), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1097), .A2(new_n1104), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1082), .A2(new_n1107), .A3(new_n1084), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1106), .A2(new_n657), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n795), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n776), .B1(new_n366), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n864), .A2(new_n819), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n729), .A2(G132), .B1(new_n720), .B2(G125), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1113), .B(new_n255), .C1(new_n201), .C2(new_n730), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n714), .A2(new_n973), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n1115), .B(KEYINPUT53), .Z(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT54), .B(G143), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n723), .A2(new_n1118), .B1(new_n747), .B2(G128), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n799), .B2(new_n724), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n807), .A2(new_n741), .ZN(new_n1121));
  NOR4_X1   g0921(.A1(new_n1114), .A2(new_n1116), .A3(new_n1120), .A4(new_n1121), .ZN(new_n1122));
  OR2_X1    g0922(.A1(new_n1122), .A2(KEYINPUT117), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(KEYINPUT117), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n730), .A2(new_n203), .B1(new_n719), .B2(new_n967), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n255), .B(new_n1125), .C1(G87), .C2(new_n750), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n734), .A2(G77), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n723), .A2(G97), .B1(new_n747), .B2(G283), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n729), .A2(G116), .B1(new_n725), .B2(G107), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1123), .A2(new_n1124), .A3(new_n1130), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1111), .B(new_n1112), .C1(new_n754), .C2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n955), .ZN(new_n1133));
  OR3_X1    g0933(.A1(new_n1105), .A2(KEYINPUT116), .A3(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(KEYINPUT116), .B1(new_n1105), .B2(new_n1133), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1132), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1109), .A2(new_n1136), .ZN(G378));
  AOI21_X1  g0937(.A(new_n708), .B1(new_n201), .B2(new_n795), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n806), .A2(G41), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n251), .A2(new_n261), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT118), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n1139), .A2(G50), .A3(new_n1141), .ZN(new_n1142));
  XOR2_X1   g0942(.A(new_n1142), .B(KEYINPUT119), .Z(new_n1143));
  INV_X1    g0943(.A(G125), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n711), .A2(new_n1144), .B1(new_n724), .B2(new_n804), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(G150), .B2(new_n734), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n729), .A2(G128), .B1(new_n750), .B2(new_n1118), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1146), .B(new_n1147), .C1(new_n799), .C2(new_n737), .ZN(new_n1148));
  OR2_X1    g0948(.A1(new_n1148), .A2(KEYINPUT59), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n720), .A2(G124), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1150), .B(new_n1141), .C1(new_n741), .C2(new_n730), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n1148), .B2(KEYINPUT59), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1143), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n737), .A2(new_n342), .B1(new_n719), .B2(new_n966), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(G97), .B2(new_n725), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n989), .B1(G58), .B2(new_n731), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n729), .A2(G107), .B1(new_n747), .B2(G116), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1156), .A2(new_n1157), .A3(new_n971), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1155), .A2(new_n1158), .A3(new_n1139), .ZN(new_n1159));
  XOR2_X1   g0959(.A(new_n1159), .B(KEYINPUT120), .Z(new_n1160));
  OAI21_X1  g0960(.A(new_n1153), .B1(new_n1160), .B2(KEYINPUT58), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(KEYINPUT58), .B2(new_n1160), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1138), .B1(new_n1162), .B2(new_n797), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n322), .A2(new_n829), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n341), .B(new_n1165), .ZN(new_n1166));
  XOR2_X1   g0966(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1167));
  XNOR2_X1  g0967(.A(new_n1166), .B(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1163), .B1(new_n1169), .B2(new_n767), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n898), .A2(new_n901), .A3(G330), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1089), .B1(new_n860), .B2(new_n863), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1173), .A2(new_n885), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1169), .B1(new_n1174), .B2(new_n884), .ZN(new_n1175));
  NOR4_X1   g0975(.A1(new_n1173), .A2(new_n883), .A3(new_n1168), .A4(new_n885), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1172), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n887), .A2(new_n1168), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1174), .A2(new_n884), .A3(new_n1169), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1178), .A2(new_n1171), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1170), .B1(new_n1181), .B2(new_n955), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT57), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1083), .B1(new_n1082), .B2(new_n1107), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1175), .A2(new_n1176), .A3(new_n1172), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1171), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  OAI211_X1 g0987(.A(KEYINPUT121), .B(new_n1183), .C1(new_n1184), .C2(new_n1187), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1057), .A2(new_n1060), .B1(new_n784), .B2(new_n789), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1072), .A2(new_n1079), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT115), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1072), .A2(KEYINPUT115), .A3(new_n1079), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1189), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1084), .B1(new_n1194), .B2(new_n1105), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1195), .A2(KEYINPUT57), .A3(new_n1181), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1188), .A2(new_n657), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1195), .A2(new_n1181), .ZN(new_n1198));
  AOI21_X1  g0998(.A(KEYINPUT121), .B1(new_n1198), .B2(new_n1183), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1182), .B1(new_n1197), .B2(new_n1199), .ZN(G375));
  OAI22_X1  g1000(.A1(new_n728), .A2(new_n799), .B1(new_n711), .B2(new_n804), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(G159), .B2(new_n750), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n723), .A2(G150), .B1(new_n731), .B2(G58), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n725), .A2(new_n1118), .B1(new_n720), .B2(G128), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n761), .B1(G50), .B2(new_n734), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n728), .A2(new_n966), .B1(new_n724), .B2(new_n439), .ZN(new_n1207));
  NOR3_X1   g1007(.A1(new_n1207), .A2(new_n255), .A3(new_n977), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(G97), .A2(new_n750), .B1(new_n720), .B2(G303), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n723), .A2(G107), .B1(new_n747), .B2(G294), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1208), .A2(new_n994), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n797), .B1(new_n1206), .B2(new_n1211), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n708), .B(new_n1212), .C1(new_n203), .C2(new_n795), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n878), .B2(new_n819), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n1194), .B2(new_n1133), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT122), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  OAI211_X1 g1017(.A(KEYINPUT122), .B(new_n1214), .C1(new_n1194), .C2(new_n1133), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1085), .A2(new_n938), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n1194), .B2(new_n1083), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1219), .A2(new_n1221), .ZN(G381));
  OR2_X1    g1022(.A1(G375), .A2(G378), .ZN(new_n1223));
  OR2_X1    g1023(.A1(G393), .A2(G396), .ZN(new_n1224));
  OR4_X1    g1024(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1224), .ZN(new_n1225));
  OR3_X1    g1025(.A1(new_n1223), .A2(new_n1225), .A3(G381), .ZN(G407));
  OAI211_X1 g1026(.A(G407), .B(G213), .C1(G343), .C2(new_n1223), .ZN(G409));
  INV_X1    g1027(.A(KEYINPUT124), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(G387), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1229), .A2(KEYINPUT125), .A3(G390), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(G393), .B(new_n779), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(G390), .A2(new_n956), .A3(new_n987), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT125), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1231), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(G390), .A2(KEYINPUT125), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1235), .A2(G387), .A3(new_n1228), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1230), .A2(new_n1234), .A3(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1232), .ZN(new_n1238));
  AOI21_X1  g1038(.A(G390), .B1(new_n956), .B2(new_n987), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1231), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1237), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT61), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT126), .ZN(new_n1244));
  OAI211_X1 g1044(.A(G378), .B(new_n1182), .C1(new_n1197), .C2(new_n1199), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1182), .B1(new_n1198), .B2(new_n939), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1246), .A2(new_n1109), .A3(new_n1136), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(G213), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1249), .A2(G343), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1244), .B1(new_n1248), .B2(new_n1251), .ZN(new_n1252));
  AOI211_X1 g1052(.A(KEYINPUT126), .B(new_n1250), .C1(new_n1245), .C2(new_n1247), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT60), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT60), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1194), .A2(new_n1256), .A3(new_n1083), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1085), .A2(new_n657), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1258), .A2(new_n1260), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1261));
  OAI21_X1  g1061(.A(KEYINPUT123), .B1(new_n1261), .B2(G384), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT123), .ZN(new_n1263));
  INV_X1    g1063(.A(G384), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1259), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1263), .B(new_n1264), .C1(new_n1219), .C2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1261), .A2(G384), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1262), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1250), .A2(G2897), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1262), .A2(new_n1266), .A3(new_n1267), .A4(new_n1269), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1243), .B1(new_n1254), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1268), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1250), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT62), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  AND2_X1   g1077(.A1(new_n1275), .A2(KEYINPUT62), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1277), .B1(new_n1254), .B2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1242), .B1(new_n1274), .B2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(KEYINPUT63), .B1(new_n1273), .B2(new_n1276), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1241), .A2(new_n1243), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1275), .A2(KEYINPUT63), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1284), .B1(new_n1254), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1283), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1280), .A2(new_n1287), .ZN(G405));
  INV_X1    g1088(.A(KEYINPUT127), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(G375), .A2(G378), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1223), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n1275), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1223), .A2(new_n1268), .A3(new_n1290), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1289), .B1(new_n1294), .B2(new_n1242), .ZN(new_n1295));
  AOI211_X1 g1095(.A(KEYINPUT127), .B(new_n1241), .C1(new_n1292), .C2(new_n1293), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1294), .A2(new_n1242), .ZN(new_n1297));
  NOR3_X1   g1097(.A1(new_n1295), .A2(new_n1296), .A3(new_n1297), .ZN(G402));
endmodule


