//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1285,
    new_n1286, new_n1287, new_n1288, new_n1289, new_n1290, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  AND2_X1   g0004(.A1(KEYINPUT64), .A2(G68), .ZN(new_n205));
  NOR2_X1   g0005(.A1(KEYINPUT64), .A2(G68), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AOI22_X1  g0007(.A1(new_n207), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G50), .A2(G226), .ZN(new_n209));
  INV_X1    g0009(.A(G244), .ZN(new_n210));
  XNOR2_X1  g0010(.A(KEYINPUT65), .B(G77), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n208), .B(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(KEYINPUT66), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G87), .B2(G250), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n212), .A2(KEYINPUT66), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n214), .B(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n218), .B1(G97), .B2(G257), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G107), .A2(G264), .ZN(new_n220));
  AOI22_X1  g0020(.A1(new_n219), .A2(new_n220), .B1(G1), .B2(G20), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT1), .Z(new_n222));
  INV_X1    g0022(.A(G1), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR3_X1   g0024(.A1(new_n223), .A2(new_n224), .A3(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT0), .Z(new_n227));
  NOR2_X1   g0027(.A1(G58), .A2(G68), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n230), .A2(new_n224), .A3(new_n231), .ZN(new_n232));
  NOR3_X1   g0032(.A1(new_n222), .A2(new_n227), .A3(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  INV_X1    g0038(.A(G264), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XOR2_X1   g0043(.A(G50), .B(G58), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  XNOR2_X1  g0049(.A(KEYINPUT3), .B(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G223), .A2(G1698), .ZN(new_n251));
  INV_X1    g0051(.A(G222), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n251), .B1(new_n252), .B2(G1698), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(new_n211), .B2(new_n250), .ZN(new_n255));
  OR2_X1    g0055(.A1(new_n255), .A2(KEYINPUT68), .ZN(new_n256));
  AND2_X1   g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  OAI21_X1  g0057(.A(KEYINPUT69), .B1(new_n257), .B2(new_n231), .ZN(new_n258));
  AND2_X1   g0058(.A1(G1), .A2(G13), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT69), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n255), .A2(KEYINPUT68), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n256), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n223), .B(G274), .C1(G41), .C2(G45), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT67), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n267), .B(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G41), .ZN(new_n270));
  INV_X1    g0070(.A(G45), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n223), .A2(new_n272), .B1(new_n259), .B2(new_n261), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n269), .B1(G226), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n266), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n275), .A2(G179), .ZN(new_n276));
  INV_X1    g0076(.A(G169), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n276), .B1(new_n277), .B2(new_n275), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n231), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n224), .A2(G33), .ZN(new_n281));
  OR2_X1    g0081(.A1(KEYINPUT8), .A2(G58), .ZN(new_n282));
  NAND2_X1  g0082(.A1(KEYINPUT8), .A2(G58), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT70), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT70), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n282), .A2(new_n286), .A3(new_n283), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n281), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(G20), .B1(new_n229), .B2(G50), .ZN(new_n289));
  INV_X1    g0089(.A(G150), .ZN(new_n290));
  INV_X1    g0090(.A(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n224), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n289), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n280), .B1(new_n288), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n280), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n223), .A2(G20), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G50), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n223), .A2(G13), .A3(G20), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n294), .B(new_n299), .C1(G50), .C2(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n278), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT9), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n275), .A2(G200), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G190), .ZN(new_n305));
  OAI221_X1 g0105(.A(new_n304), .B1(new_n303), .B2(new_n301), .C1(new_n305), .C2(new_n275), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n306), .A2(KEYINPUT10), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(KEYINPUT10), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n302), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n269), .B1(G238), .B2(new_n273), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT13), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n217), .A2(G1698), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(G226), .B2(G1698), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT3), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G33), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n291), .A2(KEYINPUT3), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G97), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n313), .A2(new_n317), .B1(new_n291), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n264), .A2(new_n319), .ZN(new_n320));
  AND3_X1   g0120(.A1(new_n310), .A2(new_n311), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n311), .B1(new_n310), .B2(new_n320), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G200), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT12), .ZN(new_n326));
  NOR3_X1   g0126(.A1(new_n207), .A2(new_n326), .A3(new_n300), .ZN(new_n327));
  INV_X1    g0127(.A(G68), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n328), .B1(new_n297), .B2(KEYINPUT12), .ZN(new_n329));
  AOI211_X1 g0129(.A(new_n327), .B(new_n329), .C1(new_n326), .C2(new_n300), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n207), .A2(new_n224), .ZN(new_n331));
  INV_X1    g0131(.A(G50), .ZN(new_n332));
  INV_X1    g0132(.A(G77), .ZN(new_n333));
  OAI22_X1  g0133(.A1(new_n292), .A2(new_n332), .B1(new_n281), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n280), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g0135(.A(new_n335), .B(KEYINPUT11), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n330), .A2(new_n336), .ZN(new_n337));
  NOR3_X1   g0137(.A1(new_n321), .A2(new_n322), .A3(new_n305), .ZN(new_n338));
  NOR3_X1   g0138(.A1(new_n325), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT72), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n323), .A2(G179), .B1(new_n340), .B2(KEYINPUT14), .ZN(new_n341));
  OAI22_X1  g0141(.A1(new_n323), .A2(new_n277), .B1(new_n340), .B2(KEYINPUT14), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n340), .A2(KEYINPUT14), .ZN(new_n343));
  OAI211_X1 g0143(.A(G169), .B(new_n343), .C1(new_n321), .C2(new_n322), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n341), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n339), .B1(new_n345), .B2(new_n337), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n269), .B1(G244), .B2(new_n273), .ZN(new_n347));
  NAND2_X1  g0147(.A1(G238), .A2(G1698), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n250), .B(new_n348), .C1(new_n217), .C2(G1698), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n264), .B(new_n349), .C1(G107), .C2(new_n250), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT71), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT71), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n347), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G190), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n352), .A2(G200), .A3(new_n354), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n284), .A2(new_n292), .B1(new_n211), .B2(new_n224), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT15), .B(G87), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(new_n281), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n280), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n298), .A2(G77), .ZN(new_n362));
  INV_X1    g0162(.A(new_n300), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n211), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n361), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n356), .A2(new_n357), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n309), .A2(new_n346), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G116), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n223), .A2(new_n369), .A3(G13), .A4(G20), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n223), .A2(G33), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n295), .A2(G116), .A3(new_n371), .A4(new_n300), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n279), .A2(new_n231), .B1(G20), .B2(new_n369), .ZN(new_n373));
  NAND2_X1  g0173(.A1(G33), .A2(G283), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n374), .B(new_n224), .C1(G33), .C2(new_n318), .ZN(new_n375));
  AND3_X1   g0175(.A1(new_n373), .A2(KEYINPUT20), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(KEYINPUT20), .B1(new_n373), .B2(new_n375), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n370), .B(new_n372), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT80), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n373), .A2(new_n375), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT20), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n373), .A2(KEYINPUT20), .A3(new_n375), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n385), .A2(KEYINPUT80), .A3(new_n370), .A4(new_n372), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT73), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n291), .B2(KEYINPUT3), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n314), .A2(KEYINPUT73), .A3(G33), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(G257), .ZN(new_n392));
  INV_X1    g0192(.A(G1698), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n239), .A2(G1698), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n391), .A2(new_n316), .A3(new_n394), .A4(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n317), .A2(G303), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n264), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT77), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n270), .A2(KEYINPUT5), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n223), .A2(G45), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n270), .A2(KEYINPUT5), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT5), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(G41), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n406), .A2(KEYINPUT77), .A3(new_n223), .A4(G45), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n403), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n259), .A2(new_n261), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(G270), .A3(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(G274), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(new_n259), .B2(new_n261), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n403), .A2(new_n407), .A3(new_n412), .A4(new_n404), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n413), .A2(KEYINPUT78), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n413), .A2(KEYINPUT78), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n399), .B(new_n410), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n387), .A2(G169), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT21), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g0219(.A(new_n413), .B(KEYINPUT78), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n399), .A2(new_n410), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n387), .A2(G179), .A3(new_n420), .A4(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n387), .A2(KEYINPUT21), .A3(new_n416), .A4(G169), .ZN(new_n423));
  AND3_X1   g0223(.A1(new_n419), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n416), .A2(G200), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n380), .A2(new_n386), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n420), .A2(G190), .A3(new_n410), .A4(new_n399), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT81), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n425), .A2(new_n426), .A3(KEYINPUT81), .A4(new_n427), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n424), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g0233(.A(KEYINPUT84), .B(KEYINPUT25), .C1(new_n300), .C2(G107), .ZN(new_n434));
  INV_X1    g0234(.A(G107), .ZN(new_n435));
  NAND2_X1  g0235(.A1(KEYINPUT84), .A2(KEYINPUT25), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n363), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(KEYINPUT84), .A2(KEYINPUT25), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n295), .A2(new_n371), .A3(new_n300), .ZN(new_n439));
  OAI221_X1 g0239(.A(new_n434), .B1(new_n437), .B2(new_n438), .C1(new_n439), .C2(new_n435), .ZN(new_n440));
  XNOR2_X1  g0240(.A(KEYINPUT82), .B(KEYINPUT24), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G87), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(G20), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n444), .A2(new_n315), .A3(new_n316), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT22), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT23), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(new_n224), .B2(G107), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n435), .A2(KEYINPUT23), .A3(G20), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G116), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(G20), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n447), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n314), .A2(G33), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n456), .B1(new_n389), .B2(new_n390), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n457), .A2(KEYINPUT22), .A3(new_n444), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n442), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n453), .B1(new_n445), .B2(new_n446), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n458), .A2(new_n460), .A3(new_n442), .A4(new_n451), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n280), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT83), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n458), .A2(new_n460), .A3(new_n451), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n441), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n461), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(KEYINPUT83), .A3(new_n280), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n440), .B1(new_n465), .B2(new_n469), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n314), .A2(KEYINPUT73), .A3(G33), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT73), .B1(new_n314), .B2(G33), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n316), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(G250), .ZN(new_n474));
  MUX2_X1   g0274(.A(new_n474), .B(new_n392), .S(G1698), .Z(new_n475));
  INV_X1    g0275(.A(G294), .ZN(new_n476));
  OAI22_X1  g0276(.A1(new_n473), .A2(new_n475), .B1(new_n291), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n264), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n408), .A2(G264), .A3(new_n409), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n480), .A2(KEYINPUT85), .A3(new_n305), .A4(new_n420), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT85), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n478), .B(new_n479), .C1(new_n414), .C2(new_n415), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n482), .B1(new_n483), .B2(new_n324), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n483), .A2(G190), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n481), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n470), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n408), .A2(G257), .A3(new_n409), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n414), .B2(new_n415), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n391), .A2(G244), .A3(new_n393), .A4(new_n316), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n393), .A2(KEYINPUT4), .A3(G244), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n493), .B1(new_n474), .B2(new_n393), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n494), .A2(new_n250), .B1(G33), .B2(G283), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n263), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(G200), .B1(new_n489), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT6), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n498), .A2(new_n318), .A3(G107), .ZN(new_n499));
  XNOR2_X1  g0299(.A(G97), .B(G107), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n499), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  OAI22_X1  g0301(.A1(new_n501), .A2(new_n224), .B1(new_n333), .B2(new_n292), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT7), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n503), .B1(new_n250), .B2(G20), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n317), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n435), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n280), .B1(new_n502), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n439), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G97), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n363), .A2(new_n318), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n507), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n492), .A2(new_n495), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n264), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n513), .A2(new_n420), .A3(G190), .A4(new_n488), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n497), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n277), .B1(new_n489), .B2(new_n496), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n507), .A2(new_n509), .A3(new_n510), .ZN(new_n517));
  INV_X1    g0317(.A(G179), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n513), .A2(new_n420), .A3(new_n518), .A4(new_n488), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n440), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT83), .B1(new_n468), .B2(new_n280), .ZN(new_n523));
  AOI211_X1 g0323(.A(new_n464), .B(new_n295), .C1(new_n467), .C2(new_n461), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n480), .A2(new_n518), .A3(new_n420), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n483), .A2(new_n277), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n359), .A2(new_n363), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n457), .A2(new_n224), .A3(G68), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT19), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n533), .A2(new_n291), .A3(new_n318), .ZN(new_n534));
  OAI22_X1  g0334(.A1(new_n534), .A2(G20), .B1(G87), .B2(new_n203), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n533), .B1(new_n281), .B2(new_n318), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n532), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n531), .B1(new_n537), .B2(new_n280), .ZN(new_n538));
  XNOR2_X1  g0338(.A(new_n359), .B(KEYINPUT79), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n508), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n402), .A2(new_n474), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n223), .A2(new_n411), .A3(G45), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n542), .A2(new_n409), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n452), .ZN(new_n545));
  NOR2_X1   g0345(.A1(G238), .A2(G1698), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(new_n210), .B2(G1698), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n545), .B1(new_n457), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n544), .B1(new_n548), .B2(new_n263), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n277), .ZN(new_n550));
  INV_X1    g0350(.A(new_n544), .ZN(new_n551));
  INV_X1    g0351(.A(new_n548), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n551), .B1(new_n552), .B2(new_n264), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n518), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n541), .A2(new_n550), .A3(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n439), .A2(new_n443), .ZN(new_n556));
  AOI211_X1 g0356(.A(new_n531), .B(new_n556), .C1(new_n537), .C2(new_n280), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n549), .A2(G200), .ZN(new_n558));
  OAI211_X1 g0358(.A(G190), .B(new_n544), .C1(new_n548), .C2(new_n263), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n487), .A2(new_n521), .A3(new_n530), .A4(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n285), .A2(new_n300), .A3(new_n287), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n285), .A2(new_n287), .B1(new_n296), .B2(new_n295), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT75), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n285), .A2(new_n287), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n297), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT75), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n570), .A3(new_n564), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT16), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n228), .B1(new_n207), .B2(G58), .ZN(new_n574));
  INV_X1    g0374(.A(G159), .ZN(new_n575));
  OAI22_X1  g0375(.A1(new_n574), .A2(new_n224), .B1(new_n575), .B2(new_n292), .ZN(new_n576));
  XNOR2_X1  g0376(.A(KEYINPUT64), .B(G68), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n577), .B1(new_n504), .B2(new_n505), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n573), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT74), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT7), .B1(new_n317), .B2(new_n224), .ZN(new_n581));
  AOI211_X1 g0381(.A(new_n503), .B(G20), .C1(new_n315), .C2(new_n316), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n207), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n292), .A2(new_n575), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n229), .B1(new_n577), .B2(new_n216), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n584), .B1(new_n585), .B2(G20), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT74), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n588), .A3(new_n573), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n580), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n473), .A2(new_n503), .A3(new_n224), .ZN(new_n591));
  OAI21_X1  g0391(.A(KEYINPUT7), .B1(new_n457), .B2(G20), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n592), .A3(G68), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(KEYINPUT16), .A3(new_n586), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n594), .A2(new_n280), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n572), .B1(new_n590), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(G226), .A2(G1698), .ZN(new_n597));
  INV_X1    g0397(.A(G223), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n597), .B1(new_n598), .B2(G1698), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n391), .A2(new_n316), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(G33), .A2(G87), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n263), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(G1), .B1(new_n270), .B2(new_n271), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n603), .A2(new_n268), .A3(G274), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n267), .A2(KEYINPUT67), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n603), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n607), .A2(G232), .A3(new_n409), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n277), .B1(new_n602), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g0410(.A1(G232), .A2(new_n273), .B1(new_n604), .B2(new_n605), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n457), .A2(new_n599), .B1(G33), .B2(G87), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n611), .B(new_n518), .C1(new_n612), .C2(new_n263), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT76), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT76), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n610), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(KEYINPUT18), .B1(new_n596), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n617), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n616), .B1(new_n610), .B2(new_n613), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT18), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n594), .A2(new_n280), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n624), .B1(new_n580), .B2(new_n589), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n622), .B(new_n623), .C1(new_n625), .C2(new_n572), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n619), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT17), .ZN(new_n629));
  OAI21_X1  g0429(.A(G200), .B1(new_n602), .B2(new_n609), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n611), .B(G190), .C1(new_n612), .C2(new_n263), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n630), .A2(new_n567), .A3(new_n631), .A4(new_n571), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n629), .B1(new_n625), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n588), .B1(new_n587), .B2(new_n573), .ZN(new_n634));
  AOI211_X1 g0434(.A(KEYINPUT74), .B(KEYINPUT16), .C1(new_n583), .C2(new_n586), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n280), .B(new_n594), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n632), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(KEYINPUT17), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n355), .A2(new_n518), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n352), .A2(new_n277), .A3(new_n354), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n365), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n628), .A2(new_n640), .A3(new_n644), .ZN(new_n645));
  NOR4_X1   g0445(.A1(new_n368), .A2(new_n433), .A3(new_n563), .A4(new_n645), .ZN(G372));
  NOR2_X1   g0446(.A1(new_n368), .A2(new_n645), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n558), .A2(KEYINPUT86), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT86), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n549), .A2(new_n649), .A3(G200), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n648), .A2(new_n557), .A3(new_n559), .A4(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n555), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n652), .B1(new_n470), .B2(new_n486), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n419), .A2(new_n422), .A3(new_n423), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n465), .A2(new_n469), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n528), .B1(new_n655), .B2(new_n522), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n653), .B(new_n521), .C1(new_n654), .C2(new_n656), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n549), .A2(new_n649), .A3(G200), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n649), .B1(new_n549), .B2(G200), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n556), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n538), .A2(new_n559), .A3(new_n661), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n538), .A2(new_n540), .B1(new_n553), .B2(new_n518), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n660), .A2(new_n662), .B1(new_n663), .B2(new_n550), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT26), .B1(new_n561), .B2(new_n520), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n667), .A2(new_n555), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n657), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n647), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT87), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n345), .A2(new_n337), .ZN(new_n673));
  AOI211_X1 g0473(.A(new_n339), .B(new_n639), .C1(new_n673), .C2(new_n644), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n672), .B1(new_n674), .B2(new_n627), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n339), .B1(new_n673), .B2(new_n644), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n640), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n677), .A2(KEYINPUT87), .A3(new_n628), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n307), .A2(new_n308), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n302), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n680), .A2(KEYINPUT88), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(KEYINPUT88), .B1(new_n680), .B2(new_n681), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n671), .B1(new_n682), .B2(new_n683), .ZN(G369));
  NAND3_X1  g0484(.A1(new_n223), .A2(new_n224), .A3(G13), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(KEYINPUT27), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G213), .A3(new_n687), .ZN(new_n688));
  XOR2_X1   g0488(.A(KEYINPUT89), .B(G343), .Z(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n487), .B1(new_n470), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n530), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n656), .A2(new_n692), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(G330), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n654), .B1(new_n430), .B2(new_n431), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n426), .B2(new_n692), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n654), .A2(new_n387), .A3(new_n691), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n697), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n701), .A2(KEYINPUT90), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(KEYINPUT90), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n696), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n654), .A2(new_n692), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n696), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(new_n695), .A3(new_n707), .ZN(G399));
  INV_X1    g0508(.A(new_n225), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(G1), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n230), .B2(new_n711), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT28), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT92), .ZN(new_n716));
  AOI21_X1  g0516(.A(G179), .B1(new_n421), .B2(new_n420), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n513), .A2(new_n420), .A3(new_n488), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n717), .A2(new_n549), .A3(new_n483), .A4(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n478), .A2(new_n479), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n416), .A2(new_n518), .A3(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n513), .A2(new_n420), .A3(new_n553), .A4(new_n488), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n720), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n421), .A2(new_n480), .A3(G179), .A4(new_n420), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n726), .A2(KEYINPUT30), .A3(new_n723), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n719), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT91), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n692), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI211_X1 g0530(.A(KEYINPUT91), .B(new_n719), .C1(new_n725), .C2(new_n727), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n563), .A2(new_n433), .A3(new_n691), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT31), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n728), .A2(KEYINPUT31), .A3(new_n691), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n716), .B1(new_n737), .B2(G330), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n515), .A2(new_n520), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n656), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n561), .B1(new_n470), .B2(new_n486), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n698), .A2(new_n740), .A3(new_n741), .A4(new_n692), .ZN(new_n742));
  AOI22_X1  g0542(.A1(new_n742), .A2(KEYINPUT31), .B1(new_n731), .B2(new_n730), .ZN(new_n743));
  INV_X1    g0543(.A(new_n736), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n716), .B(G330), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n738), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n670), .A2(new_n692), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(KEYINPUT29), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT29), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n562), .A2(new_n665), .A3(new_n666), .ZN(new_n751));
  OAI21_X1  g0551(.A(KEYINPUT26), .B1(new_n652), .B2(new_n520), .ZN(new_n752));
  AND3_X1   g0552(.A1(new_n751), .A2(new_n752), .A3(new_n555), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT93), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n739), .B(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n653), .B1(new_n654), .B2(new_n656), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n753), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n750), .B1(new_n757), .B2(new_n692), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n749), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n747), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n715), .B1(new_n761), .B2(G1), .ZN(G364));
  NOR2_X1   g0562(.A1(new_n702), .A2(new_n703), .ZN(new_n763));
  INV_X1    g0563(.A(G13), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G20), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G45), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n711), .A2(G1), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n699), .A2(new_n700), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n763), .B(new_n767), .C1(G330), .C2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n231), .B1(G20), .B2(new_n277), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n224), .A2(G179), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n771), .A2(G190), .A3(G200), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n772), .A2(KEYINPUT97), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(KEYINPUT97), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n771), .A2(new_n305), .A3(G200), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n776), .A2(G87), .B1(G107), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n224), .A2(new_n518), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT96), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(KEYINPUT96), .B1(new_n224), .B2(new_n518), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n305), .A2(G200), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G190), .A2(G200), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n782), .A2(new_n783), .A3(new_n786), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n779), .B1(new_n216), .B2(new_n785), .C1(new_n211), .C2(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n780), .A2(G190), .A3(G200), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n332), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n771), .A2(new_n786), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G159), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT32), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n780), .A2(new_n305), .A3(G200), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n784), .A2(new_n518), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G20), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n250), .B1(new_n328), .B2(new_n795), .C1(new_n798), .C2(new_n318), .ZN(new_n799));
  NOR4_X1   g0599(.A1(new_n788), .A2(new_n790), .A3(new_n794), .A4(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n789), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n801), .A2(G326), .B1(new_n792), .B2(G329), .ZN(new_n802));
  INV_X1    g0602(.A(G322), .ZN(new_n803));
  INV_X1    g0603(.A(G303), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n802), .B1(new_n803), .B2(new_n785), .C1(new_n775), .C2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G311), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n787), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G283), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n777), .A2(new_n808), .ZN(new_n809));
  XOR2_X1   g0609(.A(KEYINPUT33), .B(G317), .Z(new_n810));
  OAI221_X1 g0610(.A(new_n317), .B1(new_n795), .B2(new_n810), .C1(new_n798), .C2(new_n476), .ZN(new_n811));
  NOR4_X1   g0611(.A1(new_n805), .A2(new_n807), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n770), .B1(new_n800), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n767), .ZN(new_n814));
  AND3_X1   g0614(.A1(G355), .A2(new_n225), .A3(new_n250), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n225), .A2(G116), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n457), .A2(new_n709), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n230), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n818), .B1(new_n271), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n245), .A2(G45), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n815), .B(new_n816), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(G13), .A2(G33), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(G20), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(new_n770), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT94), .Z(new_n827));
  OAI21_X1  g0627(.A(new_n814), .B1(new_n822), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT95), .ZN(new_n829));
  INV_X1    g0629(.A(new_n825), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n813), .B(new_n829), .C1(new_n768), .C2(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n769), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G396));
  NAND2_X1  g0633(.A1(new_n365), .A2(new_n691), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT98), .Z(new_n835));
  NAND2_X1  g0635(.A1(new_n367), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n644), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n643), .A2(new_n365), .A3(new_n692), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n747), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n839), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n738), .B2(new_n746), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n748), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n840), .A2(new_n670), .A3(new_n692), .A4(new_n842), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n844), .A2(new_n767), .A3(new_n845), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n798), .A2(new_n318), .B1(new_n806), .B2(new_n791), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n317), .B1(new_n785), .B2(new_n476), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n787), .A2(new_n369), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n795), .A2(new_n808), .B1(new_n777), .B2(new_n443), .ZN(new_n850));
  NOR4_X1   g0650(.A1(new_n847), .A2(new_n848), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n851), .B1(new_n435), .B2(new_n775), .C1(new_n804), .C2(new_n789), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n798), .A2(new_n216), .ZN(new_n853));
  INV_X1    g0653(.A(new_n785), .ZN(new_n854));
  INV_X1    g0654(.A(new_n795), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n854), .A2(G143), .B1(G150), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(G137), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n856), .B1(new_n857), .B2(new_n789), .C1(new_n575), .C2(new_n787), .ZN(new_n858));
  XOR2_X1   g0658(.A(new_n858), .B(KEYINPUT34), .Z(new_n859));
  AOI211_X1 g0659(.A(new_n853), .B(new_n859), .C1(G132), .C2(new_n792), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n860), .B1(new_n332), .B2(new_n775), .C1(new_n328), .C2(new_n777), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n852), .B1(new_n861), .B2(new_n473), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n770), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n770), .A2(new_n823), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n333), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n839), .A2(new_n823), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n863), .A2(new_n814), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n846), .A2(new_n867), .ZN(G384));
  NAND2_X1  g0668(.A1(new_n337), .A2(new_n691), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n346), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n345), .A2(new_n337), .A3(new_n691), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n839), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n730), .A2(KEYINPUT31), .A3(new_n731), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n872), .B1(new_n743), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n688), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT16), .B1(new_n593), .B2(new_n586), .ZN(new_n878));
  OAI22_X1  g0678(.A1(new_n624), .A2(new_n878), .B1(new_n565), .B2(new_n566), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n877), .B(new_n879), .C1(new_n627), .C2(new_n639), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n634), .A2(new_n635), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n637), .B1(new_n881), .B2(new_n624), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT37), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n877), .B1(new_n615), .B2(new_n617), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n882), .B(new_n883), .C1(new_n596), .C2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n688), .B1(new_n620), .B2(new_n621), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n879), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n883), .B1(new_n888), .B2(new_n882), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT99), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT99), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n887), .A2(new_n879), .B1(new_n636), .B2(new_n637), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n885), .B(new_n891), .C1(new_n892), .C2(new_n883), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n880), .A2(new_n890), .A3(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n880), .A2(new_n890), .A3(KEYINPUT38), .A4(new_n893), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n876), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n629), .B(new_n632), .C1(new_n590), .C2(new_n595), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT17), .B1(new_n636), .B2(new_n637), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT100), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT100), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n633), .A2(new_n904), .A3(new_n638), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n903), .A2(new_n905), .A3(new_n619), .A4(new_n626), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n596), .A2(new_n688), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n882), .B1(new_n596), .B2(new_n884), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT37), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n906), .A2(new_n907), .B1(new_n885), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n897), .B1(new_n910), .B2(KEYINPUT38), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n911), .A2(KEYINPUT40), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n899), .A2(new_n900), .B1(new_n912), .B2(new_n876), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n735), .A2(new_n873), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n913), .A2(new_n647), .A3(new_n914), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n896), .A2(new_n897), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n900), .B1(new_n916), .B2(new_n875), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n914), .A2(new_n911), .A3(KEYINPUT40), .A4(new_n872), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n917), .A2(G330), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n697), .B1(new_n735), .B2(new_n873), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n647), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n915), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT101), .ZN(new_n924));
  INV_X1    g0724(.A(new_n759), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n647), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n682), .B2(new_n683), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n924), .B(new_n927), .Z(new_n928));
  NAND2_X1  g0728(.A1(new_n870), .A2(new_n871), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n643), .A2(new_n365), .B1(new_n367), .B2(new_n835), .ZN(new_n930));
  AOI211_X1 g0730(.A(new_n691), .B(new_n930), .C1(new_n657), .C2(new_n669), .ZN(new_n931));
  INV_X1    g0731(.A(new_n838), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n934), .A2(new_n898), .B1(new_n627), .B2(new_n688), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT39), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n911), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n896), .A2(KEYINPUT39), .A3(new_n897), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n345), .A2(new_n337), .A3(new_n692), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n935), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n928), .B(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n223), .B2(new_n765), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT35), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n224), .B(new_n231), .C1(new_n501), .C2(new_n944), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n945), .B(G116), .C1(new_n944), .C2(new_n501), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT36), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n819), .B1(new_n577), .B2(new_n216), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n948), .A2(new_n211), .B1(G50), .B2(new_n328), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(G1), .A3(new_n764), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n943), .A2(new_n947), .A3(new_n950), .ZN(G367));
  NOR2_X1   g0751(.A1(new_n775), .A2(new_n369), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT46), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT109), .ZN(new_n954));
  AOI22_X1  g0754(.A1(G97), .A2(new_n778), .B1(new_n797), .B2(G107), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n785), .A2(new_n804), .B1(new_n806), .B2(new_n789), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n473), .B(new_n955), .C1(new_n956), .C2(KEYINPUT108), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(KEYINPUT108), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n952), .B2(KEYINPUT46), .ZN(new_n959));
  INV_X1    g0759(.A(new_n787), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n957), .B(new_n959), .C1(G283), .C2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(G317), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n961), .B1(new_n962), .B2(new_n791), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n954), .B(new_n963), .C1(G294), .C2(new_n855), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n854), .A2(G150), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n960), .A2(G50), .ZN(new_n966));
  AOI22_X1  g0766(.A1(G68), .A2(new_n797), .B1(new_n792), .B2(G137), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n966), .A2(new_n250), .A3(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n775), .A2(new_n216), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n777), .A2(new_n211), .ZN(new_n970));
  INV_X1    g0770(.A(G143), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n795), .A2(new_n575), .B1(new_n789), .B2(new_n971), .ZN(new_n972));
  NOR4_X1   g0772(.A1(new_n968), .A2(new_n969), .A3(new_n970), .A4(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n964), .B1(new_n965), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT110), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT47), .Z(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n770), .ZN(new_n977));
  INV_X1    g0777(.A(new_n827), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n978), .B1(new_n225), .B2(new_n359), .C1(new_n241), .C2(new_n818), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n557), .A2(new_n692), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n980), .A2(new_n550), .A3(new_n663), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n652), .B2(new_n980), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n982), .A2(new_n830), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n977), .A2(new_n814), .A3(new_n979), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n766), .A2(G1), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n521), .A2(new_n754), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n739), .A2(KEYINPUT93), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n986), .A2(new_n987), .B1(new_n511), .B2(new_n692), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n665), .A2(new_n691), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n707), .A2(KEYINPUT45), .A3(new_n695), .A4(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT45), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n694), .A2(new_n695), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n695), .B1(new_n993), .B2(new_n705), .ZN(new_n994));
  INV_X1    g0794(.A(new_n990), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n991), .A2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n998));
  NAND3_X1  g0798(.A1(new_n994), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n994), .A2(new_n995), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n998), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n997), .A2(new_n999), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n704), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n701), .A2(KEYINPUT90), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n701), .A2(KEYINPUT90), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1006), .A2(new_n1007), .A3(new_n993), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n704), .A2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(new_n705), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n761), .B1(new_n1005), .B2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n710), .B(KEYINPUT41), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n985), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n990), .A2(KEYINPUT103), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT103), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n988), .A2(new_n1016), .A3(new_n989), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1015), .A2(new_n656), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n520), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT104), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1018), .A2(KEYINPUT104), .A3(new_n520), .ZN(new_n1022));
  AND3_X1   g0822(.A1(new_n1021), .A2(new_n692), .A3(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n707), .A2(new_n755), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT42), .Z(new_n1025));
  OAI21_X1  g0825(.A(new_n1014), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT105), .Z(new_n1028));
  NAND4_X1  g0828(.A1(new_n1004), .A2(new_n1015), .A3(new_n1017), .A4(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1028), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1030), .B1(new_n704), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1026), .B(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT107), .ZN(new_n1035));
  NOR3_X1   g0835(.A1(new_n1013), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n985), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1003), .B(new_n704), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1009), .B(new_n706), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n760), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1012), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1037), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1033), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(new_n1026), .ZN(new_n1044));
  AOI21_X1  g0844(.A(KEYINPUT107), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n984), .B1(new_n1036), .B2(new_n1045), .ZN(G387));
  NAND2_X1  g0846(.A1(new_n993), .A2(new_n825), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n712), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1048), .A2(new_n225), .A3(new_n250), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(G107), .B2(new_n225), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT111), .Z(new_n1051));
  NOR3_X1   g0851(.A1(new_n284), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1048), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(G68), .A2(G77), .ZN(new_n1054));
  OAI21_X1  g0854(.A(KEYINPUT50), .B1(new_n284), .B2(G50), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1053), .A2(new_n271), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n817), .B(new_n1056), .C1(new_n237), .C2(new_n271), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n827), .B1(new_n1051), .B2(new_n1057), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n539), .A2(new_n797), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n775), .A2(new_n211), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1059), .B(new_n1060), .C1(new_n568), .C2(new_n855), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n778), .A2(G97), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n332), .A2(new_n785), .B1(new_n787), .B2(new_n328), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(G150), .B2(new_n792), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n473), .B1(new_n801), .B2(G159), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1061), .A2(new_n1062), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n854), .A2(G317), .B1(G311), .B2(new_n855), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1067), .B1(new_n804), .B2(new_n787), .C1(new_n803), .C2(new_n789), .ZN(new_n1068));
  XOR2_X1   g0868(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n1069));
  XNOR2_X1  g0869(.A(new_n1068), .B(new_n1069), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1070), .B1(new_n808), .B2(new_n798), .C1(new_n476), .C2(new_n775), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(KEYINPUT113), .B(KEYINPUT49), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1071), .B(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n457), .B1(G326), .B2(new_n792), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n369), .B2(new_n777), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1066), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n767), .B(new_n1058), .C1(new_n1076), .C2(new_n770), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1039), .A2(new_n985), .B1(new_n1047), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n710), .B1(new_n1039), .B2(new_n761), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1010), .A2(new_n760), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1078), .B1(new_n1079), .B2(new_n1080), .ZN(G393));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1038), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1080), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n1005), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1082), .A2(new_n710), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1038), .A2(new_n985), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1031), .A2(new_n825), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n770), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n785), .A2(new_n575), .B1(new_n290), .B2(new_n789), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT51), .Z(new_n1090));
  OAI221_X1 g0890(.A(new_n457), .B1(new_n333), .B2(new_n798), .C1(new_n775), .C2(new_n577), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n777), .A2(new_n443), .B1(new_n791), .B2(new_n971), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1093), .B1(new_n332), .B2(new_n795), .C1(new_n284), .C2(new_n787), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n775), .A2(new_n808), .B1(new_n803), .B2(new_n791), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT114), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n785), .A2(new_n806), .B1(new_n962), .B2(new_n789), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT52), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n787), .A2(new_n476), .ZN(new_n1102));
  NOR4_X1   g0902(.A1(new_n1097), .A2(new_n1100), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n797), .A2(G116), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n795), .A2(new_n804), .B1(new_n777), .B2(new_n435), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1103), .A2(new_n317), .A3(new_n1104), .A4(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1088), .B1(new_n1094), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n225), .A2(new_n318), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1109), .B(new_n827), .C1(new_n248), .C2(new_n817), .ZN(new_n1110));
  NOR3_X1   g0910(.A1(new_n1108), .A2(new_n767), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1087), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1085), .A2(new_n1086), .A3(new_n1112), .ZN(G390));
  OAI211_X1 g0913(.A(new_n841), .B(new_n929), .C1(new_n738), .C2(new_n746), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n757), .A2(new_n692), .A3(new_n837), .ZN(new_n1115));
  AND2_X1   g0915(.A1(new_n1115), .A2(new_n838), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n929), .B1(new_n920), .B2(new_n841), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1114), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n872), .B(G330), .C1(new_n743), .C2(new_n874), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(KEYINPUT115), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT115), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n914), .A2(new_n1122), .A3(G330), .A4(new_n872), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n929), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1124), .B1(new_n842), .B2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n931), .A2(new_n932), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1119), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n926), .B(new_n921), .C1(new_n682), .C2(new_n683), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n933), .A2(new_n940), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n939), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n911), .A2(new_n940), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1125), .B1(new_n1115), .B2(new_n838), .ZN(new_n1135));
  OR2_X1    g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1114), .A2(new_n1133), .A3(new_n1136), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n937), .A2(new_n938), .B1(new_n940), .B2(new_n933), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1124), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1131), .A2(new_n1141), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1143), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1142), .A2(new_n710), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT120), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1147));
  OAI21_X1  g0947(.A(G330), .B1(new_n743), .B2(new_n744), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(KEYINPUT92), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n839), .B(new_n1125), .C1(new_n1149), .C2(new_n745), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1140), .B(new_n985), .C1(new_n1147), .C2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT116), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1137), .A2(KEYINPUT116), .A3(new_n985), .A4(new_n1140), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n824), .B1(new_n937), .B2(new_n938), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n864), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n568), .A2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n787), .A2(new_n318), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n317), .B1(new_n775), .B2(new_n443), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1160), .B(KEYINPUT118), .Z(new_n1161));
  OAI22_X1  g0961(.A1(new_n798), .A2(new_n333), .B1(new_n785), .B2(new_n369), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT119), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n777), .A2(new_n328), .B1(new_n791), .B2(new_n476), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G107), .B2(new_n855), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1161), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1159), .B(new_n1166), .C1(G283), .C2(new_n801), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n775), .A2(new_n290), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n1169), .A2(KEYINPUT53), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n854), .A2(G132), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(KEYINPUT54), .B(G143), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT117), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1173), .A2(new_n960), .B1(G137), .B2(new_n855), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n317), .B1(new_n797), .B2(G159), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1170), .A2(new_n1171), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1169), .A2(KEYINPUT53), .B1(G125), .B2(new_n792), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n777), .A2(new_n332), .ZN(new_n1179));
  INV_X1    g0979(.A(G128), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n789), .A2(new_n1180), .ZN(new_n1181));
  NOR4_X1   g0981(.A1(new_n1176), .A2(new_n1178), .A3(new_n1179), .A4(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n770), .B1(new_n1167), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NOR4_X1   g0984(.A1(new_n1156), .A2(new_n767), .A3(new_n1158), .A4(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1146), .B1(new_n1155), .B2(new_n1186), .ZN(new_n1187));
  AOI211_X1 g0987(.A(KEYINPUT120), .B(new_n1185), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1145), .B1(new_n1187), .B2(new_n1188), .ZN(G378));
  INV_X1    g0989(.A(KEYINPUT57), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n941), .ZN(new_n1191));
  XOR2_X1   g0991(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n309), .A2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n309), .A2(new_n1193), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n301), .A2(new_n877), .ZN(new_n1196));
  OR3_X1    g0996(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1196), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n913), .B2(G330), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1199), .A2(new_n917), .A3(G330), .A4(new_n918), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1191), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1199), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n919), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1205), .A2(new_n941), .A3(new_n1201), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1190), .B1(new_n1203), .B2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n839), .B1(new_n1149), .B2(new_n745), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1123), .B(new_n1121), .C1(new_n1208), .C2(new_n929), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1127), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1117), .B1(new_n1208), .B2(new_n929), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1209), .A2(new_n1210), .B1(new_n1211), .B2(new_n1116), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1130), .B1(new_n1212), .B2(new_n1141), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n711), .B1(new_n1207), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1129), .B1(new_n1143), .B2(new_n1128), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT121), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1205), .A2(new_n941), .A3(new_n1201), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n941), .B1(new_n1205), .B2(new_n1201), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1216), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1206), .A2(KEYINPUT121), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1215), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1214), .B1(new_n1221), .B2(KEYINPUT57), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1204), .A2(new_n824), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n391), .A2(G33), .ZN(new_n1224));
  AOI21_X1  g1024(.A(G50), .B1(new_n1224), .B2(new_n270), .ZN(new_n1225));
  AOI21_X1  g1025(.A(G33), .B1(new_n792), .B2(G124), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n776), .A2(new_n1173), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n960), .A2(G137), .B1(G132), .B2(new_n855), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n801), .A2(G125), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n797), .A2(G150), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .A4(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(G128), .B2(new_n854), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT59), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n270), .B(new_n1226), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(G159), .B2(new_n778), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1225), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1060), .B1(G107), .B2(new_n854), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n778), .A2(G58), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1238), .B(new_n1239), .C1(new_n808), .C2(new_n791), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n539), .A2(new_n960), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n797), .A2(G68), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n457), .B1(new_n801), .B2(G116), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n855), .A2(G97), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .A4(new_n1244), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1240), .A2(new_n1245), .A3(G41), .ZN(new_n1246));
  XOR2_X1   g1046(.A(new_n1246), .B(KEYINPUT58), .Z(new_n1247));
  AOI21_X1  g1047(.A(new_n1088), .B1(new_n1237), .B2(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1157), .A2(G50), .ZN(new_n1249));
  NOR4_X1   g1049(.A1(new_n1223), .A2(new_n767), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1250), .B1(new_n1251), .B2(new_n985), .ZN(new_n1252));
  AND2_X1   g1052(.A1(new_n1222), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(G375));
  OAI211_X1 g1054(.A(new_n1129), .B(new_n1119), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1131), .A2(new_n1012), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1125), .A2(new_n823), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n775), .A2(new_n575), .B1(new_n1180), .B2(new_n791), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT122), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n473), .B1(new_n1173), .B2(new_n855), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1260), .B(new_n1239), .C1(new_n332), .C2(new_n798), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n801), .A2(G132), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n960), .A2(G150), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n854), .A2(G137), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .A4(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1059), .B1(G303), .B2(new_n792), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n795), .A2(new_n369), .B1(new_n777), .B2(new_n333), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(G107), .B2(new_n960), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n250), .B1(new_n854), .B2(G283), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1267), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  OAI221_X1 g1071(.A(new_n1271), .B1(new_n318), .B2(new_n775), .C1(new_n476), .C2(new_n789), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1088), .B1(new_n1266), .B2(new_n1272), .ZN(new_n1273));
  AOI211_X1 g1073(.A(new_n767), .B(new_n1273), .C1(new_n328), .C2(new_n864), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1274), .B(KEYINPUT123), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1128), .A2(new_n985), .B1(new_n1257), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1256), .A2(new_n1276), .ZN(G381));
  AOI21_X1  g1077(.A(new_n1185), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1145), .A2(new_n1278), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1253), .A2(new_n1279), .ZN(new_n1280));
  NOR3_X1   g1080(.A1(G387), .A2(G384), .A3(G381), .ZN(new_n1281));
  OR2_X1    g1081(.A1(G393), .A2(G396), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(G390), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1280), .A2(new_n1281), .A3(new_n1283), .ZN(G407));
  INV_X1    g1084(.A(G213), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1285), .B1(new_n1280), .B2(new_n690), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(G407), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(KEYINPUT124), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT124), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1286), .A2(new_n1289), .A3(G407), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1288), .A2(new_n1290), .ZN(G409));
  INV_X1    g1091(.A(new_n984), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1035), .B1(new_n1013), .B2(new_n1034), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1042), .A2(new_n1044), .A3(KEYINPUT107), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1292), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(G390), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT125), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G393), .A2(G396), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1282), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1296), .A2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1299), .B1(new_n1295), .B2(G390), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1085), .A2(new_n1086), .A3(new_n1112), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(G393), .B(new_n832), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(G387), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1301), .A2(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1300), .B1(new_n1305), .B2(new_n1296), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT61), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n689), .A2(new_n1285), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT60), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1255), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1311), .A2(KEYINPUT60), .A3(new_n1129), .A4(new_n1119), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1310), .A2(new_n1131), .A3(new_n1312), .A4(new_n710), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1276), .ZN(new_n1314));
  INV_X1    g1114(.A(G384), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1313), .A2(G384), .A3(new_n1276), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1222), .A2(G378), .A3(new_n1252), .ZN(new_n1319));
  AOI21_X1  g1119(.A(KEYINPUT121), .B1(new_n1203), .B2(new_n1206), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1220), .ZN(new_n1321));
  OAI211_X1 g1121(.A(new_n1012), .B(new_n1213), .C1(new_n1320), .C2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1203), .A2(new_n1206), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1250), .B1(new_n1323), .B2(new_n985), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n1279), .ZN(new_n1326));
  AOI211_X1 g1126(.A(new_n1308), .B(new_n1318), .C1(new_n1319), .C2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1307), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1319), .A2(new_n1326), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1308), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1318), .ZN(new_n1332));
  XOR2_X1   g1132(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1333));
  NAND4_X1  g1133(.A1(new_n1330), .A2(new_n1331), .A3(new_n1332), .A4(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1308), .B1(new_n1319), .B2(new_n1326), .ZN(new_n1335));
  AND3_X1   g1135(.A1(new_n1313), .A2(G384), .A3(new_n1276), .ZN(new_n1336));
  AOI21_X1  g1136(.A(G384), .B1(new_n1313), .B2(new_n1276), .ZN(new_n1337));
  OAI211_X1 g1137(.A(G2897), .B(new_n1308), .C1(new_n1336), .C2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1308), .A2(G2897), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1316), .A2(new_n1317), .A3(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1338), .A2(new_n1340), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1334), .B1(new_n1335), .B2(new_n1341), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1306), .B1(new_n1329), .B2(new_n1342), .ZN(new_n1343));
  OAI21_X1  g1143(.A(KEYINPUT63), .B1(new_n1335), .B2(new_n1341), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1335), .A2(new_n1332), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  AOI22_X1  g1146(.A1(G387), .A2(new_n1302), .B1(new_n1297), .B2(new_n1303), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1282), .A2(new_n1298), .ZN(new_n1348));
  NOR3_X1   g1148(.A1(new_n1295), .A2(G390), .A3(new_n1348), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1296), .B1(new_n1347), .B2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1300), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1327), .A2(KEYINPUT63), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1346), .A2(new_n1307), .A3(new_n1352), .A4(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1343), .A2(new_n1354), .ZN(G405));
  INV_X1    g1155(.A(new_n1279), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1319), .B1(new_n1253), .B2(new_n1356), .ZN(new_n1357));
  INV_X1    g1157(.A(KEYINPUT127), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1357), .A2(new_n1358), .A3(new_n1332), .ZN(new_n1359));
  OAI221_X1 g1159(.A(new_n1319), .B1(KEYINPUT127), .B2(new_n1318), .C1(new_n1253), .C2(new_n1356), .ZN(new_n1360));
  AND3_X1   g1160(.A1(new_n1306), .A2(new_n1359), .A3(new_n1360), .ZN(new_n1361));
  AOI21_X1  g1161(.A(new_n1306), .B1(new_n1359), .B2(new_n1360), .ZN(new_n1362));
  NOR2_X1   g1162(.A1(new_n1361), .A2(new_n1362), .ZN(G402));
endmodule


