//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n578, new_n579, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n452), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND3_X1   g037(.A1(new_n462), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(KEYINPUT67), .B1(new_n462), .B2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(G101), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI211_X1 g042(.A(G137), .B(new_n462), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g044(.A(G125), .B1(new_n466), .B2(new_n467), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n462), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n469), .A2(new_n472), .ZN(G160));
  OR2_X1    g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n462), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n462), .B1(new_n474), .B2(new_n475), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  OAI211_X1 g060(.A(G138), .B(new_n462), .C1(new_n466), .C2(new_n467), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT4), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n466), .A2(new_n467), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n490), .A2(new_n462), .A3(G138), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n488), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AND3_X1   g067(.A1(new_n490), .A2(new_n462), .A3(G138), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n476), .A2(KEYINPUT69), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n487), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n462), .A2(G114), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n497), .A2(new_n499), .A3(KEYINPUT68), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n501), .B1(new_n496), .B2(new_n498), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n500), .A2(new_n502), .B1(new_n480), .B2(G126), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n495), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  NAND2_X1  g080(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n509));
  OR2_X1    g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  XOR2_X1   g087(.A(KEYINPUT71), .B(G88), .Z(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G50), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n508), .A2(new_n509), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n514), .B(new_n516), .C1(new_n518), .C2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  NAND2_X1  g096(.A1(new_n515), .A2(G51), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  AND2_X1   g099(.A1(G63), .A2(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n517), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n522), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n512), .A2(G89), .ZN(new_n528));
  OAI21_X1  g103(.A(KEYINPUT72), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n515), .A2(G51), .B1(new_n517), .B2(new_n525), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n512), .A2(G89), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT72), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n530), .A2(new_n531), .A3(new_n532), .A4(new_n524), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n529), .A2(new_n533), .ZN(G168));
  XNOR2_X1  g109(.A(KEYINPUT6), .B(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n517), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n535), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G52), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n536), .A2(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n517), .A2(G64), .ZN(new_n541));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G651), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n540), .B1(new_n544), .B2(KEYINPUT73), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT73), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n543), .A2(new_n546), .A3(G651), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n545), .A2(new_n547), .ZN(G171));
  AOI22_X1  g123(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n519), .ZN(new_n550));
  INV_X1    g125(.A(G81), .ZN(new_n551));
  INV_X1    g126(.A(G43), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n536), .A2(new_n551), .B1(new_n538), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  INV_X1    g134(.A(G53), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT9), .B1(new_n538), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n515), .A2(new_n562), .A3(G53), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n561), .A2(new_n563), .B1(G91), .B2(new_n512), .ZN(new_n564));
  AND2_X1   g139(.A1(G78), .A2(G543), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n565), .B1(new_n517), .B2(G65), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(KEYINPUT74), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(new_n508), .B2(new_n509), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n568), .B1(new_n570), .B2(new_n565), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n567), .A2(G651), .A3(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n573));
  AND3_X1   g148(.A1(new_n564), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n573), .B1(new_n564), .B2(new_n572), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n574), .A2(new_n575), .ZN(G299));
  NAND2_X1  g151(.A1(new_n545), .A2(new_n547), .ZN(G301));
  AND3_X1   g152(.A1(new_n529), .A2(KEYINPUT76), .A3(new_n533), .ZN(new_n578));
  AOI21_X1  g153(.A(KEYINPUT76), .B1(new_n529), .B2(new_n533), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(G286));
  NAND2_X1  g155(.A1(new_n512), .A2(G87), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n515), .A2(G49), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(G288));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n585), .B1(new_n508), .B2(new_n509), .ZN(new_n586));
  AND2_X1   g161(.A1(G73), .A2(G543), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT77), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI211_X1 g165(.A(KEYINPUT77), .B(G651), .C1(new_n586), .C2(new_n587), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n512), .A2(G86), .B1(new_n515), .B2(G48), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(G305));
  AOI22_X1  g168(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(new_n519), .ZN(new_n595));
  INV_X1    g170(.A(G85), .ZN(new_n596));
  INV_X1    g171(.A(G47), .ZN(new_n597));
  OAI22_X1  g172(.A1(new_n536), .A2(new_n596), .B1(new_n538), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(KEYINPUT78), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT78), .ZN(new_n600));
  OAI221_X1 g175(.A(new_n600), .B1(new_n538), .B2(new_n597), .C1(new_n536), .C2(new_n596), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n595), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(new_n512), .A2(G92), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n604), .B(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n517), .A2(G66), .ZN(new_n607));
  INV_X1    g182(.A(G79), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(new_n507), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n609), .A2(G651), .B1(G54), .B2(new_n515), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G171), .B2(new_n612), .ZN(G284));
  OAI21_X1  g189(.A(new_n613), .B1(G171), .B2(new_n612), .ZN(G321));
  MUX2_X1   g190(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g191(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g192(.A(G860), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n611), .B1(G559), .B2(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT79), .ZN(G148));
  OAI21_X1  g195(.A(KEYINPUT80), .B1(new_n554), .B2(G868), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n611), .A2(G559), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  MUX2_X1   g198(.A(KEYINPUT80), .B(new_n621), .S(new_n623), .Z(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g200(.A1(new_n463), .A2(new_n464), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(new_n476), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT13), .Z(new_n630));
  INV_X1    g205(.A(G2100), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n480), .A2(G123), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n462), .A2(G111), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  INV_X1    g211(.A(G135), .ZN(new_n637));
  OAI221_X1 g212(.A(new_n634), .B1(new_n635), .B2(new_n636), .C1(new_n637), .C2(new_n477), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(G2096), .Z(new_n639));
  NAND3_X1  g214(.A1(new_n632), .A2(new_n633), .A3(new_n639), .ZN(G156));
  XOR2_X1   g215(.A(KEYINPUT15), .B(G2435), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2438), .ZN(new_n642));
  XOR2_X1   g217(.A(G2427), .B(G2430), .Z(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT83), .B(KEYINPUT14), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n642), .A2(new_n643), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G1341), .B(G1348), .Z(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(KEYINPUT82), .B(KEYINPUT16), .Z(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(G14), .B1(new_n652), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n656), .B2(new_n652), .ZN(G401));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(KEYINPUT18), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2072), .B(G2078), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2096), .B(G2100), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT84), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n664), .B(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT18), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n661), .A2(KEYINPUT17), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n659), .A2(new_n660), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n667), .B(new_n671), .Z(G227));
  XNOR2_X1  g247(.A(G1981), .B(G1986), .ZN(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT85), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1956), .B(G2474), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT20), .Z(new_n682));
  OR2_X1    g257(.A1(new_n675), .A2(new_n677), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n683), .A2(new_n680), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n683), .A2(new_n680), .A3(new_n678), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n682), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT86), .Z(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n686), .A2(new_n689), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n673), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n692), .ZN(new_n694));
  INV_X1    g269(.A(new_n673), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n694), .A2(new_n695), .A3(new_n690), .ZN(new_n696));
  XOR2_X1   g271(.A(G1991), .B(G1996), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT88), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT87), .ZN(new_n699));
  AND3_X1   g274(.A1(new_n693), .A2(new_n696), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n699), .B1(new_n693), .B2(new_n696), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(G229));
  AND2_X1   g277(.A1(new_n606), .A2(new_n610), .ZN(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G4), .B2(new_n704), .ZN(new_n706));
  INV_X1    g281(.A(G1348), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G2072), .ZN(new_n709));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n710), .A2(G33), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT25), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G139), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n477), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n717), .A2(new_n462), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT92), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n711), .B1(new_n721), .B2(G29), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n708), .B1(new_n709), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(new_n709), .B2(new_n722), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n710), .A2(G32), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n478), .A2(G141), .B1(new_n626), .B2(G105), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n480), .A2(G129), .ZN(new_n727));
  NAND3_X1  g302(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT26), .Z(new_n729));
  NAND3_X1  g304(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n725), .B1(new_n731), .B2(new_n710), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT27), .Z(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(G1996), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n704), .A2(G19), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n554), .B2(new_n704), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1341), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n706), .A2(new_n707), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n710), .A2(G35), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G162), .B2(new_n710), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT29), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n738), .B1(G2090), .B2(new_n741), .ZN(new_n742));
  NOR4_X1   g317(.A1(new_n724), .A2(new_n734), .A3(new_n737), .A4(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(G16), .A2(G21), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G168), .B2(G16), .ZN(new_n745));
  INV_X1    g320(.A(G1966), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n741), .A2(G2090), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT95), .Z(new_n749));
  NAND3_X1  g324(.A1(new_n743), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(G299), .A2(G16), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n704), .A2(G20), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT23), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1956), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT31), .B(G11), .Z(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT94), .B(KEYINPUT30), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n757), .A2(G28), .ZN(new_n758));
  AOI21_X1  g333(.A(G29), .B1(new_n757), .B2(G28), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n756), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G34), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(KEYINPUT24), .ZN(new_n762));
  AOI21_X1  g337(.A(G29), .B1(new_n761), .B2(KEYINPUT24), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n762), .B1(new_n763), .B2(KEYINPUT93), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(KEYINPUT93), .B2(new_n763), .ZN(new_n765));
  INV_X1    g340(.A(G160), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n765), .B1(new_n766), .B2(new_n710), .ZN(new_n767));
  INV_X1    g342(.A(G2084), .ZN(new_n768));
  OAI221_X1 g343(.A(new_n760), .B1(new_n710), .B2(new_n638), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n710), .A2(G26), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT91), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT28), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n478), .A2(G140), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n480), .A2(G128), .ZN(new_n774));
  OR2_X1    g349(.A1(G104), .A2(G2105), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n775), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n773), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n772), .B1(new_n778), .B2(new_n710), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G2067), .ZN(new_n780));
  AOI211_X1 g355(.A(new_n769), .B(new_n780), .C1(new_n768), .C2(new_n767), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n710), .A2(G27), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G164), .B2(new_n710), .ZN(new_n783));
  INV_X1    g358(.A(G2078), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n733), .A2(G1996), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n704), .A2(G5), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G171), .B2(new_n704), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(G1961), .Z(new_n789));
  NAND4_X1  g364(.A1(new_n781), .A2(new_n785), .A3(new_n786), .A4(new_n789), .ZN(new_n790));
  NOR3_X1   g365(.A1(new_n750), .A2(new_n755), .A3(new_n790), .ZN(new_n791));
  MUX2_X1   g366(.A(G6), .B(G305), .S(G16), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT90), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT32), .B(G1981), .Z(new_n794));
  OR2_X1    g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n704), .A2(G22), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G166), .B2(new_n704), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(G1971), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n704), .A2(G23), .ZN(new_n800));
  INV_X1    g375(.A(G288), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(new_n704), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT33), .B(G1976), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n795), .A2(new_n796), .A3(new_n799), .A4(new_n804), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(KEYINPUT34), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(KEYINPUT34), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n710), .A2(G25), .ZN(new_n808));
  OAI21_X1  g383(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n809));
  INV_X1    g384(.A(G107), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n809), .B1(new_n810), .B2(G2105), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n480), .A2(G119), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT89), .ZN(new_n813));
  AOI211_X1 g388(.A(new_n811), .B(new_n813), .C1(G131), .C2(new_n478), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n808), .B1(new_n814), .B2(new_n710), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT35), .B(G1991), .Z(new_n816));
  XOR2_X1   g391(.A(new_n815), .B(new_n816), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n704), .A2(G24), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n602), .B2(new_n704), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(G1986), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n819), .A2(G1986), .ZN(new_n821));
  NOR3_X1   g396(.A1(new_n817), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n806), .A2(new_n807), .A3(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT36), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n791), .A2(new_n824), .ZN(G150));
  INV_X1    g400(.A(G150), .ZN(G311));
  AOI22_X1  g401(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n827), .A2(new_n519), .ZN(new_n828));
  INV_X1    g403(.A(G93), .ZN(new_n829));
  INV_X1    g404(.A(G55), .ZN(new_n830));
  OAI22_X1  g405(.A1(new_n536), .A2(new_n829), .B1(new_n538), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n832), .A2(new_n618), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT37), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n703), .A2(G559), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT96), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT38), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n554), .B(new_n832), .Z(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n837), .B(new_n839), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n618), .B1(new_n840), .B2(KEYINPUT39), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n834), .B1(new_n841), .B2(new_n842), .ZN(G145));
  XNOR2_X1  g418(.A(new_n638), .B(G160), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(G162), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n777), .B(new_n504), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n721), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n730), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n480), .A2(G130), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n462), .A2(G118), .ZN(new_n850));
  OAI21_X1  g425(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(G142), .B2(new_n478), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n629), .B(new_n853), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n814), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n848), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT97), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n848), .A2(new_n855), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT98), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n845), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n856), .A2(new_n845), .ZN(new_n862));
  AOI21_X1  g437(.A(G37), .B1(new_n862), .B2(new_n858), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n861), .A2(new_n863), .A3(new_n865), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(G395));
  OR2_X1    g444(.A1(new_n602), .A2(G305), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n602), .A2(G305), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(G303), .B(G288), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n870), .A2(new_n873), .A3(new_n871), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n564), .A2(new_n572), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(KEYINPUT75), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n564), .A2(new_n572), .A3(new_n573), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n703), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n611), .B1(new_n574), .B2(new_n575), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n881), .A2(new_n882), .A3(KEYINPUT41), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT41), .B1(new_n881), .B2(new_n882), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n838), .B(new_n622), .ZN(new_n887));
  MUX2_X1   g462(.A(new_n883), .B(new_n886), .S(new_n887), .Z(new_n888));
  AND2_X1   g463(.A1(new_n888), .A2(KEYINPUT42), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(KEYINPUT42), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n877), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n888), .A2(KEYINPUT42), .ZN(new_n892));
  INV_X1    g467(.A(new_n877), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n888), .A2(KEYINPUT42), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AND4_X1   g470(.A1(KEYINPUT100), .A2(new_n891), .A3(new_n895), .A4(G868), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n891), .A2(new_n895), .A3(G868), .ZN(new_n897));
  INV_X1    g472(.A(new_n832), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT100), .B1(new_n898), .B2(new_n612), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n896), .B1(new_n897), .B2(new_n899), .ZN(G295));
  AOI21_X1  g475(.A(new_n896), .B1(new_n897), .B2(new_n899), .ZN(G331));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n903));
  INV_X1    g478(.A(G37), .ZN(new_n904));
  OAI21_X1  g479(.A(G171), .B1(new_n578), .B2(new_n579), .ZN(new_n905));
  NAND3_X1  g480(.A1(G301), .A2(new_n533), .A3(new_n529), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI22_X1  g482(.A1(new_n907), .A2(new_n839), .B1(new_n881), .B2(new_n882), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n905), .A2(new_n838), .A3(new_n906), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n905), .A2(new_n838), .A3(KEYINPUT101), .A4(new_n906), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n908), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n909), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n838), .B1(new_n905), .B2(new_n906), .ZN(new_n915));
  OAI22_X1  g490(.A1(new_n914), .A2(new_n915), .B1(new_n884), .B2(new_n885), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n913), .A2(new_n916), .A3(new_n877), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n907), .A2(new_n839), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n911), .A2(new_n918), .A3(new_n912), .ZN(new_n919));
  AOI22_X1  g494(.A1(new_n919), .A2(new_n886), .B1(new_n909), .B2(new_n908), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n875), .A2(KEYINPUT102), .A3(new_n876), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT102), .B1(new_n875), .B2(new_n876), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n904), .B(new_n917), .C1(new_n920), .C2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n903), .B1(new_n924), .B2(KEYINPUT43), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n917), .A2(new_n904), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n913), .A2(new_n916), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n921), .A2(new_n922), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n927), .A2(KEYINPUT103), .A3(new_n928), .A4(new_n931), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n931), .A2(new_n928), .A3(new_n904), .A4(new_n917), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT103), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n925), .A2(new_n932), .A3(new_n935), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n920), .A2(new_n923), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n937), .A2(new_n927), .A3(new_n928), .ZN(new_n938));
  INV_X1    g513(.A(new_n931), .ZN(new_n939));
  OAI21_X1  g514(.A(KEYINPUT43), .B1(new_n939), .B2(new_n926), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT44), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n902), .B1(new_n936), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n938), .A2(new_n940), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n903), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n925), .A2(new_n932), .A3(new_n935), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(KEYINPUT104), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n942), .A2(new_n946), .ZN(G397));
  NAND2_X1  g522(.A1(new_n515), .A2(G48), .ZN(new_n948));
  INV_X1    g523(.A(G86), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n948), .B1(new_n536), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT113), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n948), .B(KEYINPUT113), .C1(new_n536), .C2(new_n949), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n952), .A2(new_n591), .A3(new_n590), .A4(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(G1981), .ZN(new_n955));
  INV_X1    g530(.A(G1981), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n590), .A2(new_n956), .A3(new_n591), .A4(new_n592), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n957), .A2(KEYINPUT112), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(KEYINPUT112), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n955), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT49), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n955), .B(KEYINPUT49), .C1(new_n958), .C2(new_n959), .ZN(new_n963));
  INV_X1    g538(.A(G8), .ZN(new_n964));
  AOI21_X1  g539(.A(G1384), .B1(new_n495), .B2(new_n503), .ZN(new_n965));
  XOR2_X1   g540(.A(KEYINPUT105), .B(G40), .Z(new_n966));
  NOR3_X1   g541(.A1(new_n469), .A2(new_n472), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n964), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n962), .A2(new_n963), .A3(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n970));
  NAND3_X1  g545(.A1(G303), .A2(G8), .A3(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  AOI22_X1  g547(.A1(G303), .A2(G8), .B1(KEYINPUT109), .B2(KEYINPUT55), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n975), .A2(G1384), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n504), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n977), .B(new_n967), .C1(KEYINPUT45), .C2(new_n965), .ZN(new_n978));
  XOR2_X1   g553(.A(KEYINPUT108), .B(G1971), .Z(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G1384), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n504), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT50), .ZN(new_n983));
  INV_X1    g558(.A(G2090), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT50), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n965), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n983), .A2(new_n984), .A3(new_n967), .A4(new_n986), .ZN(new_n987));
  AOI211_X1 g562(.A(new_n964), .B(new_n974), .C1(new_n980), .C2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n504), .A2(new_n967), .A3(new_n981), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n581), .A2(G1976), .A3(new_n582), .A4(new_n583), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n990), .A2(G8), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT110), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n989), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n968), .A2(KEYINPUT110), .A3(new_n991), .ZN(new_n995));
  INV_X1    g570(.A(G1976), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT52), .B1(G288), .B2(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n990), .A2(G8), .A3(new_n991), .A4(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT111), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n968), .A2(new_n1000), .A3(new_n991), .A4(new_n997), .ZN(new_n1001));
  AOI22_X1  g576(.A1(new_n994), .A2(new_n995), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n969), .A2(new_n988), .A3(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n969), .A2(new_n996), .A3(new_n801), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n958), .A2(new_n959), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1003), .B1(new_n1006), .B2(new_n968), .ZN(new_n1007));
  INV_X1    g582(.A(new_n472), .ZN(new_n1008));
  INV_X1    g583(.A(new_n966), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1008), .A2(new_n465), .A3(new_n468), .A4(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1010), .B1(new_n982), .B2(KEYINPUT50), .ZN(new_n1011));
  XOR2_X1   g586(.A(KEYINPUT116), .B(G2084), .Z(new_n1012));
  AOI21_X1  g587(.A(new_n1012), .B1(new_n965), .B2(new_n985), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n746), .A2(new_n978), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  NOR3_X1   g589(.A1(new_n1014), .A2(new_n964), .A3(G286), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n964), .B1(new_n980), .B2(new_n987), .ZN(new_n1016));
  INV_X1    g591(.A(new_n974), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n969), .A2(new_n1002), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT63), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n967), .B1(new_n965), .B2(new_n985), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g598(.A(KEYINPUT114), .B(new_n967), .C1(new_n965), .C2(new_n985), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1023), .A2(new_n984), .A3(new_n986), .A4(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n980), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(G8), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n988), .B1(new_n1027), .B2(new_n974), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n969), .A2(KEYINPUT115), .A3(new_n1002), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT115), .B1(new_n969), .B2(new_n1002), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1028), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OR4_X1    g606(.A1(KEYINPUT63), .A2(new_n1014), .A3(new_n964), .A4(G286), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1007), .B(new_n1020), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(G168), .A2(new_n964), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1014), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT51), .ZN(new_n1037));
  AOI211_X1 g612(.A(new_n1037), .B(new_n964), .C1(new_n1014), .C2(G168), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT121), .B1(new_n1014), .B2(new_n964), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT121), .ZN(new_n1040));
  INV_X1    g615(.A(new_n986), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1041), .A2(new_n1021), .A3(new_n1012), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n982), .A2(new_n975), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1010), .B1(new_n504), .B2(new_n976), .ZN(new_n1044));
  AOI21_X1  g619(.A(G1966), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1040), .B(G8), .C1(new_n1042), .C2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1034), .A2(KEYINPUT51), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1039), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1038), .B1(new_n1048), .B2(KEYINPUT122), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT122), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1039), .A2(new_n1046), .A3(new_n1050), .A4(new_n1047), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1036), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g627(.A(G301), .B(KEYINPUT54), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n977), .A2(new_n967), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n965), .A2(KEYINPUT45), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT53), .B1(new_n1056), .B2(new_n784), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1058), .A2(G2078), .ZN(new_n1059));
  AND4_X1   g634(.A1(G40), .A2(new_n977), .A3(G160), .A4(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1057), .B1(new_n1043), .B2(new_n1060), .ZN(new_n1061));
  XOR2_X1   g636(.A(KEYINPUT123), .B(G1961), .Z(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(new_n1041), .B2(new_n1021), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1053), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT124), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1062), .B1(new_n1011), .B2(new_n986), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1059), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1054), .A2(new_n1055), .A3(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1066), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1043), .A2(new_n1044), .A3(new_n1059), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1064), .A2(new_n1071), .A3(KEYINPUT124), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1057), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1065), .B1(new_n1073), .B2(new_n1053), .ZN(new_n1074));
  NOR3_X1   g649(.A1(new_n1052), .A2(new_n1031), .A3(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1023), .A2(new_n986), .A3(new_n1024), .ZN(new_n1076));
  INV_X1    g651(.A(G1956), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  XOR2_X1   g653(.A(new_n878), .B(KEYINPUT57), .Z(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT56), .B(G2072), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1056), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1078), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1079), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n707), .B1(new_n1041), .B2(new_n1021), .ZN(new_n1084));
  INV_X1    g659(.A(new_n990), .ZN(new_n1085));
  INV_X1    g660(.A(G2067), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n611), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1082), .B1(new_n1083), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OR2_X1    g666(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1079), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1041), .B1(new_n1022), .B2(new_n1021), .ZN(new_n1094));
  AOI21_X1  g669(.A(G1956), .B1(new_n1094), .B2(new_n1024), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1081), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1093), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT61), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1097), .A2(new_n1098), .A3(new_n1082), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1098), .B1(new_n1097), .B2(new_n1082), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1102), .B1(new_n606), .B2(new_n610), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT60), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1103), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n611), .A2(KEYINPUT119), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1108), .A2(new_n1103), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1109), .A2(KEYINPUT60), .A3(new_n1087), .A4(new_n1084), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1106), .A2(new_n1107), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT120), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1106), .A2(new_n1107), .A3(KEYINPUT120), .A4(new_n1110), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT118), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n978), .A2(G1996), .ZN(new_n1116));
  XNOR2_X1  g691(.A(KEYINPUT58), .B(G1341), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1085), .A2(new_n1117), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1115), .B(new_n554), .C1(new_n1116), .C2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n1119), .B(KEYINPUT59), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1113), .A2(new_n1114), .A3(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1091), .B(new_n1092), .C1(new_n1101), .C2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1033), .B1(new_n1075), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1057), .ZN(new_n1125));
  AOI21_X1  g700(.A(G301), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1028), .B(new_n1126), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT62), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1128), .B1(new_n1052), .B2(new_n1129), .ZN(new_n1130));
  AOI211_X1 g705(.A(KEYINPUT62), .B(new_n1036), .C1(new_n1049), .C2(new_n1051), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT125), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1048), .A2(KEYINPUT122), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1038), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1133), .A2(new_n1134), .A3(new_n1051), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1036), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT62), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1052), .A2(new_n1129), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT125), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .A4(new_n1128), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1123), .A2(new_n1132), .A3(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1043), .A2(new_n1010), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1143), .B(KEYINPUT106), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n777), .B(new_n1086), .ZN(new_n1145));
  INV_X1    g720(.A(G1996), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1145), .B1(new_n1146), .B2(new_n731), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1148), .B1(new_n730), .B2(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n814), .B(new_n816), .ZN(new_n1151));
  XOR2_X1   g726(.A(new_n1151), .B(KEYINPUT107), .Z(new_n1152));
  AOI21_X1  g727(.A(new_n1150), .B1(new_n1152), .B2(new_n1144), .ZN(new_n1153));
  XOR2_X1   g728(.A(new_n602), .B(G1986), .Z(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(new_n1143), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1142), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT46), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1149), .A2(new_n1158), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n1159), .B(KEYINPUT126), .Z(new_n1160));
  INV_X1    g735(.A(new_n1145), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1144), .B1(new_n730), .B2(new_n1161), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1160), .B(new_n1162), .C1(new_n1158), .C2(new_n1149), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1163), .B(KEYINPUT47), .ZN(new_n1164));
  NOR4_X1   g739(.A1(G290), .A2(new_n1043), .A3(G1986), .A4(new_n1010), .ZN(new_n1165));
  XOR2_X1   g740(.A(new_n1165), .B(KEYINPUT48), .Z(new_n1166));
  NAND2_X1  g741(.A1(new_n1153), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n814), .A2(new_n816), .ZN(new_n1169));
  OAI22_X1  g744(.A1(new_n1150), .A2(new_n1169), .B1(G2067), .B2(new_n777), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1168), .B1(new_n1144), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1157), .A2(new_n1171), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g747(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1174));
  OAI21_X1  g748(.A(new_n1174), .B1(new_n700), .B2(new_n701), .ZN(new_n1175));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n1176));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  OAI211_X1 g751(.A(KEYINPUT127), .B(new_n1174), .C1(new_n700), .C2(new_n701), .ZN(new_n1178));
  NAND2_X1  g752(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g753(.A1(new_n864), .A2(new_n1179), .A3(new_n943), .ZN(G225));
  INV_X1    g754(.A(G225), .ZN(G308));
endmodule


