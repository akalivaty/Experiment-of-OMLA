//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020;
  INV_X1    g000(.A(G134), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT11), .B1(new_n187), .B2(G137), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G134), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT66), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n193), .B1(new_n190), .B2(G134), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n187), .A2(KEYINPUT66), .A3(G137), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G131), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n192), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n197), .B1(new_n192), .B2(new_n196), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT65), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT64), .B(G143), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(new_n203), .ZN(new_n207));
  AND2_X1   g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(KEYINPUT64), .ZN(new_n212));
  OAI211_X1 g026(.A(KEYINPUT65), .B(G146), .C1(new_n210), .C2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n207), .A2(new_n208), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(KEYINPUT64), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n209), .A2(G143), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(new_n203), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n211), .A2(G146), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(KEYINPUT0), .A2(G128), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n208), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n214), .A2(KEYINPUT67), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(KEYINPUT67), .B1(new_n214), .B2(new_n222), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n202), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(G116), .B(G119), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT2), .B(G113), .ZN(new_n227));
  XNOR2_X1  g041(.A(new_n226), .B(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G128), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n229), .B1(new_n204), .B2(KEYINPUT1), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n207), .A2(new_n213), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n230), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n219), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n190), .A2(G134), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n187), .A2(G137), .ZN(new_n236));
  OAI21_X1  g050(.A(G131), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n234), .A2(new_n198), .A3(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n225), .A2(new_n228), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G237), .ZN(new_n240));
  INV_X1    g054(.A(G953), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n240), .A2(new_n241), .A3(G210), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT27), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n244), .B(KEYINPUT26), .ZN(new_n245));
  INV_X1    g059(.A(G101), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n245), .B(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n239), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT68), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n225), .A2(KEYINPUT30), .A3(new_n238), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT30), .ZN(new_n251));
  INV_X1    g065(.A(new_n238), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n214), .A2(new_n222), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n201), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n251), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n228), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n250), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n239), .A2(new_n258), .A3(new_n247), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n249), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT31), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n247), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n256), .B1(new_n252), .B2(new_n254), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n239), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT28), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT28), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n239), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n265), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n269), .B1(new_n239), .B2(new_n266), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n272), .A2(KEYINPUT70), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n264), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n249), .A2(new_n257), .A3(new_n259), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT31), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n260), .A2(KEYINPUT69), .A3(KEYINPUT31), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n263), .A2(new_n274), .A3(new_n277), .A4(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(G472), .A2(G902), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT32), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n279), .A2(KEYINPUT32), .A3(new_n280), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT29), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n257), .A2(new_n239), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n264), .ZN(new_n287));
  INV_X1    g101(.A(new_n270), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT70), .B1(new_n288), .B2(new_n272), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n268), .A2(new_n265), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n285), .B(new_n287), .C1(new_n291), .C2(new_n264), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT67), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n253), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n214), .A2(KEYINPUT67), .A3(new_n222), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n201), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n256), .B1(new_n296), .B2(new_n252), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n269), .B1(new_n297), .B2(new_n239), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n298), .A2(new_n288), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n264), .A2(new_n285), .ZN(new_n300));
  AOI21_X1  g114(.A(G902), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n292), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G472), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n283), .A2(new_n284), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n229), .A2(G119), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n229), .A2(G119), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT23), .ZN(new_n307));
  OAI211_X1 g121(.A(KEYINPUT71), .B(new_n305), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n307), .A2(KEYINPUT71), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n308), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n305), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n311), .A2(new_n306), .ZN(new_n312));
  XOR2_X1   g126(.A(KEYINPUT24), .B(G110), .Z(new_n313));
  OAI22_X1  g127(.A1(new_n310), .A2(G110), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G125), .ZN(new_n315));
  NOR3_X1   g129(.A1(new_n315), .A2(KEYINPUT16), .A3(G140), .ZN(new_n316));
  NAND2_X1  g130(.A1(KEYINPUT73), .A2(G125), .ZN(new_n317));
  INV_X1    g131(.A(G140), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n317), .B(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n316), .B1(new_n319), .B2(KEYINPUT16), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G146), .ZN(new_n321));
  XOR2_X1   g135(.A(G125), .B(G140), .Z(new_n322));
  OR2_X1    g136(.A1(new_n322), .A2(G146), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n314), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n317), .B(G140), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT16), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n203), .B1(new_n327), .B2(new_n316), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(new_n321), .A3(KEYINPUT74), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT74), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n320), .A2(new_n330), .A3(G146), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n312), .A2(new_n313), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n329), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n310), .A2(G110), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(KEYINPUT72), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n324), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n241), .A2(G221), .A3(G234), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n337), .B(KEYINPUT75), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(KEYINPUT22), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n339), .B(new_n190), .ZN(new_n340));
  OR2_X1    g154(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n336), .A2(new_n340), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G217), .ZN(new_n345));
  INV_X1    g159(.A(G902), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n345), .B1(G234), .B2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n347), .A2(G902), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n348), .B(KEYINPUT76), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n341), .A2(new_n346), .A3(new_n342), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT25), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n341), .A2(KEYINPUT25), .A3(new_n346), .A4(new_n342), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n347), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n350), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n304), .A2(new_n358), .ZN(new_n359));
  XOR2_X1   g173(.A(KEYINPUT9), .B(G234), .Z(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(G221), .B1(new_n361), .B2(G902), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G469), .ZN(new_n364));
  INV_X1    g178(.A(G104), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT3), .B1(new_n365), .B2(G107), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT3), .ZN(new_n367));
  INV_X1    g181(.A(G107), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n368), .A3(G104), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n365), .A2(G107), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n370), .A2(KEYINPUT77), .A3(new_n246), .A4(new_n371), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n366), .A2(new_n369), .A3(new_n246), .A4(new_n371), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT77), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n368), .A2(G104), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n371), .A2(new_n376), .ZN(new_n377));
  AOI22_X1  g191(.A1(new_n372), .A2(new_n375), .B1(G101), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n379));
  AOI22_X1  g193(.A1(new_n207), .A2(new_n213), .B1(new_n379), .B2(G128), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT78), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n231), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n207), .A2(new_n213), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n379), .A2(G128), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(new_n381), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n378), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT10), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n378), .A2(KEYINPUT10), .A3(new_n234), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT79), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n378), .A2(KEYINPUT79), .A3(new_n234), .A4(KEYINPUT10), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n373), .B(KEYINPUT77), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n366), .A2(new_n369), .A3(new_n371), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G101), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT4), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  OR2_X1    g213(.A1(new_n397), .A2(KEYINPUT4), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n294), .A2(new_n295), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n389), .A2(new_n394), .A3(new_n201), .A4(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(G110), .B(G140), .ZN(new_n406));
  INV_X1    g220(.A(G227), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n407), .A2(G953), .ZN(new_n408));
  XOR2_X1   g222(.A(new_n406), .B(new_n408), .Z(new_n409));
  NOR2_X1   g223(.A1(new_n378), .A2(new_n234), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n387), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(KEYINPUT12), .B1(new_n412), .B2(new_n202), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT12), .ZN(new_n414));
  AOI211_X1 g228(.A(new_n414), .B(new_n201), .C1(new_n387), .C2(new_n411), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n405), .B(new_n409), .C1(new_n413), .C2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n389), .A2(new_n394), .A3(new_n404), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n202), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n409), .B1(new_n419), .B2(new_n405), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n364), .B(new_n346), .C1(new_n417), .C2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT80), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n405), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n387), .A2(new_n388), .B1(new_n402), .B2(new_n403), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n201), .B1(new_n425), .B2(new_n394), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n416), .B1(new_n427), .B2(new_n409), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n428), .A2(KEYINPUT80), .A3(new_n364), .A4(new_n346), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n423), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n419), .A2(new_n405), .A3(new_n409), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n389), .A2(new_n394), .A3(new_n404), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n412), .A2(KEYINPUT12), .A3(new_n202), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n383), .A2(new_n384), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT78), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(new_n231), .A3(new_n385), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n410), .B1(new_n436), .B2(new_n378), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n414), .B1(new_n437), .B2(new_n201), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n432), .A2(new_n201), .B1(new_n433), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n431), .B1(new_n439), .B2(new_n409), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n346), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G469), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n363), .B1(new_n430), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(G214), .B1(G237), .B2(G902), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT85), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n256), .B(new_n400), .C1(new_n395), .C2(new_n398), .ZN(new_n446));
  INV_X1    g260(.A(new_n226), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(new_n227), .ZN(new_n448));
  INV_X1    g262(.A(G116), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n449), .A2(KEYINPUT5), .A3(G119), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n450), .B1(new_n226), .B2(KEYINPUT5), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n448), .B1(G113), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n378), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g267(.A(G110), .B(G122), .Z(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n446), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT81), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n446), .A2(new_n453), .A3(KEYINPUT81), .A4(new_n455), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n231), .A2(new_n315), .A3(new_n233), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n315), .B1(new_n214), .B2(new_n222), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT84), .ZN(new_n465));
  XOR2_X1   g279(.A(KEYINPUT82), .B(G224), .Z(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n241), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT7), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n253), .A2(G125), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n469), .A2(KEYINPUT7), .A3(new_n461), .A4(new_n467), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(KEYINPUT84), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  XOR2_X1   g286(.A(new_n454), .B(KEYINPUT8), .Z(new_n473));
  INV_X1    g287(.A(KEYINPUT83), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n377), .A2(G101), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n373), .A2(new_n374), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n373), .A2(new_n374), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n451), .A2(G113), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n479), .B1(new_n447), .B2(new_n227), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n474), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n478), .A2(new_n480), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR3_X1   g297(.A1(new_n478), .A2(new_n480), .A3(new_n474), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n473), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n464), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n467), .A2(KEYINPUT7), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n460), .A2(new_n472), .A3(new_n485), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n346), .ZN(new_n490));
  INV_X1    g304(.A(new_n467), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n491), .B1(new_n462), .B2(new_n463), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n469), .A2(new_n461), .A3(new_n467), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI211_X1 g308(.A(KEYINPUT6), .B(new_n455), .C1(new_n446), .C2(new_n453), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n455), .B1(new_n446), .B2(new_n453), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT6), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI211_X1 g312(.A(new_n494), .B(new_n495), .C1(new_n460), .C2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n445), .B1(new_n490), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(G210), .B1(G237), .B2(G902), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  AOI22_X1  g316(.A1(new_n458), .A2(new_n459), .B1(new_n468), .B2(new_n471), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT83), .B1(new_n378), .B2(new_n452), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n453), .ZN(new_n505));
  INV_X1    g319(.A(new_n484), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n507), .A2(new_n473), .B1(new_n486), .B2(new_n487), .ZN(new_n508));
  AOI21_X1  g322(.A(G902), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n460), .A2(new_n498), .ZN(new_n510));
  INV_X1    g324(.A(new_n494), .ZN(new_n511));
  INV_X1    g325(.A(new_n495), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n509), .A2(new_n513), .A3(KEYINPUT85), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n500), .A2(new_n502), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT86), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n509), .A2(new_n513), .A3(new_n501), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT86), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n500), .A2(new_n518), .A3(new_n502), .A4(new_n514), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n443), .A2(new_n444), .A3(new_n520), .ZN(new_n521));
  XOR2_X1   g335(.A(KEYINPUT91), .B(KEYINPUT13), .Z(new_n522));
  OAI211_X1 g336(.A(new_n522), .B(G128), .C1(new_n210), .C2(new_n212), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n229), .A2(G143), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n524), .B1(new_n206), .B2(new_n229), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n523), .B(G134), .C1(new_n525), .C2(new_n522), .ZN(new_n526));
  INV_X1    g340(.A(G122), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(G116), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(KEYINPUT90), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n529), .B1(new_n449), .B2(G122), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n530), .A2(new_n368), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT90), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n528), .B(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n533), .B1(G116), .B2(new_n527), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(G107), .ZN(new_n535));
  OAI221_X1 g349(.A(new_n526), .B1(G134), .B2(new_n525), .C1(new_n531), .C2(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n530), .B1(KEYINPUT14), .B2(new_n368), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n533), .A2(KEYINPUT14), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n534), .A2(G107), .A3(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n525), .A2(G134), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n525), .A2(G134), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n537), .B(new_n539), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n361), .A2(new_n345), .A3(G953), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT92), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n536), .A2(new_n542), .A3(new_n544), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n536), .A2(KEYINPUT92), .A3(new_n542), .A4(new_n544), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(new_n346), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G478), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(KEYINPUT15), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n551), .B(new_n553), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n240), .A2(new_n241), .A3(G214), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT87), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n555), .B(new_n211), .C1(new_n209), .C2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n240), .A2(new_n241), .A3(G214), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n558), .B1(new_n206), .B2(KEYINPUT87), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n557), .A2(new_n559), .A3(G131), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n329), .A2(new_n331), .B1(KEYINPUT17), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT88), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n557), .A2(new_n559), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n197), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n560), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n563), .B1(new_n566), .B2(KEYINPUT17), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT17), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n565), .A2(KEYINPUT88), .A3(new_n568), .A4(new_n560), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n562), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(G113), .B(G122), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(new_n365), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n561), .A2(KEYINPUT18), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n323), .B1(new_n319), .B2(new_n203), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT18), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n564), .B1(new_n575), .B2(new_n197), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n573), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n570), .A2(new_n572), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n572), .B1(new_n570), .B2(new_n577), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n346), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(G475), .ZN(new_n582));
  NOR2_X1   g396(.A1(G475), .A2(G902), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n572), .ZN(new_n585));
  INV_X1    g399(.A(new_n577), .ZN(new_n586));
  MUX2_X1   g400(.A(new_n322), .B(new_n319), .S(KEYINPUT19), .Z(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n203), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n566), .A2(new_n321), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n585), .B1(new_n586), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n584), .B1(new_n578), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT20), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n578), .A2(new_n590), .ZN(new_n594));
  XOR2_X1   g408(.A(new_n583), .B(KEYINPUT89), .Z(new_n595));
  AND3_X1   g409(.A1(new_n594), .A2(new_n592), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n582), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(G234), .A2(G237), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(G952), .A3(new_n241), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT21), .B(G898), .Z(new_n600));
  NAND3_X1  g414(.A1(new_n598), .A2(G902), .A3(G953), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n554), .A2(new_n597), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n359), .A2(new_n521), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(new_n246), .ZN(G3));
  INV_X1    g421(.A(G472), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n279), .B2(new_n346), .ZN(new_n609));
  INV_X1    g423(.A(new_n280), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n260), .A2(KEYINPUT69), .A3(KEYINPUT31), .ZN(new_n611));
  AOI21_X1  g425(.A(KEYINPUT69), .B1(new_n260), .B2(KEYINPUT31), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n291), .A2(new_n264), .B1(new_n275), .B2(new_n276), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n610), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n609), .A2(new_n615), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n443), .A2(new_n616), .A3(new_n358), .ZN(new_n617));
  INV_X1    g431(.A(new_n444), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n502), .B1(new_n490), .B2(new_n499), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n618), .B1(new_n619), .B2(new_n517), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n549), .A2(new_n622), .A3(new_n550), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n546), .A2(KEYINPUT33), .A3(new_n548), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n623), .A2(G478), .A3(new_n346), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n551), .A2(new_n552), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n597), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n621), .A2(new_n628), .A3(new_n603), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n617), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT94), .B(G104), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT93), .B(KEYINPUT34), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  INV_X1    g448(.A(new_n582), .ZN(new_n635));
  OR3_X1    g449(.A1(new_n591), .A2(KEYINPUT95), .A3(new_n592), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n594), .A2(new_n592), .A3(new_n583), .ZN(new_n637));
  OAI21_X1  g451(.A(KEYINPUT95), .B1(new_n591), .B2(new_n592), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT96), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n636), .A2(new_n638), .A3(KEYINPUT96), .A4(new_n637), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n635), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n621), .A2(new_n603), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n643), .A2(new_n644), .A3(new_n554), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n617), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT35), .B(G107), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  INV_X1    g462(.A(new_n521), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n356), .B1(new_n353), .B2(new_n354), .ZN(new_n650));
  OR2_X1    g464(.A1(new_n336), .A2(KEYINPUT97), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n340), .A2(KEYINPUT36), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n336), .A2(KEYINPUT97), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n652), .B1(new_n651), .B2(new_n653), .ZN(new_n655));
  INV_X1    g469(.A(new_n349), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n650), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n605), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n649), .A2(new_n616), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n660), .B(KEYINPUT37), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G110), .ZN(G12));
  INV_X1    g476(.A(new_n658), .ZN(new_n663));
  AND4_X1   g477(.A1(new_n304), .A2(new_n443), .A3(new_n620), .A4(new_n663), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n599), .B1(new_n601), .B2(G900), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n643), .A2(new_n554), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G128), .ZN(G30));
  XNOR2_X1  g482(.A(new_n520), .B(KEYINPUT38), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n554), .A2(new_n597), .A3(new_n444), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT99), .ZN(new_n671));
  OR3_X1    g485(.A1(new_n670), .A2(new_n663), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n671), .B1(new_n670), .B2(new_n663), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n665), .B(KEYINPUT100), .Z(new_n676));
  XOR2_X1   g490(.A(new_n676), .B(KEYINPUT39), .Z(new_n677));
  NAND2_X1  g491(.A1(new_n443), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT40), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n283), .A2(new_n284), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n247), .B1(new_n297), .B2(new_n239), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT98), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n346), .B1(new_n683), .B2(new_n275), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(G472), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n675), .A2(new_n680), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(new_n206), .ZN(G45));
  INV_X1    g502(.A(new_n665), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n628), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n664), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  NAND2_X1  g506(.A1(new_n428), .A2(new_n346), .ZN(new_n693));
  AOI22_X1  g507(.A1(new_n423), .A2(new_n429), .B1(G469), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n362), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n696), .A2(new_n304), .A3(new_n358), .A4(new_n629), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT41), .B(G113), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT101), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n697), .B(new_n699), .ZN(G15));
  NAND4_X1  g514(.A1(new_n645), .A2(new_n358), .A3(new_n304), .A4(new_n696), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G116), .ZN(G18));
  NAND2_X1  g516(.A1(new_n693), .A2(G469), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n430), .A2(new_n362), .A3(new_n620), .A4(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(KEYINPUT102), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT102), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n694), .A2(new_n706), .A3(new_n362), .A4(new_n620), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n304), .A3(new_n659), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G119), .ZN(G21));
  XNOR2_X1  g524(.A(new_n260), .B(new_n276), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT103), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n299), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g527(.A(KEYINPUT103), .B1(new_n298), .B2(new_n288), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n713), .A2(new_n264), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n610), .B1(new_n711), .B2(new_n715), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n609), .A2(new_n357), .A3(new_n716), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n619), .A2(new_n517), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n670), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n696), .A2(new_n717), .A3(new_n602), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G122), .ZN(G24));
  INV_X1    g535(.A(new_n716), .ZN(new_n722));
  AOI21_X1  g536(.A(G902), .B1(new_n613), .B2(new_n614), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n722), .B(new_n663), .C1(new_n723), .C2(new_n608), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(KEYINPUT104), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n279), .A2(new_n346), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n716), .B1(new_n726), .B2(G472), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT104), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(new_n728), .A3(new_n663), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n708), .A3(new_n690), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G125), .ZN(G27));
  NAND4_X1  g546(.A1(new_n516), .A2(new_n444), .A3(new_n517), .A4(new_n519), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n304), .A2(new_n734), .A3(new_n358), .A4(new_n443), .ZN(new_n735));
  INV_X1    g549(.A(new_n690), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT106), .B1(new_n737), .B2(KEYINPUT42), .ZN(new_n738));
  AOI22_X1  g552(.A1(new_n423), .A2(new_n429), .B1(G469), .B2(new_n441), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n733), .A2(new_n363), .A3(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n740), .A2(new_n358), .A3(new_n304), .A4(new_n690), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT106), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT42), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT105), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n745), .B(new_n743), .C1(new_n735), .C2(new_n736), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n745), .B1(new_n741), .B2(new_n743), .ZN(new_n748));
  OAI22_X1  g562(.A1(new_n738), .A2(new_n744), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G131), .ZN(G33));
  INV_X1    g564(.A(new_n359), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n666), .A3(new_n740), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G134), .ZN(G36));
  OAI21_X1  g567(.A(new_n663), .B1(new_n609), .B2(new_n615), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT43), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n625), .A2(new_n626), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n755), .B1(new_n756), .B2(new_n597), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT108), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT108), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n759), .B(new_n755), .C1(new_n756), .C2(new_n597), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n597), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(KEYINPUT43), .A3(new_n627), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(KEYINPUT109), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT109), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n762), .A2(new_n765), .A3(KEYINPUT43), .A4(new_n627), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n754), .B1(new_n761), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(KEYINPUT44), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n733), .B1(new_n768), .B2(KEYINPUT44), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT45), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n440), .A2(new_n772), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n431), .B(KEYINPUT45), .C1(new_n439), .C2(new_n409), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(G469), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(G469), .A2(G902), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT46), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n775), .A2(KEYINPUT46), .A3(new_n776), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n779), .A2(new_n430), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n362), .ZN(new_n782));
  INV_X1    g596(.A(new_n677), .ZN(new_n783));
  OAI21_X1  g597(.A(KEYINPUT107), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n782), .A2(KEYINPUT107), .A3(new_n783), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n770), .B(new_n771), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G137), .ZN(G39));
  INV_X1    g602(.A(new_n304), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n736), .A2(new_n733), .A3(new_n358), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT110), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n781), .A2(new_n791), .A3(new_n362), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT47), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n791), .B1(new_n781), .B2(new_n362), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n782), .A2(KEYINPUT110), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT47), .B1(new_n797), .B2(new_n792), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n789), .B(new_n790), .C1(new_n796), .C2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G140), .ZN(G42));
  OAI21_X1  g614(.A(new_n794), .B1(new_n793), .B2(new_n795), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n797), .A2(KEYINPUT47), .A3(new_n792), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n694), .A2(new_n363), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n599), .B1(new_n761), .B2(new_n767), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n805), .A2(new_n717), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n804), .A2(new_n806), .A3(new_n734), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n696), .A2(new_n717), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT38), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n520), .B(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n805), .A2(new_n808), .A3(new_n618), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT116), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT50), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT50), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n811), .A2(KEYINPUT116), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n695), .A2(new_n733), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n805), .A2(new_n730), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n358), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n819), .A2(new_n599), .A3(new_n686), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n762), .A3(new_n756), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n807), .A2(new_n816), .A3(new_n818), .A4(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT51), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n806), .A2(new_n708), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n805), .A2(new_n751), .A3(new_n817), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT48), .ZN(new_n827));
  INV_X1    g641(.A(G952), .ZN(new_n828));
  INV_X1    g642(.A(new_n628), .ZN(new_n829));
  AOI211_X1 g643(.A(new_n828), .B(G953), .C1(new_n820), .C2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n831), .B1(new_n822), .B2(new_n823), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n824), .A2(new_n825), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n824), .A2(new_n832), .A3(KEYINPUT117), .A4(new_n825), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n728), .B1(new_n727), .B2(new_n663), .ZN(new_n838));
  NOR4_X1   g652(.A1(new_n609), .A2(new_n716), .A3(new_n658), .A4(KEYINPUT104), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n740), .B(new_n690), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT114), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n730), .A2(KEYINPUT114), .A3(new_n690), .A4(new_n740), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n304), .A2(new_n443), .A3(new_n663), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n733), .A2(new_n554), .A3(new_n689), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n845), .A2(KEYINPUT113), .A3(new_n643), .A4(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT113), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n304), .A2(new_n443), .A3(new_n643), .A4(new_n663), .ZN(new_n849));
  OR3_X1    g663(.A1(new_n733), .A2(new_n554), .A3(new_n689), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n844), .A2(new_n752), .A3(new_n852), .ZN(new_n853));
  NOR4_X1   g667(.A1(new_n609), .A2(new_n615), .A3(new_n357), .A4(new_n603), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n649), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n762), .A2(new_n554), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n660), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n520), .A2(new_n444), .ZN(new_n858));
  AND4_X1   g672(.A1(new_n858), .A2(new_n854), .A3(new_n443), .A4(new_n829), .ZN(new_n859));
  OAI21_X1  g673(.A(KEYINPUT112), .B1(new_n606), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n751), .A2(new_n604), .A3(new_n649), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT112), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n649), .A2(new_n829), .A3(new_n854), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n857), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n853), .A2(KEYINPUT53), .A3(new_n749), .A4(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n709), .A2(new_n701), .A3(new_n697), .A4(new_n720), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n670), .A2(new_n663), .A3(new_n718), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n686), .A2(new_n870), .A3(new_n443), .A4(new_n665), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n667), .A2(new_n691), .A3(new_n731), .A4(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT52), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n872), .A2(KEYINPUT115), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n872), .A2(new_n873), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n736), .B1(new_n725), .B2(new_n729), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n708), .A2(new_n876), .B1(new_n664), .B2(new_n666), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n877), .A2(KEYINPUT52), .A3(new_n691), .A4(new_n871), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT115), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n875), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n867), .A2(new_n869), .A3(new_n874), .A4(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT54), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n868), .A2(KEYINPUT111), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n697), .A2(new_n720), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT111), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n885), .A2(new_n886), .A3(new_n701), .A4(new_n709), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n853), .A2(new_n888), .A3(new_n749), .A4(new_n865), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n875), .A2(new_n878), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n883), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n881), .A2(new_n882), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT53), .B1(new_n889), .B2(new_n891), .ZN(new_n894));
  AND4_X1   g708(.A1(new_n749), .A2(new_n853), .A3(new_n888), .A4(new_n865), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n883), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n880), .A2(new_n874), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n893), .B1(new_n898), .B2(new_n882), .ZN(new_n899));
  OAI22_X1  g713(.A1(new_n837), .A2(new_n899), .B1(G952), .B2(G953), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n669), .A2(new_n597), .A3(new_n756), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT49), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n358), .B(new_n362), .C1(new_n694), .C2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n902), .B2(new_n694), .ZN(new_n904));
  INV_X1    g718(.A(new_n686), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n901), .A2(new_n444), .A3(new_n904), .A4(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n900), .A2(new_n906), .ZN(G75));
  AOI21_X1  g721(.A(KEYINPUT53), .B1(new_n895), .B2(new_n890), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n897), .A2(new_n866), .A3(new_n868), .ZN(new_n909));
  OAI211_X1 g723(.A(G210), .B(G902), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT119), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT56), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n495), .B1(new_n460), .B2(new_n498), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n913), .A2(new_n511), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n914), .A2(new_n499), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT118), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT55), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n910), .A2(new_n911), .A3(new_n912), .A4(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n828), .A2(G953), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT120), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n346), .B1(new_n881), .B2(new_n892), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT56), .B1(new_n922), .B2(G210), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n917), .B1(new_n923), .B2(new_n911), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n911), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n921), .B1(new_n924), .B2(new_n925), .ZN(G51));
  INV_X1    g740(.A(new_n920), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n776), .B(KEYINPUT57), .Z(new_n928));
  INV_X1    g742(.A(new_n893), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n882), .B1(new_n881), .B2(new_n892), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n428), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n922), .A2(G469), .A3(new_n774), .A4(new_n773), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n927), .B1(new_n932), .B2(new_n933), .ZN(G54));
  INV_X1    g748(.A(new_n594), .ZN(new_n935));
  OAI211_X1 g749(.A(KEYINPUT58), .B(G902), .C1(new_n908), .C2(new_n909), .ZN(new_n936));
  INV_X1    g750(.A(G475), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n920), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n922), .A2(KEYINPUT58), .A3(G475), .ZN(new_n940));
  OAI21_X1  g754(.A(KEYINPUT121), .B1(new_n940), .B2(new_n935), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n936), .A2(new_n937), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT121), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n942), .A2(new_n943), .A3(new_n594), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n939), .B1(new_n941), .B2(new_n944), .ZN(G60));
  NAND2_X1  g759(.A1(new_n623), .A2(new_n624), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(G478), .A2(G902), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT59), .Z(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n947), .B1(new_n899), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n947), .A2(new_n950), .ZN(new_n952));
  INV_X1    g766(.A(new_n930), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n952), .B1(new_n953), .B2(new_n893), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n951), .A2(new_n954), .A3(new_n927), .ZN(G63));
  INV_X1    g769(.A(KEYINPUT61), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n881), .A2(new_n892), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n654), .A2(new_n655), .ZN(new_n958));
  XNOR2_X1  g772(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n345), .A2(new_n346), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n957), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n920), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n344), .B1(new_n957), .B2(new_n961), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n956), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n964), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n966), .A2(KEYINPUT61), .A3(new_n920), .A4(new_n962), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n965), .A2(new_n967), .ZN(G66));
  AOI21_X1  g782(.A(new_n241), .B1(new_n600), .B2(new_n466), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n888), .A2(new_n865), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n969), .B1(new_n970), .B2(new_n241), .ZN(new_n971));
  INV_X1    g785(.A(G898), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n913), .B1(new_n972), .B2(G953), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT123), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n971), .B(new_n974), .ZN(G69));
  NOR2_X1   g789(.A1(new_n678), .A2(new_n733), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n856), .A2(new_n628), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n751), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n687), .A2(new_n691), .A3(new_n877), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT62), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n667), .A2(new_n691), .A3(new_n731), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n983), .A2(KEYINPUT62), .A3(new_n687), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n979), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n799), .A2(new_n787), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n250), .A2(new_n255), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(new_n587), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n751), .B(new_n719), .C1(new_n785), .C2(new_n786), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n799), .A2(new_n752), .A3(new_n787), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n749), .A2(new_n983), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n241), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n989), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(G953), .B1(new_n990), .B2(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(G900), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(G953), .B1(new_n407), .B2(new_n998), .ZN(new_n1000));
  OAI22_X1  g814(.A1(new_n997), .A2(new_n999), .B1(KEYINPUT124), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(KEYINPUT124), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1001), .B(new_n1002), .ZN(G72));
  INV_X1    g817(.A(new_n286), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n992), .A2(new_n970), .A3(new_n993), .ZN(new_n1005));
  NAND2_X1  g819(.A1(G472), .A2(G902), .ZN(new_n1006));
  XOR2_X1   g820(.A(new_n1006), .B(KEYINPUT63), .Z(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(new_n1008));
  OAI211_X1 g822(.A(new_n264), .B(new_n1004), .C1(new_n1005), .C2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n920), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT126), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n985), .A2(new_n888), .A3(new_n865), .A4(new_n986), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n264), .B1(new_n1013), .B2(new_n1007), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT125), .ZN(new_n1015));
  AND3_X1   g829(.A1(new_n1014), .A2(new_n1015), .A3(new_n286), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1015), .B1(new_n1014), .B2(new_n286), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n287), .B(KEYINPUT127), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1007), .B1(new_n1018), .B2(new_n275), .ZN(new_n1019));
  OAI22_X1  g833(.A1(new_n1016), .A2(new_n1017), .B1(new_n898), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n1012), .A2(new_n1020), .ZN(G57));
endmodule


