

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580;

  XOR2_X1 U322 ( .A(n380), .B(n379), .Z(n514) );
  XOR2_X1 U323 ( .A(n442), .B(n441), .Z(n290) );
  XOR2_X1 U324 ( .A(n437), .B(n436), .Z(n291) );
  INV_X1 U325 ( .A(G197GAT), .ZN(n353) );
  XNOR2_X1 U326 ( .A(n354), .B(n353), .ZN(n356) );
  XNOR2_X1 U327 ( .A(n443), .B(n290), .ZN(n444) );
  XNOR2_X1 U328 ( .A(n356), .B(n355), .ZN(n373) );
  XNOR2_X1 U329 ( .A(n445), .B(n444), .ZN(n446) );
  INV_X1 U330 ( .A(G190GAT), .ZN(n468) );
  NOR2_X1 U331 ( .A1(n523), .A2(n467), .ZN(n561) );
  XOR2_X1 U332 ( .A(n570), .B(KEYINPUT41), .Z(n556) );
  INV_X1 U333 ( .A(G43GAT), .ZN(n449) );
  XNOR2_X1 U334 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U335 ( .A(n449), .B(KEYINPUT40), .ZN(n450) );
  XNOR2_X1 U336 ( .A(n471), .B(n470), .ZN(G1351GAT) );
  XNOR2_X1 U337 ( .A(n451), .B(n450), .ZN(G1330GAT) );
  XOR2_X1 U338 ( .A(G120GAT), .B(G71GAT), .Z(n437) );
  XOR2_X1 U339 ( .A(G99GAT), .B(G15GAT), .Z(n293) );
  XNOR2_X1 U340 ( .A(G169GAT), .B(G43GAT), .ZN(n292) );
  XNOR2_X1 U341 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U342 ( .A(n437), .B(n294), .Z(n296) );
  NAND2_X1 U343 ( .A1(G227GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U344 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U345 ( .A(G176GAT), .B(KEYINPUT20), .Z(n298) );
  XNOR2_X1 U346 ( .A(KEYINPUT87), .B(KEYINPUT85), .ZN(n297) );
  XNOR2_X1 U347 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U348 ( .A(n300), .B(n299), .Z(n309) );
  XNOR2_X1 U349 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n301), .B(KEYINPUT86), .ZN(n302) );
  XOR2_X1 U351 ( .A(n302), .B(KEYINPUT18), .Z(n304) );
  XNOR2_X1 U352 ( .A(G183GAT), .B(G190GAT), .ZN(n303) );
  XNOR2_X1 U353 ( .A(n304), .B(n303), .ZN(n380) );
  XOR2_X1 U354 ( .A(KEYINPUT84), .B(G134GAT), .Z(n306) );
  XNOR2_X1 U355 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n305) );
  XNOR2_X1 U356 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U357 ( .A(G113GAT), .B(n307), .ZN(n345) );
  XOR2_X1 U358 ( .A(n380), .B(n345), .Z(n308) );
  XOR2_X1 U359 ( .A(n309), .B(n308), .Z(n484) );
  INV_X1 U360 ( .A(n484), .ZN(n523) );
  XOR2_X1 U361 ( .A(G155GAT), .B(G78GAT), .Z(n311) );
  XNOR2_X1 U362 ( .A(G22GAT), .B(G211GAT), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U364 ( .A(G71GAT), .B(G127GAT), .Z(n313) );
  XNOR2_X1 U365 ( .A(G8GAT), .B(G183GAT), .ZN(n312) );
  XNOR2_X1 U366 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U367 ( .A(n315), .B(n314), .Z(n320) );
  XOR2_X1 U368 ( .A(KEYINPUT81), .B(KEYINPUT83), .Z(n317) );
  NAND2_X1 U369 ( .A1(G231GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U370 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U371 ( .A(KEYINPUT82), .B(n318), .ZN(n319) );
  XNOR2_X1 U372 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U373 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n322) );
  XNOR2_X1 U374 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U376 ( .A(n324), .B(n323), .Z(n328) );
  XNOR2_X1 U377 ( .A(G15GAT), .B(G1GAT), .ZN(n325) );
  XNOR2_X1 U378 ( .A(n325), .B(KEYINPUT68), .ZN(n426) );
  XNOR2_X1 U379 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n326), .B(KEYINPUT13), .ZN(n432) );
  XNOR2_X1 U381 ( .A(n426), .B(n432), .ZN(n327) );
  XOR2_X1 U382 ( .A(n328), .B(n327), .Z(n573) );
  INV_X1 U383 ( .A(n573), .ZN(n472) );
  XOR2_X1 U384 ( .A(G155GAT), .B(KEYINPUT2), .Z(n330) );
  XNOR2_X1 U385 ( .A(G162GAT), .B(KEYINPUT3), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n330), .B(n329), .ZN(n367) );
  XOR2_X1 U387 ( .A(G85GAT), .B(n367), .Z(n332) );
  NAND2_X1 U388 ( .A1(G225GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U389 ( .A(n332), .B(n331), .ZN(n352) );
  XOR2_X1 U390 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n334) );
  XNOR2_X1 U391 ( .A(KEYINPUT94), .B(KEYINPUT96), .ZN(n333) );
  XNOR2_X1 U392 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U393 ( .A(KEYINPUT95), .B(G148GAT), .Z(n336) );
  XNOR2_X1 U394 ( .A(G141GAT), .B(G120GAT), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n338), .B(n337), .ZN(n349) );
  XOR2_X1 U397 ( .A(G57GAT), .B(KEYINPUT97), .Z(n340) );
  XNOR2_X1 U398 ( .A(KEYINPUT92), .B(KEYINPUT98), .ZN(n339) );
  XNOR2_X1 U399 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U400 ( .A(KEYINPUT1), .B(KEYINPUT93), .Z(n342) );
  XNOR2_X1 U401 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n341) );
  XNOR2_X1 U402 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U403 ( .A(n344), .B(n343), .ZN(n347) );
  INV_X1 U404 ( .A(n345), .ZN(n346) );
  XOR2_X1 U405 ( .A(n347), .B(n346), .Z(n348) );
  XNOR2_X1 U406 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U407 ( .A(G29GAT), .B(n350), .Z(n351) );
  XOR2_X1 U408 ( .A(n352), .B(n351), .Z(n478) );
  XNOR2_X1 U409 ( .A(KEYINPUT90), .B(G211GAT), .ZN(n354) );
  XOR2_X1 U410 ( .A(KEYINPUT21), .B(G218GAT), .Z(n355) );
  XOR2_X1 U411 ( .A(G141GAT), .B(G22GAT), .Z(n429) );
  XOR2_X1 U412 ( .A(G204GAT), .B(KEYINPUT89), .Z(n358) );
  XNOR2_X1 U413 ( .A(G50GAT), .B(KEYINPUT91), .ZN(n357) );
  XNOR2_X1 U414 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U415 ( .A(n429), .B(n359), .Z(n361) );
  NAND2_X1 U416 ( .A1(G228GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n361), .B(n360), .ZN(n365) );
  XOR2_X1 U418 ( .A(KEYINPUT88), .B(KEYINPUT22), .Z(n363) );
  XNOR2_X1 U419 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n362) );
  XNOR2_X1 U420 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U421 ( .A(n365), .B(n364), .Z(n369) );
  XNOR2_X1 U422 ( .A(G106GAT), .B(G78GAT), .ZN(n366) );
  XNOR2_X1 U423 ( .A(n366), .B(G148GAT), .ZN(n440) );
  XNOR2_X1 U424 ( .A(n440), .B(n367), .ZN(n368) );
  XNOR2_X1 U425 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U426 ( .A(n373), .B(n370), .ZN(n465) );
  XOR2_X1 U427 ( .A(G169GAT), .B(G8GAT), .Z(n428) );
  XOR2_X1 U428 ( .A(G64GAT), .B(G92GAT), .Z(n372) );
  XNOR2_X1 U429 ( .A(G176GAT), .B(G204GAT), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n372), .B(n371), .ZN(n433) );
  XOR2_X1 U431 ( .A(n433), .B(KEYINPUT99), .Z(n375) );
  XNOR2_X1 U432 ( .A(G36GAT), .B(n373), .ZN(n374) );
  XNOR2_X1 U433 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U434 ( .A(n428), .B(n376), .Z(n378) );
  NAND2_X1 U435 ( .A1(G226GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U436 ( .A(n378), .B(n377), .ZN(n379) );
  NOR2_X1 U437 ( .A1(n523), .A2(n514), .ZN(n381) );
  NOR2_X1 U438 ( .A1(n465), .A2(n381), .ZN(n382) );
  XOR2_X1 U439 ( .A(KEYINPUT25), .B(n382), .Z(n386) );
  NAND2_X1 U440 ( .A1(n465), .A2(n523), .ZN(n383) );
  XNOR2_X1 U441 ( .A(n383), .B(KEYINPUT26), .ZN(n384) );
  XNOR2_X1 U442 ( .A(KEYINPUT102), .B(n384), .ZN(n563) );
  XNOR2_X1 U443 ( .A(KEYINPUT27), .B(n514), .ZN(n388) );
  NOR2_X1 U444 ( .A1(n563), .A2(n388), .ZN(n385) );
  NOR2_X1 U445 ( .A1(n386), .A2(n385), .ZN(n387) );
  NOR2_X1 U446 ( .A1(n478), .A2(n387), .ZN(n393) );
  XOR2_X1 U447 ( .A(KEYINPUT28), .B(n465), .Z(n518) );
  INV_X1 U448 ( .A(n518), .ZN(n526) );
  INV_X1 U449 ( .A(n478), .ZN(n512) );
  NOR2_X1 U450 ( .A1(n388), .A2(n512), .ZN(n389) );
  XNOR2_X1 U451 ( .A(n389), .B(KEYINPUT100), .ZN(n521) );
  NAND2_X1 U452 ( .A1(n521), .A2(n523), .ZN(n390) );
  NOR2_X1 U453 ( .A1(n526), .A2(n390), .ZN(n391) );
  XOR2_X1 U454 ( .A(KEYINPUT101), .B(n391), .Z(n392) );
  NOR2_X1 U455 ( .A1(n393), .A2(n392), .ZN(n475) );
  XOR2_X1 U456 ( .A(KEYINPUT78), .B(KEYINPUT77), .Z(n395) );
  XNOR2_X1 U457 ( .A(KEYINPUT9), .B(KEYINPUT11), .ZN(n394) );
  XNOR2_X1 U458 ( .A(n395), .B(n394), .ZN(n409) );
  XOR2_X1 U459 ( .A(KEYINPUT10), .B(KEYINPUT79), .Z(n397) );
  XNOR2_X1 U460 ( .A(G190GAT), .B(G106GAT), .ZN(n396) );
  XNOR2_X1 U461 ( .A(n397), .B(n396), .ZN(n401) );
  XOR2_X1 U462 ( .A(KEYINPUT64), .B(G92GAT), .Z(n399) );
  XNOR2_X1 U463 ( .A(G134GAT), .B(G162GAT), .ZN(n398) );
  XNOR2_X1 U464 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U465 ( .A(n401), .B(n400), .Z(n407) );
  XNOR2_X1 U466 ( .A(G99GAT), .B(G85GAT), .ZN(n402) );
  XNOR2_X1 U467 ( .A(n402), .B(KEYINPUT73), .ZN(n439) );
  XOR2_X1 U468 ( .A(KEYINPUT80), .B(n439), .Z(n404) );
  NAND2_X1 U469 ( .A1(G232GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U470 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U471 ( .A(G218GAT), .B(n405), .ZN(n406) );
  XNOR2_X1 U472 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U473 ( .A(n409), .B(n408), .ZN(n414) );
  XNOR2_X1 U474 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n410) );
  XNOR2_X1 U475 ( .A(n410), .B(G29GAT), .ZN(n411) );
  XOR2_X1 U476 ( .A(n411), .B(KEYINPUT8), .Z(n413) );
  XNOR2_X1 U477 ( .A(G43GAT), .B(G50GAT), .ZN(n412) );
  XOR2_X1 U478 ( .A(n413), .B(n412), .Z(n423) );
  XNOR2_X1 U479 ( .A(n414), .B(n423), .ZN(n550) );
  XOR2_X1 U480 ( .A(KEYINPUT36), .B(n550), .Z(n578) );
  NOR2_X1 U481 ( .A1(n475), .A2(n578), .ZN(n415) );
  NAND2_X1 U482 ( .A1(n472), .A2(n415), .ZN(n416) );
  XNOR2_X1 U483 ( .A(KEYINPUT37), .B(n416), .ZN(n511) );
  XOR2_X1 U484 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n418) );
  NAND2_X1 U485 ( .A1(G229GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U486 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U487 ( .A(n419), .B(KEYINPUT66), .Z(n425) );
  XOR2_X1 U488 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n421) );
  XNOR2_X1 U489 ( .A(G197GAT), .B(G113GAT), .ZN(n420) );
  XNOR2_X1 U490 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U491 ( .A(n423), .B(n422), .Z(n424) );
  XNOR2_X1 U492 ( .A(n425), .B(n424), .ZN(n427) );
  XOR2_X1 U493 ( .A(n427), .B(n426), .Z(n431) );
  XNOR2_X1 U494 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U495 ( .A(n431), .B(n430), .ZN(n565) );
  XNOR2_X1 U496 ( .A(n565), .B(KEYINPUT69), .ZN(n527) );
  XNOR2_X1 U497 ( .A(n433), .B(n432), .ZN(n447) );
  XOR2_X1 U498 ( .A(KEYINPUT32), .B(KEYINPUT76), .Z(n435) );
  XNOR2_X1 U499 ( .A(KEYINPUT75), .B(KEYINPUT71), .ZN(n434) );
  XNOR2_X1 U500 ( .A(n435), .B(n434), .ZN(n436) );
  NAND2_X1 U501 ( .A1(G230GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U502 ( .A(n291), .B(n438), .ZN(n445) );
  XNOR2_X1 U503 ( .A(n440), .B(n439), .ZN(n443) );
  XOR2_X1 U504 ( .A(KEYINPUT72), .B(KEYINPUT33), .Z(n442) );
  XNOR2_X1 U505 ( .A(KEYINPUT74), .B(KEYINPUT31), .ZN(n441) );
  XOR2_X1 U506 ( .A(n447), .B(n446), .Z(n570) );
  NOR2_X1 U507 ( .A1(n527), .A2(n570), .ZN(n476) );
  NAND2_X1 U508 ( .A1(n511), .A2(n476), .ZN(n448) );
  XNOR2_X1 U509 ( .A(KEYINPUT38), .B(n448), .ZN(n494) );
  NOR2_X1 U510 ( .A1(n523), .A2(n494), .ZN(n451) );
  NAND2_X1 U511 ( .A1(n565), .A2(n556), .ZN(n452) );
  XNOR2_X1 U512 ( .A(KEYINPUT46), .B(n452), .ZN(n453) );
  NAND2_X1 U513 ( .A1(n453), .A2(n472), .ZN(n454) );
  NOR2_X1 U514 ( .A1(n550), .A2(n454), .ZN(n455) );
  XNOR2_X1 U515 ( .A(n455), .B(KEYINPUT47), .ZN(n460) );
  NOR2_X1 U516 ( .A1(n472), .A2(n578), .ZN(n456) );
  XOR2_X1 U517 ( .A(KEYINPUT45), .B(n456), .Z(n457) );
  NOR2_X1 U518 ( .A1(n570), .A2(n457), .ZN(n458) );
  NAND2_X1 U519 ( .A1(n458), .A2(n527), .ZN(n459) );
  NAND2_X1 U520 ( .A1(n460), .A2(n459), .ZN(n461) );
  XNOR2_X1 U521 ( .A(KEYINPUT48), .B(n461), .ZN(n522) );
  INV_X1 U522 ( .A(n514), .ZN(n482) );
  NAND2_X1 U523 ( .A1(n522), .A2(n482), .ZN(n463) );
  XOR2_X1 U524 ( .A(KEYINPUT54), .B(KEYINPUT122), .Z(n462) );
  XNOR2_X1 U525 ( .A(n463), .B(n462), .ZN(n464) );
  NAND2_X1 U526 ( .A1(n512), .A2(n464), .ZN(n564) );
  NOR2_X1 U527 ( .A1(n465), .A2(n564), .ZN(n466) );
  XNOR2_X1 U528 ( .A(n466), .B(KEYINPUT55), .ZN(n467) );
  NAND2_X1 U529 ( .A1(n561), .A2(n550), .ZN(n471) );
  XOR2_X1 U530 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n469) );
  XOR2_X1 U531 ( .A(KEYINPUT34), .B(KEYINPUT104), .Z(n480) );
  NOR2_X1 U532 ( .A1(n472), .A2(n550), .ZN(n473) );
  XOR2_X1 U533 ( .A(KEYINPUT16), .B(n473), .Z(n474) );
  NOR2_X1 U534 ( .A1(n475), .A2(n474), .ZN(n498) );
  NAND2_X1 U535 ( .A1(n476), .A2(n498), .ZN(n477) );
  XNOR2_X1 U536 ( .A(KEYINPUT103), .B(n477), .ZN(n488) );
  NAND2_X1 U537 ( .A1(n488), .A2(n478), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U539 ( .A(G1GAT), .B(n481), .Z(G1324GAT) );
  NAND2_X1 U540 ( .A1(n482), .A2(n488), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n483), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U542 ( .A(KEYINPUT105), .B(KEYINPUT35), .Z(n486) );
  NAND2_X1 U543 ( .A1(n488), .A2(n484), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U545 ( .A(G15GAT), .B(n487), .Z(G1326GAT) );
  NAND2_X1 U546 ( .A1(n488), .A2(n526), .ZN(n489) );
  XNOR2_X1 U547 ( .A(n489), .B(G22GAT), .ZN(G1327GAT) );
  XNOR2_X1 U548 ( .A(KEYINPUT39), .B(KEYINPUT106), .ZN(n491) );
  NOR2_X1 U549 ( .A1(n512), .A2(n494), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U551 ( .A(G29GAT), .B(n492), .ZN(G1328GAT) );
  NOR2_X1 U552 ( .A1(n514), .A2(n494), .ZN(n493) );
  XOR2_X1 U553 ( .A(G36GAT), .B(n493), .Z(G1329GAT) );
  NOR2_X1 U554 ( .A1(n494), .A2(n518), .ZN(n496) );
  XNOR2_X1 U555 ( .A(G50GAT), .B(KEYINPUT107), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n496), .B(n495), .ZN(G1331GAT) );
  INV_X1 U557 ( .A(n556), .ZN(n497) );
  NOR2_X1 U558 ( .A1(n565), .A2(n497), .ZN(n510) );
  NAND2_X1 U559 ( .A1(n510), .A2(n498), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n499), .B(KEYINPUT108), .ZN(n506) );
  NOR2_X1 U561 ( .A1(n512), .A2(n506), .ZN(n502) );
  XNOR2_X1 U562 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n500), .B(KEYINPUT109), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(G1332GAT) );
  NOR2_X1 U565 ( .A1(n514), .A2(n506), .ZN(n503) );
  XOR2_X1 U566 ( .A(G64GAT), .B(n503), .Z(G1333GAT) );
  NOR2_X1 U567 ( .A1(n523), .A2(n506), .ZN(n504) );
  XOR2_X1 U568 ( .A(KEYINPUT110), .B(n504), .Z(n505) );
  XNOR2_X1 U569 ( .A(G71GAT), .B(n505), .ZN(G1334GAT) );
  NOR2_X1 U570 ( .A1(n506), .A2(n518), .ZN(n508) );
  XNOR2_X1 U571 ( .A(KEYINPUT43), .B(KEYINPUT111), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U573 ( .A(G78GAT), .B(n509), .Z(G1335GAT) );
  NAND2_X1 U574 ( .A1(n511), .A2(n510), .ZN(n517) );
  NOR2_X1 U575 ( .A1(n512), .A2(n517), .ZN(n513) );
  XOR2_X1 U576 ( .A(G85GAT), .B(n513), .Z(G1336GAT) );
  NOR2_X1 U577 ( .A1(n514), .A2(n517), .ZN(n515) );
  XOR2_X1 U578 ( .A(G92GAT), .B(n515), .Z(G1337GAT) );
  NOR2_X1 U579 ( .A1(n523), .A2(n517), .ZN(n516) );
  XOR2_X1 U580 ( .A(G99GAT), .B(n516), .Z(G1338GAT) );
  NOR2_X1 U581 ( .A1(n518), .A2(n517), .ZN(n519) );
  XOR2_X1 U582 ( .A(KEYINPUT44), .B(n519), .Z(n520) );
  XNOR2_X1 U583 ( .A(G106GAT), .B(n520), .ZN(G1339GAT) );
  XOR2_X1 U584 ( .A(G113GAT), .B(KEYINPUT113), .Z(n529) );
  NAND2_X1 U585 ( .A1(n522), .A2(n521), .ZN(n540) );
  NOR2_X1 U586 ( .A1(n523), .A2(n540), .ZN(n524) );
  XOR2_X1 U587 ( .A(KEYINPUT112), .B(n524), .Z(n525) );
  NOR2_X1 U588 ( .A1(n526), .A2(n525), .ZN(n535) );
  INV_X1 U589 ( .A(n527), .ZN(n554) );
  NAND2_X1 U590 ( .A1(n535), .A2(n554), .ZN(n528) );
  XNOR2_X1 U591 ( .A(n529), .B(n528), .ZN(G1340GAT) );
  XOR2_X1 U592 ( .A(G120GAT), .B(KEYINPUT49), .Z(n531) );
  NAND2_X1 U593 ( .A1(n535), .A2(n556), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT114), .B(KEYINPUT50), .Z(n533) );
  NAND2_X1 U596 ( .A1(n535), .A2(n573), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U598 ( .A(G127GAT), .B(n534), .Z(G1342GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n537) );
  NAND2_X1 U600 ( .A1(n535), .A2(n550), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n537), .B(n536), .ZN(n539) );
  XOR2_X1 U602 ( .A(G134GAT), .B(KEYINPUT115), .Z(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(G1343GAT) );
  XOR2_X1 U604 ( .A(G141GAT), .B(KEYINPUT117), .Z(n542) );
  NOR2_X1 U605 ( .A1(n540), .A2(n563), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n551), .A2(n565), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(G1344GAT) );
  XNOR2_X1 U608 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n546) );
  XOR2_X1 U609 ( .A(KEYINPUT52), .B(KEYINPUT118), .Z(n544) );
  NAND2_X1 U610 ( .A1(n551), .A2(n556), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(G1345GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n548) );
  NAND2_X1 U614 ( .A1(n551), .A2(n573), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(G155GAT), .B(n549), .ZN(G1346GAT) );
  XOR2_X1 U617 ( .A(G162GAT), .B(KEYINPUT121), .Z(n553) );
  NAND2_X1 U618 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1347GAT) );
  NAND2_X1 U620 ( .A1(n561), .A2(n554), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n558) );
  NAND2_X1 U623 ( .A1(n561), .A2(n556), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(n560) );
  XOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT56), .Z(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1349GAT) );
  NAND2_X1 U627 ( .A1(n573), .A2(n561), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U629 ( .A(G197GAT), .B(KEYINPUT125), .Z(n567) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n576) );
  NAND2_X1 U631 ( .A1(n576), .A2(n565), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .Z(n572) );
  NAND2_X1 U636 ( .A1(n576), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1353GAT) );
  NAND2_X1 U638 ( .A1(n573), .A2(n576), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(KEYINPUT126), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G211GAT), .B(n575), .ZN(G1354GAT) );
  INV_X1 U641 ( .A(n576), .ZN(n577) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U643 ( .A(KEYINPUT62), .B(n579), .Z(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(n580), .ZN(G1355GAT) );
endmodule

