//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 1 0 0 0 0 1 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 0 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n575, new_n577, new_n578, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n641, new_n644, new_n646, new_n647,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1217, new_n1218;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  XOR2_X1   g011(.A(new_n436), .B(KEYINPUT64), .Z(G220));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G96), .Z(G221));
  XNOR2_X1  g013(.A(KEYINPUT66), .B(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n452), .A2(G2106), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT68), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(new_n454), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT69), .Z(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G137), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n463), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT72), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT72), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n470), .A2(new_n473), .A3(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n477));
  AND3_X1   g052(.A1(new_n464), .A2(new_n466), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n477), .B1(new_n464), .B2(new_n466), .ZN(new_n479));
  OAI21_X1  g054(.A(G125), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(KEYINPUT71), .ZN(new_n481));
  NAND2_X1  g056(.A1(G113), .A2(G2104), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT71), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G125), .C1(new_n478), .C2(new_n479), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n476), .B1(new_n485), .B2(G2105), .ZN(G160));
  NAND2_X1  g061(.A1(new_n468), .A2(G136), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT73), .ZN(new_n488));
  INV_X1    g063(.A(G2105), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n467), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  NOR2_X1   g066(.A1(G100), .A2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(new_n489), .B2(G112), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OR2_X1    g069(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  OAI211_X1 g071(.A(G138), .B(new_n489), .C1(new_n478), .C2(new_n479), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n464), .A2(new_n466), .A3(G126), .ZN(new_n500));
  NAND2_X1  g075(.A1(G114), .A2(G2104), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n489), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n470), .A2(G102), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT74), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT4), .A2(G138), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n468), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT74), .ZN(new_n508));
  INV_X1    g083(.A(new_n501), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT3), .B(G2104), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(G126), .ZN(new_n511));
  OAI211_X1 g086(.A(new_n508), .B(new_n503), .C1(new_n511), .C2(new_n489), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n499), .A2(new_n505), .A3(new_n507), .A4(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(G164));
  AND2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  OAI21_X1  g091(.A(G543), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n521), .A2(KEYINPUT5), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT5), .ZN(new_n523));
  OAI21_X1  g098(.A(KEYINPUT75), .B1(new_n523), .B2(G543), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT75), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n525), .A2(new_n521), .A3(KEYINPUT5), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n522), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n527), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT6), .B(G651), .ZN(new_n529));
  INV_X1    g104(.A(new_n522), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n525), .B1(KEYINPUT5), .B2(new_n521), .ZN(new_n531));
  NOR3_X1   g106(.A1(new_n523), .A2(KEYINPUT75), .A3(G543), .ZN(new_n532));
  OAI211_X1 g107(.A(new_n529), .B(new_n530), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n527), .A2(KEYINPUT76), .A3(new_n529), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G88), .ZN(new_n538));
  OAI221_X1 g113(.A(new_n519), .B1(new_n520), .B2(new_n528), .C1(new_n537), .C2(new_n538), .ZN(G303));
  INV_X1    g114(.A(G303), .ZN(G166));
  AND3_X1   g115(.A1(new_n535), .A2(G89), .A3(new_n536), .ZN(new_n541));
  AOI21_X1  g116(.A(KEYINPUT77), .B1(new_n529), .B2(G543), .ZN(new_n542));
  OAI211_X1 g117(.A(KEYINPUT77), .B(G543), .C1(new_n515), .C2(new_n516), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g119(.A(G51), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n527), .A2(G63), .A3(G651), .ZN(new_n546));
  NAND3_X1  g121(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n547));
  XOR2_X1   g122(.A(new_n547), .B(KEYINPUT7), .Z(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n545), .A2(new_n546), .A3(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n541), .A2(new_n550), .ZN(G168));
  AOI22_X1  g126(.A1(new_n527), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(new_n520), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n535), .A2(G90), .A3(new_n536), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT79), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT77), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n517), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(new_n543), .ZN(new_n558));
  XOR2_X1   g133(.A(KEYINPUT78), .B(G52), .Z(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AND3_X1   g135(.A1(new_n554), .A2(new_n555), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n555), .B1(new_n554), .B2(new_n560), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n553), .B1(new_n561), .B2(new_n562), .ZN(G301));
  INV_X1    g138(.A(G301), .ZN(G171));
  NAND3_X1  g139(.A1(new_n535), .A2(G81), .A3(new_n536), .ZN(new_n565));
  NAND2_X1  g140(.A1(G68), .A2(G543), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n567));
  INV_X1    g142(.A(G56), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G651), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n558), .A2(G43), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n565), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G860), .ZN(G153));
  AND3_X1   g149(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G36), .ZN(G176));
  NAND2_X1  g151(.A1(G1), .A2(G3), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT8), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n575), .A2(new_n578), .ZN(G188));
  INV_X1    g154(.A(G91), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT80), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n533), .A2(new_n534), .ZN(new_n582));
  AOI21_X1  g157(.A(KEYINPUT76), .B1(new_n527), .B2(new_n529), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n535), .A2(KEYINPUT80), .A3(new_n536), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n580), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AND2_X1   g161(.A1(G78), .A2(G543), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(new_n527), .B2(G65), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT81), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI211_X1 g165(.A(KEYINPUT81), .B(new_n587), .C1(new_n527), .C2(G65), .ZN(new_n591));
  NOR3_X1   g166(.A1(new_n590), .A2(new_n591), .A3(new_n520), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n518), .A2(G53), .ZN(new_n593));
  XOR2_X1   g168(.A(new_n593), .B(KEYINPUT9), .Z(new_n594));
  NOR3_X1   g169(.A1(new_n586), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G299));
  OAI21_X1  g171(.A(KEYINPUT82), .B1(new_n541), .B2(new_n550), .ZN(new_n597));
  INV_X1    g172(.A(G51), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(new_n557), .B2(new_n543), .ZN(new_n599));
  NAND2_X1  g174(.A1(G63), .A2(G651), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n567), .A2(new_n600), .ZN(new_n601));
  NOR3_X1   g176(.A1(new_n599), .A2(new_n601), .A3(new_n548), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT82), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n535), .A2(G89), .A3(new_n536), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n597), .A2(new_n605), .ZN(G286));
  NOR3_X1   g181(.A1(new_n582), .A2(new_n583), .A3(new_n581), .ZN(new_n607));
  AOI21_X1  g182(.A(KEYINPUT80), .B1(new_n535), .B2(new_n536), .ZN(new_n608));
  OAI21_X1  g183(.A(G87), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(G651), .B1(new_n527), .B2(G74), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n518), .A2(G49), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(G288));
  NAND2_X1  g187(.A1(new_n584), .A2(new_n585), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G86), .ZN(new_n614));
  NAND2_X1  g189(.A1(G73), .A2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G61), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n567), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n617), .A2(G651), .B1(G48), .B2(new_n518), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n614), .A2(new_n618), .ZN(G305));
  INV_X1    g194(.A(new_n537), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n620), .A2(G85), .B1(G47), .B2(new_n558), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n527), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT83), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n624), .A2(new_n625), .A3(G651), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n621), .A2(new_n626), .ZN(G290));
  NAND2_X1  g202(.A1(G301), .A2(G868), .ZN(new_n628));
  OAI21_X1  g203(.A(G92), .B1(new_n607), .B2(new_n608), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(KEYINPUT10), .ZN(new_n630));
  AOI22_X1  g205(.A1(new_n527), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT84), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  AOI22_X1  g208(.A1(new_n633), .A2(G651), .B1(G54), .B2(new_n558), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT10), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n613), .A2(new_n635), .A3(G92), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n630), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n628), .B1(new_n638), .B2(G868), .ZN(G284));
  OAI21_X1  g214(.A(new_n628), .B1(new_n638), .B2(G868), .ZN(G321));
  NAND2_X1  g215(.A1(G286), .A2(G868), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(G868), .B2(new_n595), .ZN(G297));
  OAI21_X1  g217(.A(new_n641), .B1(G868), .B2(new_n595), .ZN(G280));
  INV_X1    g218(.A(G559), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n638), .B1(new_n644), .B2(G860), .ZN(G148));
  NAND2_X1  g220(.A1(new_n638), .A2(new_n644), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(G868), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(G868), .B2(new_n573), .ZN(G323));
  XNOR2_X1  g223(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g224(.A(new_n470), .B1(new_n478), .B2(new_n479), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT12), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT13), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2100), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n490), .A2(G123), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n468), .A2(G135), .ZN(new_n655));
  NOR2_X1   g230(.A1(G99), .A2(G2105), .ZN(new_n656));
  OAI21_X1  g231(.A(G2104), .B1(new_n489), .B2(G111), .ZN(new_n657));
  OAI211_X1 g232(.A(new_n654), .B(new_n655), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(G2096), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n653), .A2(new_n660), .ZN(G156));
  XOR2_X1   g236(.A(KEYINPUT15), .B(G2435), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2438), .ZN(new_n663));
  XOR2_X1   g238(.A(G2427), .B(G2430), .Z(new_n664));
  OAI21_X1  g239(.A(KEYINPUT14), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT86), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n664), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT16), .Z(new_n669));
  XNOR2_X1  g244(.A(G2451), .B(G2454), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT85), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2443), .B(G2446), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1341), .B(G1348), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n669), .B(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(G14), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT87), .Z(G401));
  XOR2_X1   g254(.A(G2084), .B(G2090), .Z(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G2067), .B(G2678), .Z(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G2072), .B(G2078), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n681), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT88), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n684), .B(KEYINPUT89), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT17), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n686), .B1(new_n688), .B2(new_n682), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n688), .A2(new_n682), .A3(new_n680), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n683), .A2(new_n684), .A3(new_n680), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT18), .Z(new_n692));
  NAND3_X1  g267(.A1(new_n689), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(new_n659), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G2100), .ZN(G227));
  XOR2_X1   g270(.A(G1956), .B(G2474), .Z(new_n696));
  XOR2_X1   g271(.A(G1961), .B(G1966), .Z(new_n697));
  NOR2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1971), .B(G1976), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT19), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n696), .A2(new_n697), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n698), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n700), .A2(KEYINPUT92), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n700), .A2(new_n701), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT90), .B(KEYINPUT91), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT20), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n706), .B(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT21), .B(G1986), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1991), .B(G1996), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT22), .B(G1981), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n714), .B(new_n715), .Z(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(G229));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G4), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(new_n638), .B2(new_n718), .ZN(new_n720));
  INV_X1    g295(.A(G1348), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT95), .B(G16), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G20), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT103), .B(KEYINPUT23), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G299), .B2(G16), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G1956), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n723), .A2(G19), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n573), .B2(new_n723), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT28), .ZN(new_n732));
  INV_X1    g307(.A(G26), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(G29), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(G29), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n490), .A2(G128), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n468), .A2(G140), .ZN(new_n737));
  OR2_X1    g312(.A1(G104), .A2(G2105), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n738), .B(G2104), .C1(G116), .C2(new_n489), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n736), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n735), .B1(new_n740), .B2(G29), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n734), .B1(new_n741), .B2(new_n732), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n731), .A2(G1341), .B1(G2067), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n722), .A2(new_n729), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(G301), .A2(G16), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n718), .A2(G5), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(KEYINPUT100), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT100), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n745), .A2(new_n749), .A3(new_n746), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G1961), .ZN(new_n752));
  INV_X1    g327(.A(G1961), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n748), .A2(new_n753), .A3(new_n750), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(G29), .A2(G32), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n468), .A2(G141), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n490), .A2(G129), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n470), .A2(G105), .ZN(new_n759));
  NAND3_X1  g334(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT26), .Z(new_n761));
  NAND4_X1  g336(.A1(new_n757), .A2(new_n758), .A3(new_n759), .A4(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G29), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n756), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT27), .B(G1996), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT30), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n767), .A2(G28), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(G28), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n768), .A2(new_n769), .A3(new_n763), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n658), .B2(new_n763), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n766), .A2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT101), .ZN(new_n773));
  INV_X1    g348(.A(G27), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n774), .B2(G29), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n774), .A2(G29), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n513), .B2(G29), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n775), .B1(new_n777), .B2(new_n773), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G2078), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n470), .A2(G103), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT25), .ZN(new_n781));
  OAI21_X1  g356(.A(G127), .B1(new_n478), .B2(new_n479), .ZN(new_n782));
  INV_X1    g357(.A(G115), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n463), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n781), .B1(new_n784), .B2(G2105), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n468), .A2(G139), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT98), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n763), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n763), .A2(G33), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n791), .A2(G2072), .ZN(new_n792));
  INV_X1    g367(.A(G2072), .ZN(new_n793));
  NOR3_X1   g368(.A1(new_n788), .A2(new_n793), .A3(new_n790), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n772), .B(new_n779), .C1(new_n792), .C2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(G16), .A2(G21), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G168), .B2(G16), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n797), .A2(G1966), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(G1966), .ZN(new_n799));
  INV_X1    g374(.A(G2078), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n800), .B(new_n775), .C1(new_n777), .C2(new_n773), .ZN(new_n801));
  NAND2_X1  g376(.A1(G160), .A2(G29), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT99), .B(KEYINPUT24), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G34), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(new_n763), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n802), .A2(G2084), .A3(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n798), .A2(new_n799), .A3(new_n801), .A4(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(G2084), .B1(new_n802), .B2(new_n805), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT31), .B(G11), .Z(new_n809));
  NOR4_X1   g384(.A1(new_n795), .A2(new_n807), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n755), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(KEYINPUT102), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT102), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n755), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n744), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n742), .A2(G2067), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n731), .A2(G1341), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n763), .A2(G35), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G162), .B2(new_n763), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT29), .Z(new_n820));
  INV_X1    g395(.A(G2090), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n815), .A2(new_n816), .A3(new_n817), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(KEYINPUT104), .ZN(new_n825));
  AOI211_X1 g400(.A(new_n744), .B(new_n822), .C1(new_n812), .C2(new_n814), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT104), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n826), .A2(new_n827), .A3(new_n816), .A4(new_n817), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n724), .A2(G22), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(G303), .B2(new_n723), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT97), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(G1971), .ZN(new_n835));
  MUX2_X1   g410(.A(G6), .B(G305), .S(G16), .Z(new_n836));
  XOR2_X1   g411(.A(KEYINPUT32), .B(G1981), .Z(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(G1976), .ZN(new_n839));
  INV_X1    g414(.A(G288), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(G16), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n842));
  OR2_X1    g417(.A1(G16), .A2(G23), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n842), .B1(new_n841), .B2(new_n843), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n839), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n845), .A2(new_n839), .A3(new_n846), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n835), .B(new_n838), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  XOR2_X1   g425(.A(KEYINPUT96), .B(KEYINPUT34), .Z(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n849), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(new_n847), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n855), .A2(new_n851), .A3(new_n835), .A4(new_n838), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n763), .A2(G25), .ZN(new_n858));
  OAI21_X1  g433(.A(G2104), .B1(new_n489), .B2(G107), .ZN(new_n859));
  INV_X1    g434(.A(G95), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n859), .B1(new_n860), .B2(new_n489), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT93), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n862), .B1(G131), .B2(new_n468), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n490), .A2(G119), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n858), .B1(new_n866), .B2(new_n763), .ZN(new_n867));
  XNOR2_X1  g442(.A(KEYINPUT35), .B(G1991), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT94), .Z(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n867), .B(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(G290), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(new_n723), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(G24), .B2(new_n723), .ZN(new_n874));
  INV_X1    g449(.A(G1986), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n871), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n876), .B1(new_n875), .B2(new_n874), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n857), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(KEYINPUT36), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT36), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n857), .A2(new_n880), .A3(new_n877), .ZN(new_n881));
  AOI22_X1  g456(.A1(new_n825), .A2(new_n828), .B1(new_n879), .B2(new_n881), .ZN(G311));
  NAND2_X1  g457(.A1(new_n825), .A2(new_n828), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n879), .A2(new_n881), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(G150));
  NAND3_X1  g460(.A1(new_n535), .A2(G93), .A3(new_n536), .ZN(new_n886));
  INV_X1    g461(.A(G67), .ZN(new_n887));
  AOI211_X1 g462(.A(new_n887), .B(new_n522), .C1(new_n524), .C2(new_n526), .ZN(new_n888));
  AND2_X1   g463(.A1(G80), .A2(G543), .ZN(new_n889));
  OAI21_X1  g464(.A(G651), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n558), .A2(G55), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n886), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(G860), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n893), .B(KEYINPUT37), .Z(new_n894));
  NOR2_X1   g469(.A1(new_n637), .A2(new_n644), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n572), .B(new_n892), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n895), .B(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n898), .B(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(KEYINPUT39), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT106), .ZN(new_n902));
  INV_X1    g477(.A(G860), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(new_n900), .B2(KEYINPUT39), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n894), .B1(new_n902), .B2(new_n904), .ZN(G145));
  XNOR2_X1  g480(.A(new_n762), .B(new_n740), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n502), .A2(new_n504), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n499), .A2(new_n507), .A3(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n906), .B(new_n908), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n785), .A2(new_n787), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n909), .B(new_n910), .ZN(new_n911));
  AOI22_X1  g486(.A1(G130), .A2(new_n490), .B1(new_n468), .B2(G142), .ZN(new_n912));
  OAI21_X1  g487(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n489), .A2(G118), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(KEYINPUT107), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n912), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n651), .B(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(new_n865), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT108), .ZN(new_n919));
  XOR2_X1   g494(.A(new_n911), .B(new_n919), .Z(new_n920));
  XNOR2_X1  g495(.A(new_n495), .B(new_n658), .ZN(new_n921));
  XOR2_X1   g496(.A(new_n921), .B(G160), .Z(new_n922));
  OR2_X1    g497(.A1(new_n922), .A2(KEYINPUT109), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(KEYINPUT109), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n920), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  XOR2_X1   g500(.A(new_n911), .B(new_n918), .Z(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(new_n922), .ZN(new_n927));
  INV_X1    g502(.A(G37), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n925), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT110), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT110), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n925), .A2(new_n927), .A3(new_n931), .A4(new_n928), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n930), .A2(KEYINPUT40), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT40), .B1(new_n930), .B2(new_n932), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(G395));
  INV_X1    g510(.A(G868), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n892), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n840), .A2(G290), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n872), .A2(G288), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(G305), .B(G303), .ZN(new_n941));
  OR3_X1    g516(.A1(new_n940), .A2(new_n941), .A3(KEYINPUT112), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(KEYINPUT112), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT112), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n938), .A2(new_n939), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n943), .A2(new_n945), .A3(new_n941), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n942), .A2(new_n946), .ZN(new_n947));
  XOR2_X1   g522(.A(new_n947), .B(KEYINPUT42), .Z(new_n948));
  NAND2_X1  g523(.A1(new_n637), .A2(G299), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n595), .A2(new_n634), .A3(new_n630), .A4(new_n636), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT111), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT41), .ZN(new_n953));
  AOI211_X1 g528(.A(new_n952), .B(new_n953), .C1(new_n949), .C2(new_n950), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n949), .A2(new_n953), .A3(new_n950), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n953), .B1(new_n949), .B2(new_n950), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n954), .B1(new_n957), .B2(new_n952), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n646), .B(new_n897), .ZN(new_n959));
  MUX2_X1   g534(.A(new_n951), .B(new_n958), .S(new_n959), .Z(new_n960));
  XNOR2_X1  g535(.A(new_n948), .B(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n937), .B1(new_n961), .B2(new_n936), .ZN(G295));
  OAI21_X1  g537(.A(new_n937), .B1(new_n961), .B2(new_n936), .ZN(G331));
  INV_X1    g538(.A(KEYINPUT114), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n548), .B1(new_n558), .B2(G51), .ZN(new_n965));
  AND4_X1   g540(.A1(new_n603), .A2(new_n604), .A3(new_n965), .A4(new_n546), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n603), .B1(new_n602), .B2(new_n604), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n968), .A2(G301), .ZN(new_n969));
  INV_X1    g544(.A(G168), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n554), .A2(new_n560), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT79), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n554), .A2(new_n555), .A3(new_n560), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n970), .B1(new_n974), .B2(new_n553), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n897), .B1(new_n969), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(G286), .A2(new_n974), .A3(new_n553), .ZN(new_n977));
  NAND2_X1  g552(.A1(G301), .A2(G168), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(new_n978), .A3(new_n896), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n949), .A2(new_n950), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n964), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n951), .A2(KEYINPUT114), .A3(new_n976), .A4(new_n979), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n976), .A2(KEYINPUT113), .A3(new_n979), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n896), .B1(new_n977), .B2(new_n978), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n984), .B1(new_n958), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n947), .ZN(new_n992));
  AOI21_X1  g567(.A(G37), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n977), .A2(new_n978), .A3(new_n896), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n994), .A2(new_n986), .A3(new_n987), .ZN(new_n995));
  INV_X1    g570(.A(new_n988), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n951), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT116), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n980), .B1(new_n955), .B2(new_n956), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT115), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n980), .B(KEYINPUT115), .C1(new_n955), .C2(new_n956), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n989), .A2(new_n1003), .A3(new_n951), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n998), .A2(new_n1001), .A3(new_n1002), .A4(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n947), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n993), .A2(new_n1006), .A3(KEYINPUT43), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n982), .A2(new_n983), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n981), .A2(KEYINPUT41), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n949), .A2(new_n953), .A3(new_n950), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(new_n952), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n956), .A2(KEYINPUT111), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1011), .A2(new_n1012), .A3(new_n988), .A4(new_n985), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n992), .B1(new_n1008), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT43), .B1(new_n993), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(KEYINPUT44), .B1(new_n1007), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT43), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n993), .A2(new_n1006), .A3(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1008), .A2(new_n992), .A3(new_n1013), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n928), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT43), .B1(new_n1021), .B2(new_n1014), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT44), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1017), .A2(new_n1025), .ZN(G397));
  INV_X1    g601(.A(G1996), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n762), .B(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G2067), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n740), .B(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1031), .B1(new_n869), .B2(new_n865), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n866), .A2(new_n870), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1034), .B1(new_n875), .B2(new_n872), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(new_n875), .B2(new_n872), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n485), .A2(G2105), .ZN(new_n1037));
  INV_X1    g612(.A(new_n476), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(G40), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1384), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n908), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT45), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1039), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1036), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G1966), .ZN(new_n1046));
  INV_X1    g621(.A(G40), .ZN(new_n1047));
  AOI211_X1 g622(.A(new_n1047), .B(new_n476), .C1(new_n485), .C2(G2105), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT123), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n513), .A2(new_n1049), .A3(KEYINPUT45), .A4(new_n1040), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1048), .A2(new_n1043), .A3(new_n1050), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n513), .A2(new_n1040), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1049), .B1(new_n1052), .B2(KEYINPUT45), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1046), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n513), .A2(new_n1040), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT50), .ZN(new_n1056));
  INV_X1    g631(.A(G2084), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n497), .A2(new_n498), .B1(new_n468), .B2(new_n506), .ZN(new_n1058));
  AOI21_X1  g633(.A(G1384), .B1(new_n1058), .B2(new_n907), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT118), .B(KEYINPUT50), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1056), .A2(new_n1048), .A3(new_n1057), .A4(new_n1062), .ZN(new_n1063));
  XOR2_X1   g638(.A(KEYINPUT119), .B(G8), .Z(new_n1064));
  NAND2_X1  g639(.A1(new_n970), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1054), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT123), .B1(new_n1055), .B2(new_n1042), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1067), .A2(new_n1048), .A3(new_n1043), .A4(new_n1050), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n1056), .A2(new_n1048), .A3(new_n1062), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1046), .A2(new_n1068), .B1(new_n1069), .B2(new_n1057), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n1065), .A2(G8), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1066), .B(KEYINPUT51), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1064), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1073), .B(new_n1065), .C1(new_n1070), .C2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT62), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT45), .B1(new_n513), .B2(new_n1040), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1039), .B1(KEYINPUT117), .B2(new_n1077), .ZN(new_n1078));
  AOI211_X1 g653(.A(new_n1042), .B(G1384), .C1(new_n1058), .C2(new_n907), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1055), .A2(new_n1042), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(G1971), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT50), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n513), .A2(new_n1084), .A3(new_n1040), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT122), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1041), .A2(new_n1060), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n513), .A2(new_n1088), .A3(new_n1084), .A4(new_n1040), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1086), .A2(new_n1048), .A3(new_n1087), .A4(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1090), .A2(G2090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1064), .B1(new_n1083), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(G303), .A2(G8), .ZN(new_n1093));
  XOR2_X1   g668(.A(new_n1093), .B(KEYINPUT55), .Z(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT49), .ZN(new_n1097));
  INV_X1    g672(.A(G86), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1098), .B1(new_n584), .B2(new_n585), .ZN(new_n1099));
  INV_X1    g674(.A(new_n618), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n1099), .A2(G1981), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(G1981), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n620), .A2(G86), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1102), .B1(new_n1103), .B2(new_n618), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1097), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n614), .A2(new_n1102), .A3(new_n618), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1103), .A2(new_n618), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(G1981), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1106), .A2(KEYINPUT49), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1074), .B1(new_n1048), .B2(new_n1059), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1105), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT120), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n609), .A2(G1976), .A3(new_n610), .A4(new_n611), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1110), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(G160), .A2(G40), .A3(new_n1059), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1115), .A2(G288), .A3(new_n839), .A4(new_n1064), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT52), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1114), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1119));
  AND4_X1   g694(.A1(new_n1112), .A2(new_n1113), .A3(new_n1115), .A4(new_n1064), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1111), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1056), .A2(new_n1048), .A3(new_n1062), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1123), .A2(G2090), .ZN(new_n1124));
  OAI211_X1 g699(.A(G8), .B(new_n1094), .C1(new_n1083), .C2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1096), .A2(new_n1122), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n800), .A2(KEYINPUT53), .ZN(new_n1127));
  OR2_X1    g702(.A1(new_n1068), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1123), .A2(new_n753), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1078), .A2(new_n1082), .A3(new_n800), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1128), .B(new_n1129), .C1(new_n1130), .C2(KEYINPUT53), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(G171), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1076), .A2(new_n1126), .A3(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1133), .A2(KEYINPUT127), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1136), .A2(KEYINPUT62), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT127), .ZN(new_n1138));
  NOR4_X1   g713(.A1(new_n1076), .A2(new_n1126), .A3(new_n1132), .A4(new_n1138), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1134), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(KEYINPUT125), .A2(KEYINPUT63), .ZN(new_n1141));
  OR2_X1    g716(.A1(KEYINPUT125), .A2(KEYINPUT63), .ZN(new_n1142));
  NOR4_X1   g717(.A1(new_n1070), .A2(KEYINPUT124), .A3(G286), .A4(new_n1074), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1074), .B1(new_n1054), .B2(new_n1063), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1144), .B1(new_n1145), .B2(new_n968), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1141), .B(new_n1142), .C1(new_n1147), .C2(new_n1126), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT63), .ZN(new_n1150));
  OAI21_X1  g725(.A(G8), .B1(new_n1083), .B2(new_n1124), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1150), .B1(new_n1151), .B2(new_n1095), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1149), .B(new_n1152), .C1(new_n1143), .C2(new_n1146), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1148), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1105), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1155), .A2(new_n839), .A3(new_n840), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n1106), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT121), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1125), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1158), .A2(new_n1110), .B1(new_n1159), .B2(new_n1122), .ZN(new_n1160));
  XNOR2_X1  g735(.A(KEYINPUT56), .B(G2072), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1078), .A2(new_n1082), .A3(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n595), .B(KEYINPUT57), .ZN(new_n1163));
  INV_X1    g738(.A(G1956), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1090), .A2(KEYINPUT126), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(KEYINPUT126), .B1(new_n1090), .B2(new_n1164), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1162), .B(new_n1163), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1123), .A2(new_n721), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1048), .A2(new_n1029), .A3(new_n1059), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n637), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1162), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1163), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1078), .A2(new_n1082), .A3(new_n1027), .ZN(new_n1176));
  XOR2_X1   g751(.A(KEYINPUT58), .B(G1341), .Z(new_n1177));
  NAND2_X1  g752(.A1(new_n1115), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n572), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1179), .B(KEYINPUT59), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1168), .A2(new_n637), .A3(new_n1169), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(KEYINPUT60), .B1(new_n1182), .B2(new_n1170), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n637), .A2(KEYINPUT60), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1184), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1180), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT61), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n1167), .B(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1175), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1126), .ZN(new_n1191));
  XOR2_X1   g766(.A(G301), .B(KEYINPUT54), .Z(new_n1192));
  INV_X1    g767(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1131), .A2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1079), .A2(new_n1127), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1195), .A2(new_n1048), .A3(new_n1043), .ZN(new_n1196));
  AND2_X1   g771(.A1(new_n1192), .A2(new_n1196), .ZN(new_n1197));
  OAI211_X1 g772(.A(new_n1197), .B(new_n1129), .C1(KEYINPUT53), .C2(new_n1130), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1191), .A2(new_n1136), .A3(new_n1194), .A4(new_n1198), .ZN(new_n1199));
  OAI211_X1 g774(.A(new_n1154), .B(new_n1160), .C1(new_n1190), .C2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1045), .B1(new_n1140), .B2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1044), .A2(new_n875), .A3(new_n872), .ZN(new_n1202));
  XOR2_X1   g777(.A(new_n1202), .B(KEYINPUT48), .Z(new_n1203));
  AOI21_X1  g778(.A(new_n1203), .B1(new_n1044), .B2(new_n1034), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT46), .ZN(new_n1205));
  INV_X1    g780(.A(new_n1044), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1205), .B1(new_n1206), .B2(G1996), .ZN(new_n1207));
  INV_X1    g782(.A(new_n1030), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1044), .B1(new_n762), .B2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1044), .A2(KEYINPUT46), .A3(new_n1027), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1207), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  XOR2_X1   g786(.A(new_n1211), .B(KEYINPUT47), .Z(new_n1212));
  OAI22_X1  g787(.A1(new_n1033), .A2(new_n1031), .B1(G2067), .B2(new_n740), .ZN(new_n1213));
  AOI211_X1 g788(.A(new_n1204), .B(new_n1212), .C1(new_n1044), .C2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1201), .A2(new_n1214), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g790(.A1(new_n678), .A2(G227), .ZN(new_n1217));
  AND2_X1   g791(.A1(new_n929), .A2(new_n1217), .ZN(new_n1218));
  AND4_X1   g792(.A1(G319), .A2(new_n1023), .A3(new_n716), .A4(new_n1218), .ZN(G308));
  NAND4_X1  g793(.A1(new_n1023), .A2(G319), .A3(new_n1218), .A4(new_n716), .ZN(G225));
endmodule


