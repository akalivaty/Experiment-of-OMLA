//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G107), .ZN(new_n188));
  OR2_X1    g002(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G104), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n188), .B1(new_n189), .B2(new_n191), .ZN(new_n192));
  NOR2_X1   g006(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n187), .A2(G107), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n193), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(G101), .B1(new_n192), .B2(new_n196), .ZN(new_n197));
  AND2_X1   g011(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n189), .B1(new_n191), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G101), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n194), .A2(new_n193), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n199), .A2(new_n200), .A3(new_n188), .A4(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n197), .A2(KEYINPUT4), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G143), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(G143), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT0), .A2(G128), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT0), .ZN(new_n213));
  INV_X1    g027(.A(G128), .ZN(new_n214));
  AOI22_X1  g028(.A1(new_n211), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n204), .A2(G143), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n217), .B1(new_n207), .B2(G146), .ZN(new_n218));
  INV_X1    g032(.A(new_n209), .ZN(new_n219));
  AOI22_X1  g033(.A1(new_n208), .A2(new_n215), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT4), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n221), .B(G101), .C1(new_n192), .C2(new_n196), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n203), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n191), .A2(new_n188), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G101), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n202), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n214), .B1(new_n216), .B2(KEYINPUT1), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n208), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G143), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT65), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT65), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G143), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n231), .A2(new_n233), .A3(G146), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n214), .A2(KEYINPUT1), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n216), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n229), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n226), .A2(new_n237), .A3(KEYINPUT10), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n223), .A2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n232), .A2(G143), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n230), .A2(KEYINPUT65), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n204), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n214), .B1(new_n242), .B2(KEYINPUT1), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n236), .B1(new_n243), .B2(new_n218), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(new_n226), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT10), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT78), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT78), .ZN(new_n248));
  AOI211_X1 g062(.A(new_n248), .B(KEYINPUT10), .C1(new_n244), .C2(new_n226), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n239), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT11), .ZN(new_n251));
  INV_X1    g065(.A(G134), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n251), .B1(new_n252), .B2(G137), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(G137), .ZN(new_n254));
  INV_X1    g068(.A(G137), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(KEYINPUT11), .A3(G134), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n253), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(KEYINPUT66), .A2(G131), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n253), .A2(new_n256), .A3(new_n258), .A4(new_n254), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n250), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n262), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n264), .B(new_n239), .C1(new_n247), .C2(new_n249), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(G110), .B(G140), .ZN(new_n267));
  INV_X1    g081(.A(G953), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n268), .A2(G227), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n267), .B(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT79), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n272), .B1(new_n226), .B2(new_n237), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n202), .A2(new_n225), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n274), .A2(KEYINPUT79), .A3(new_n229), .A4(new_n236), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n273), .A2(new_n245), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n262), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT12), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n276), .A2(KEYINPUT12), .A3(new_n262), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n223), .A2(new_n238), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n234), .A2(new_n216), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT1), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n231), .A2(new_n233), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n284), .B1(new_n285), .B2(new_n204), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n283), .B1(new_n286), .B2(new_n214), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n274), .B1(new_n236), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n248), .B1(new_n288), .B2(KEYINPUT10), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n245), .A2(KEYINPUT78), .A3(new_n246), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n282), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n270), .B1(new_n291), .B2(new_n264), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n281), .B1(new_n292), .B2(KEYINPUT80), .ZN(new_n293));
  INV_X1    g107(.A(new_n270), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n265), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT80), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n271), .B1(new_n293), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G469), .ZN(new_n299));
  INV_X1    g113(.A(G902), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n299), .A2(new_n300), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n281), .A2(new_n265), .ZN(new_n304));
  XOR2_X1   g118(.A(new_n270), .B(KEYINPUT76), .Z(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n292), .A2(new_n263), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(G469), .A3(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n301), .A2(new_n303), .A3(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT9), .B(G234), .ZN(new_n310));
  OAI21_X1  g124(.A(G221), .B1(new_n310), .B2(G902), .ZN(new_n311));
  OAI21_X1  g125(.A(G214), .B1(G237), .B2(G902), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n234), .A2(new_n219), .A3(new_n216), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n205), .B1(new_n285), .B2(new_n204), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n211), .A2(new_n212), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n213), .A2(new_n214), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n314), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G125), .ZN(new_n320));
  INV_X1    g134(.A(G125), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n229), .A2(new_n321), .A3(new_n236), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n268), .A2(G224), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n323), .B(new_n324), .ZN(new_n325));
  XOR2_X1   g139(.A(G116), .B(G119), .Z(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT2), .B(G113), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AND2_X1   g142(.A1(KEYINPUT2), .A2(G113), .ZN(new_n329));
  NOR2_X1   g143(.A1(KEYINPUT2), .A2(G113), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(G116), .B(G119), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n331), .A2(new_n332), .A3(KEYINPUT67), .ZN(new_n333));
  AOI21_X1  g147(.A(KEYINPUT67), .B1(new_n331), .B2(new_n332), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n328), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n203), .A2(new_n335), .A3(new_n222), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT67), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n337), .B1(new_n326), .B2(new_n327), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n331), .A2(new_n332), .A3(KEYINPUT67), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT5), .ZN(new_n341));
  INV_X1    g155(.A(G119), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n342), .A3(G116), .ZN(new_n343));
  OAI211_X1 g157(.A(G113), .B(new_n343), .C1(new_n326), .C2(new_n341), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n340), .A2(new_n202), .A3(new_n225), .A4(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n336), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(G110), .B(G122), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n336), .A2(new_n347), .A3(new_n345), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(KEYINPUT6), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT6), .ZN(new_n352));
  AND4_X1   g166(.A1(KEYINPUT81), .A2(new_n346), .A3(new_n352), .A4(new_n348), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n347), .B1(new_n336), .B2(new_n345), .ZN(new_n354));
  AOI21_X1  g168(.A(KEYINPUT81), .B1(new_n354), .B2(new_n352), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n325), .B(new_n351), .C1(new_n353), .C2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n320), .A2(KEYINPUT82), .A3(new_n322), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT82), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n229), .A2(new_n358), .A3(new_n321), .A4(new_n236), .ZN(new_n359));
  INV_X1    g173(.A(new_n324), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT7), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n357), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n347), .B(KEYINPUT8), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n344), .B1(new_n333), .B2(new_n334), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(new_n274), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n340), .A2(new_n344), .B1(new_n202), .B2(new_n225), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n363), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT83), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT7), .B1(new_n324), .B2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n369), .B1(new_n368), .B2(new_n324), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n320), .A2(new_n322), .A3(new_n370), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n362), .A2(new_n367), .A3(new_n350), .A4(new_n371), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n372), .A2(new_n300), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n356), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(G210), .B1(G237), .B2(G902), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n356), .A2(new_n373), .A3(new_n375), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n313), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G475), .ZN(new_n380));
  INV_X1    g194(.A(G237), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n381), .A2(new_n268), .A3(G143), .A4(G214), .ZN(new_n382));
  INV_X1    g196(.A(G214), .ZN(new_n383));
  NOR3_X1   g197(.A1(new_n383), .A2(G237), .A3(G953), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n382), .B1(new_n285), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G131), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT17), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n381), .A2(new_n268), .A3(G214), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(new_n231), .A3(new_n233), .ZN(new_n389));
  INV_X1    g203(.A(G131), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(new_n382), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n386), .A2(new_n387), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G140), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G125), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n321), .A2(G140), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n395), .A3(KEYINPUT16), .ZN(new_n396));
  OR3_X1    g210(.A1(new_n321), .A2(KEYINPUT16), .A3(G140), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n396), .A2(G146), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(G146), .B1(new_n396), .B2(new_n397), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n390), .B1(new_n389), .B2(new_n382), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT17), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n392), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n321), .A2(G140), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n393), .A2(G125), .ZN(new_n405));
  OAI21_X1  g219(.A(G146), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n394), .A2(new_n395), .A3(new_n204), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(KEYINPUT18), .A2(G131), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n389), .A2(new_n409), .A3(new_n382), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  AOI211_X1 g225(.A(KEYINPUT84), .B(new_n409), .C1(new_n389), .C2(new_n382), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT84), .ZN(new_n413));
  INV_X1    g227(.A(new_n409), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n413), .B1(new_n385), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n411), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n403), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G113), .B(G122), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(KEYINPUT86), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G104), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT86), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n418), .B(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n187), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n417), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n403), .A2(new_n416), .A3(new_n424), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n380), .B1(new_n428), .B2(new_n300), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT89), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n394), .A2(new_n395), .A3(KEYINPUT19), .ZN(new_n432));
  AOI21_X1  g246(.A(KEYINPUT19), .B1(new_n394), .B2(new_n395), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n204), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT85), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT19), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n436), .B1(new_n404), .B2(new_n405), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n394), .A2(new_n395), .A3(KEYINPUT19), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT85), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n440), .A3(new_n204), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n435), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n398), .B1(new_n386), .B2(new_n391), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n424), .B1(new_n444), .B2(new_n416), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT87), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n427), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n415), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n385), .A2(new_n413), .A3(new_n414), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n450), .A2(new_n411), .B1(new_n442), .B2(new_n443), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n451), .A2(KEYINPUT87), .A3(new_n424), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n431), .B1(new_n447), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT20), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT87), .B1(new_n451), .B2(new_n424), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n396), .A2(new_n397), .A3(G146), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n389), .A2(new_n390), .A3(new_n382), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n456), .B1(new_n457), .B2(new_n401), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n458), .B1(new_n441), .B2(new_n435), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n408), .A2(new_n410), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n460), .B1(new_n448), .B2(new_n449), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n446), .B(new_n425), .C1(new_n459), .C2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n455), .A2(new_n427), .A3(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(G475), .A2(G902), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(KEYINPUT88), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n453), .A2(new_n454), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  AND4_X1   g280(.A1(KEYINPUT89), .A2(new_n463), .A3(new_n454), .A4(new_n465), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n430), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G217), .ZN(new_n469));
  NOR3_X1   g283(.A1(new_n310), .A2(new_n469), .A3(G953), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(G116), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G122), .ZN(new_n473));
  INV_X1    g287(.A(G122), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(G116), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT90), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n473), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n476), .B1(new_n473), .B2(new_n475), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n190), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n231), .A2(new_n233), .A3(G128), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n214), .A2(G143), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n480), .A2(new_n252), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n252), .B1(new_n480), .B2(new_n481), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n479), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(KEYINPUT14), .B1(new_n474), .B2(G116), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT91), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n473), .A2(KEYINPUT91), .A3(KEYINPUT14), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n488), .A3(new_n475), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT92), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT92), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n487), .A2(new_n488), .A3(new_n491), .A4(new_n475), .ZN(new_n492));
  INV_X1    g306(.A(new_n473), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT14), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n490), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n484), .B1(new_n496), .B2(G107), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n477), .A2(new_n478), .A3(new_n190), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n473), .A2(new_n475), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT90), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n473), .A2(new_n475), .A3(new_n476), .ZN(new_n501));
  AOI21_X1  g315(.A(G107), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n480), .A2(new_n252), .A3(new_n481), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n480), .A2(KEYINPUT13), .A3(new_n481), .ZN(new_n505));
  OAI21_X1  g319(.A(G134), .B1(new_n480), .B2(KEYINPUT13), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n471), .B1(new_n497), .B2(new_n508), .ZN(new_n509));
  OAI221_X1 g323(.A(new_n504), .B1(new_n505), .B2(new_n506), .C1(new_n498), .C2(new_n502), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n489), .A2(KEYINPUT92), .B1(new_n494), .B2(new_n493), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n190), .B1(new_n511), .B2(new_n492), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n510), .B(new_n470), .C1(new_n512), .C2(new_n484), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n509), .A2(new_n513), .A3(KEYINPUT93), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n497), .A2(new_n508), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT93), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n516), .A3(new_n470), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n300), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT15), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT94), .B1(new_n519), .B2(G478), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(G478), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(KEYINPUT94), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n514), .A2(new_n517), .A3(new_n300), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n268), .A2(G952), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n526), .B1(G234), .B2(G237), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  AOI211_X1 g342(.A(new_n300), .B(new_n268), .C1(G234), .C2(G237), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  XOR2_X1   g344(.A(KEYINPUT21), .B(G898), .Z(new_n531));
  OAI21_X1  g345(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n525), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n468), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n309), .A2(new_n311), .A3(new_n379), .A4(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n208), .A2(new_n215), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n262), .A2(new_n536), .A3(new_n314), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n253), .A2(new_n256), .A3(new_n390), .A4(new_n254), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n252), .A2(G137), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n255), .A2(G134), .ZN(new_n540));
  OAI21_X1  g354(.A(G131), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n227), .B1(new_n242), .B2(new_n206), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n234), .A2(new_n216), .A3(new_n235), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n537), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n335), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n537), .A2(new_n545), .A3(new_n328), .A4(new_n340), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n547), .B1(new_n548), .B2(KEYINPUT70), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n548), .A2(KEYINPUT70), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT28), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n335), .B1(new_n546), .B2(KEYINPUT68), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT68), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n537), .A2(new_n545), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT28), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n381), .A2(new_n268), .A3(G210), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT27), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT26), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(new_n200), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(KEYINPUT29), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n300), .B1(new_n557), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT30), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n546), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n537), .A2(new_n545), .A3(KEYINPUT30), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(new_n335), .A3(new_n567), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n568), .A2(new_n548), .ZN(new_n569));
  INV_X1    g383(.A(new_n562), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT28), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n572), .B1(new_n547), .B2(new_n548), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n562), .B1(new_n555), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT29), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(G472), .B1(new_n564), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n568), .A2(new_n562), .A3(new_n548), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT31), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n570), .B1(new_n555), .B2(new_n573), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT31), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n568), .A2(new_n562), .A3(new_n580), .A4(new_n548), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(G472), .A2(G902), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT69), .ZN(new_n585));
  AOI21_X1  g399(.A(KEYINPUT32), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT32), .ZN(new_n587));
  AOI211_X1 g401(.A(KEYINPUT69), .B(new_n587), .C1(new_n582), .C2(new_n583), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n576), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n342), .A2(G128), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n214), .A2(KEYINPUT23), .A3(G119), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n342), .A2(G128), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n590), .B(new_n591), .C1(new_n592), .C2(KEYINPUT23), .ZN(new_n593));
  XOR2_X1   g407(.A(KEYINPUT24), .B(G110), .Z(new_n594));
  XNOR2_X1  g408(.A(G119), .B(G128), .ZN(new_n595));
  OAI22_X1  g409(.A1(new_n593), .A2(G110), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n596), .A2(new_n456), .A3(new_n407), .ZN(new_n597));
  OR2_X1    g411(.A1(new_n398), .A2(new_n399), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n593), .A2(G110), .B1(new_n594), .B2(new_n595), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT72), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n599), .B(KEYINPUT72), .C1(new_n399), .C2(new_n398), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n597), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT73), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT73), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n605), .B(new_n597), .C1(new_n600), .C2(new_n602), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n268), .A2(G221), .A3(G234), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(KEYINPUT74), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(KEYINPUT22), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(new_n255), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n604), .A2(new_n606), .A3(new_n610), .ZN(new_n611));
  OR2_X1    g425(.A1(new_n610), .A2(new_n603), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(G217), .A2(G902), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n614), .B1(new_n469), .B2(G234), .ZN(new_n615));
  XOR2_X1   g429(.A(new_n615), .B(KEYINPUT71), .Z(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n300), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT75), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n613), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n611), .A2(new_n300), .A3(new_n612), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n617), .B1(new_n621), .B2(KEYINPUT25), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT25), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n611), .A2(new_n612), .A3(new_n623), .A4(new_n300), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n620), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n589), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n535), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(new_n200), .ZN(G3));
  AND2_X1   g442(.A1(new_n309), .A2(new_n311), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n379), .A2(new_n532), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n465), .B1(new_n447), .B2(new_n452), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n403), .A2(new_n424), .A3(new_n416), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n425), .B1(new_n459), .B2(new_n461), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n632), .B1(new_n633), .B2(KEYINPUT87), .ZN(new_n634));
  AOI21_X1  g448(.A(KEYINPUT89), .B1(new_n634), .B2(new_n462), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n631), .B1(new_n635), .B2(KEYINPUT20), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n463), .A2(KEYINPUT89), .A3(new_n454), .A4(new_n465), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n429), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT33), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n514), .A2(new_n639), .A3(new_n517), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n509), .A2(new_n513), .A3(KEYINPUT33), .ZN(new_n641));
  INV_X1    g455(.A(G478), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(G902), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n518), .A2(new_n642), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g460(.A(KEYINPUT95), .B1(new_n638), .B2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT95), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n644), .A2(new_n645), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n468), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n630), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(G472), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n582), .B2(new_n300), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n653), .B1(new_n583), .B2(new_n582), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n629), .A2(new_n651), .A3(new_n625), .A4(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT34), .B(G104), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G6));
  XOR2_X1   g471(.A(new_n532), .B(KEYINPUT96), .Z(new_n658));
  AND3_X1   g472(.A1(new_n356), .A2(new_n375), .A3(new_n373), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n375), .B1(new_n356), .B2(new_n373), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n312), .B(new_n658), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n521), .A2(new_n524), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n463), .A2(KEYINPUT20), .A3(new_n465), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n429), .B1(new_n631), .B2(new_n454), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(KEYINPUT97), .B1(new_n661), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n631), .A2(new_n454), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n667), .A2(new_n430), .A3(new_n663), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n668), .A2(new_n525), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT97), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n379), .A2(new_n669), .A3(new_n670), .A4(new_n658), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n309), .A2(new_n625), .A3(new_n654), .A4(new_n311), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT35), .B(G107), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G9));
  INV_X1    g490(.A(new_n619), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n604), .A2(new_n606), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n678), .B1(KEYINPUT36), .B2(new_n610), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n610), .A2(KEYINPUT36), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n680), .A2(new_n604), .A3(new_n606), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  AOI22_X1  g496(.A1(new_n622), .A2(new_n624), .B1(new_n677), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n654), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n535), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT37), .B(G110), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G12));
  AND2_X1   g502(.A1(new_n589), .A2(new_n684), .ZN(new_n689));
  INV_X1    g503(.A(G900), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n527), .B1(new_n529), .B2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n662), .A2(new_n663), .A3(new_n664), .A4(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n312), .B1(new_n659), .B2(new_n660), .ZN(new_n694));
  OAI21_X1  g508(.A(KEYINPUT98), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n667), .A2(new_n430), .A3(new_n663), .A4(new_n692), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(new_n525), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT98), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n379), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n689), .A2(new_n629), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT99), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n214), .ZN(G30));
  NAND2_X1  g517(.A1(new_n377), .A2(new_n378), .ZN(new_n704));
  XOR2_X1   g518(.A(new_n704), .B(KEYINPUT38), .Z(new_n705));
  OR2_X1    g519(.A1(new_n569), .A2(new_n570), .ZN(new_n706));
  OR3_X1    g520(.A1(new_n549), .A2(new_n550), .A3(new_n562), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n706), .A2(new_n300), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(G472), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n709), .B1(new_n586), .B2(new_n588), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n525), .A2(new_n313), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n683), .A2(new_n468), .A3(new_n712), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n705), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(new_n691), .B(KEYINPUT39), .Z(new_n715));
  AND2_X1   g529(.A1(new_n629), .A2(new_n715), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n716), .A2(KEYINPUT40), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(KEYINPUT40), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n714), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(new_n285), .ZN(G45));
  NAND3_X1  g534(.A1(new_n468), .A2(new_n649), .A3(new_n692), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(KEYINPUT100), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT100), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n468), .A2(new_n723), .A3(new_n649), .A4(new_n692), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n722), .A2(new_n379), .A3(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n589), .A2(new_n309), .A3(new_n311), .A4(new_n684), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n204), .ZN(G48));
  AOI21_X1  g542(.A(new_n294), .B1(new_n263), .B2(new_n265), .ZN(new_n729));
  AOI22_X1  g543(.A1(new_n295), .A2(new_n296), .B1(new_n280), .B2(new_n279), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n292), .A2(KEYINPUT80), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(G469), .B1(new_n732), .B2(G902), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n733), .A2(new_n311), .A3(new_n301), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n651), .A2(new_n625), .A3(new_n589), .A4(new_n734), .ZN(new_n735));
  XOR2_X1   g549(.A(KEYINPUT41), .B(G113), .Z(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(KEYINPUT101), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n735), .B(new_n737), .ZN(G15));
  INV_X1    g552(.A(KEYINPUT102), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n733), .A2(new_n301), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n740), .A2(new_n625), .A3(new_n589), .A4(new_n311), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n739), .B1(new_n741), .B2(new_n672), .ZN(new_n742));
  INV_X1    g556(.A(new_n626), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n666), .A2(new_n671), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n743), .A2(KEYINPUT102), .A3(new_n744), .A4(new_n734), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G116), .ZN(G18));
  NAND4_X1  g561(.A1(new_n733), .A2(new_n301), .A3(new_n311), .A4(new_n379), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n749), .A2(new_n589), .A3(new_n534), .A4(new_n684), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G119), .ZN(G21));
  INV_X1    g565(.A(new_n625), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n583), .B(KEYINPUT103), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n578), .A2(new_n581), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n557), .A2(new_n570), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n752), .A2(new_n653), .A3(new_n757), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n468), .A2(new_n712), .A3(new_n704), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n758), .A2(new_n734), .A3(new_n658), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G122), .ZN(G24));
  NAND2_X1  g575(.A1(new_n636), .A2(new_n637), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n646), .B1(new_n762), .B2(new_n430), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n723), .B1(new_n763), .B2(new_n692), .ZN(new_n764));
  INV_X1    g578(.A(new_n724), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n683), .A2(new_n757), .A3(new_n653), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n766), .A2(KEYINPUT104), .A3(new_n749), .A4(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT104), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n722), .A2(new_n767), .A3(new_n724), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n769), .B1(new_n770), .B2(new_n748), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G125), .ZN(G27));
  NAND3_X1  g587(.A1(new_n304), .A2(KEYINPUT105), .A3(new_n305), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT105), .ZN(new_n775));
  AOI22_X1  g589(.A1(new_n279), .A2(new_n280), .B1(new_n264), .B2(new_n291), .ZN(new_n776));
  INV_X1    g590(.A(new_n305), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n774), .A2(new_n778), .A3(G469), .A4(new_n307), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n301), .A2(new_n303), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n311), .A2(new_n312), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n704), .A2(new_n781), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n766), .A2(new_n743), .A3(KEYINPUT106), .A4(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT42), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT106), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n589), .A2(new_n780), .A3(new_n625), .A4(new_n782), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n722), .A2(new_n724), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n784), .A2(new_n785), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n584), .A2(new_n587), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n576), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n584), .A2(new_n587), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n625), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n766), .A2(KEYINPUT42), .A3(new_n783), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n790), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT107), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(new_n390), .ZN(G33));
  NAND3_X1  g613(.A1(new_n743), .A2(new_n783), .A3(new_n697), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G134), .ZN(G36));
  NAND2_X1  g615(.A1(new_n638), .A2(new_n649), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT43), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n802), .B(new_n803), .C1(KEYINPUT109), .C2(new_n468), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT109), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n638), .B(new_n649), .C1(new_n805), .C2(KEYINPUT43), .ZN(new_n806));
  AOI211_X1 g620(.A(new_n654), .B(new_n683), .C1(new_n804), .C2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(KEYINPUT44), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n704), .A2(new_n313), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n311), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n306), .A2(new_n307), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT45), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n299), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n774), .A2(new_n778), .A3(KEYINPUT45), .A4(new_n307), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n817), .A2(KEYINPUT46), .A3(new_n303), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(KEYINPUT108), .A3(new_n301), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n302), .B1(new_n815), .B2(new_n816), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n820), .A2(KEYINPUT46), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT108), .B1(new_n818), .B2(new_n301), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n812), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n807), .A2(KEYINPUT44), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n811), .A2(new_n825), .A3(new_n715), .A4(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G137), .ZN(G39));
  XNOR2_X1  g642(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n819), .A2(new_n821), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n311), .B(new_n829), .C1(new_n830), .C2(new_n823), .ZN(new_n831));
  NOR4_X1   g645(.A1(new_n788), .A2(new_n625), .A3(new_n589), .A4(new_n810), .ZN(new_n832));
  NOR2_X1   g646(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n831), .B(new_n832), .C1(new_n825), .C2(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(G140), .ZN(G42));
  AND3_X1   g649(.A1(new_n740), .A2(new_n527), .A3(new_n782), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n804), .A2(new_n806), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n795), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(KEYINPUT48), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n528), .B1(new_n804), .B2(new_n806), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n841), .A2(new_n749), .A3(new_n758), .ZN(new_n842));
  XOR2_X1   g656(.A(new_n526), .B(KEYINPUT116), .Z(new_n843));
  AND3_X1   g657(.A1(new_n836), .A2(new_n625), .A3(new_n711), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n647), .A2(new_n650), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n840), .A2(new_n842), .A3(new_n843), .A4(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT51), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n831), .B1(new_n825), .B2(new_n833), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n740), .A2(new_n812), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n841), .A2(new_n758), .A3(new_n809), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT115), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n841), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n705), .A2(new_n313), .A3(new_n734), .A4(new_n758), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT50), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n838), .A2(new_n767), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n844), .A2(new_n638), .A3(new_n646), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n848), .B1(new_n855), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n853), .B1(new_n849), .B2(new_n850), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n865), .A2(new_n862), .A3(KEYINPUT51), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n847), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI211_X1 g683(.A(KEYINPUT117), .B(new_n847), .C1(new_n864), .C2(new_n866), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n683), .A2(new_n311), .A3(new_n692), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n873), .A2(new_n710), .A3(new_n759), .A4(new_n780), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n693), .A2(new_n694), .A3(KEYINPUT98), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n698), .B1(new_n697), .B2(new_n379), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n874), .B1(new_n726), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n878), .A2(new_n727), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n879), .A2(new_n772), .A3(KEYINPUT52), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT52), .B1(new_n879), .B2(new_n772), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n880), .A2(new_n881), .A3(KEYINPUT113), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT52), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n768), .A2(new_n771), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n701), .B(new_n874), .C1(new_n726), .C2(new_n725), .ZN(new_n885));
  OAI211_X1 g699(.A(KEYINPUT113), .B(new_n883), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n735), .A2(new_n750), .A3(new_n760), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n535), .B1(new_n626), .B2(new_n685), .ZN(new_n888));
  INV_X1    g702(.A(new_n661), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n638), .A2(KEYINPUT112), .A3(new_n662), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT112), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n891), .B1(new_n468), .B2(new_n525), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n889), .B(new_n890), .C1(new_n892), .C2(new_n763), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(new_n673), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n888), .A2(new_n894), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n887), .A2(new_n746), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n766), .A2(new_n767), .A3(new_n783), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n810), .A2(new_n662), .A3(new_n696), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n689), .A2(new_n898), .A3(new_n629), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n897), .A2(new_n800), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n790), .B2(new_n796), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n886), .A2(new_n896), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n872), .B1(new_n882), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT114), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n896), .B(new_n901), .C1(new_n880), .C2(new_n881), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n904), .B1(new_n905), .B2(new_n872), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n896), .A2(new_n901), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n879), .A2(new_n772), .A3(KEYINPUT52), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n907), .A2(KEYINPUT114), .A3(KEYINPUT53), .A4(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n903), .A2(new_n906), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT54), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT113), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n908), .A2(new_n914), .A3(new_n909), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n907), .A2(new_n915), .A3(KEYINPUT53), .A4(new_n886), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT54), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n905), .A2(new_n872), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n913), .A2(new_n919), .ZN(new_n920));
  OAI22_X1  g734(.A1(new_n871), .A2(new_n920), .B1(G952), .B2(G953), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n802), .A2(new_n752), .A3(new_n781), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT49), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n922), .B1(new_n923), .B2(new_n740), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT111), .Z(new_n925));
  NAND2_X1  g739(.A1(new_n740), .A2(new_n923), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n925), .A2(new_n705), .A3(new_n711), .A4(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n921), .A2(new_n927), .ZN(G75));
  NOR2_X1   g742(.A1(new_n268), .A2(G952), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n300), .B1(new_n916), .B2(new_n918), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT56), .B1(new_n931), .B2(G210), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n351), .B1(new_n353), .B2(new_n355), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(new_n325), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT55), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n930), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n932), .A2(new_n935), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT118), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n932), .A2(KEYINPUT118), .A3(new_n935), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n936), .B1(new_n939), .B2(new_n940), .ZN(G51));
  NAND2_X1  g755(.A1(new_n916), .A2(new_n918), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(KEYINPUT54), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n919), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n302), .B(KEYINPUT57), .Z(new_n946));
  OAI21_X1  g760(.A(new_n298), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n931), .A2(new_n816), .A3(new_n815), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n929), .B1(new_n947), .B2(new_n948), .ZN(G54));
  NAND3_X1  g763(.A1(new_n931), .A2(KEYINPUT58), .A3(G475), .ZN(new_n950));
  INV_X1    g764(.A(new_n463), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n929), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n950), .A2(new_n951), .ZN(new_n954));
  OAI21_X1  g768(.A(KEYINPUT119), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT119), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n952), .B(new_n956), .C1(new_n951), .C2(new_n950), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n955), .A2(new_n957), .ZN(G60));
  NAND2_X1  g772(.A1(new_n640), .A2(new_n641), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT120), .Z(new_n960));
  NAND2_X1  g774(.A1(G478), .A2(G902), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT59), .Z(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n960), .B1(new_n920), .B2(new_n963), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n960), .A2(new_n963), .ZN(new_n965));
  INV_X1    g779(.A(new_n919), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n917), .B1(new_n916), .B2(new_n918), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n930), .ZN(new_n969));
  OAI21_X1  g783(.A(KEYINPUT121), .B1(new_n964), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n929), .B1(new_n944), .B2(new_n965), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT121), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n962), .B1(new_n913), .B2(new_n919), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n971), .B(new_n972), .C1(new_n960), .C2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n970), .A2(new_n974), .ZN(G63));
  XNOR2_X1  g789(.A(new_n614), .B(KEYINPUT122), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT60), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n942), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n929), .B1(new_n978), .B2(new_n613), .ZN(new_n979));
  INV_X1    g793(.A(new_n682), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n979), .B1(new_n980), .B2(new_n978), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT61), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(G66));
  NAND3_X1  g797(.A1(new_n531), .A2(G224), .A3(G953), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n896), .B(KEYINPUT123), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n984), .B1(new_n985), .B2(G953), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n933), .B1(G898), .B2(new_n268), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n986), .B(new_n987), .Z(G69));
  NAND2_X1  g802(.A1(new_n797), .A2(new_n800), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT126), .Z(new_n990));
  AOI21_X1  g804(.A(new_n726), .B1(new_n725), .B2(new_n877), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n884), .A2(new_n991), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n825), .A2(new_n715), .A3(new_n759), .A4(new_n795), .ZN(new_n993));
  AND4_X1   g807(.A1(new_n827), .A2(new_n834), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n990), .A2(new_n268), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n566), .A2(new_n567), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(new_n439), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n997), .B1(G900), .B2(G953), .ZN(new_n998));
  AOI21_X1  g812(.A(KEYINPUT124), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n268), .B1(G227), .B2(G900), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(KEYINPUT125), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n992), .A2(new_n719), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n890), .B1(new_n892), .B2(new_n763), .ZN(new_n1004));
  NOR4_X1   g818(.A1(new_n1004), .A2(new_n626), .A3(new_n313), .A4(new_n704), .ZN(new_n1005));
  AOI22_X1  g819(.A1(new_n1003), .A2(KEYINPUT62), .B1(new_n716), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1006), .B1(KEYINPUT62), .B2(new_n1003), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n834), .A2(new_n827), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n268), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AOI22_X1  g823(.A1(new_n1009), .A2(new_n997), .B1(new_n995), .B2(new_n998), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1002), .B(new_n1010), .ZN(G72));
  XNOR2_X1  g825(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1012));
  NAND2_X1  g826(.A1(G472), .A2(G902), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  OR2_X1    g828(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1014), .B1(new_n1015), .B2(new_n985), .ZN(new_n1016));
  INV_X1    g830(.A(new_n706), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n912), .A2(new_n571), .A3(new_n706), .A4(new_n1014), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n990), .A2(new_n994), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1014), .B1(new_n1020), .B2(new_n985), .ZN(new_n1021));
  INV_X1    g835(.A(new_n571), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n929), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AND3_X1   g837(.A1(new_n1018), .A2(new_n1019), .A3(new_n1023), .ZN(G57));
endmodule


