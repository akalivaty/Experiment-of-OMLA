//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 0 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0008(.A(G77), .ZN(new_n209));
  INV_X1    g0009(.A(G244), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G107), .A2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n212), .B(new_n213), .C1(new_n202), .C2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n211), .B(new_n215), .C1(G116), .C2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n201), .C2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G1), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n220), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT1), .Z(new_n226));
  INV_X1    g0026(.A(new_n206), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n227), .A2(KEYINPUT67), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(KEYINPUT67), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n228), .A2(G50), .A3(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT68), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(KEYINPUT65), .ZN(new_n233));
  INV_X1    g0033(.A(KEYINPUT65), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n234), .A2(G1), .A3(G13), .ZN(new_n235));
  AND2_X1   g0035(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n222), .A2(KEYINPUT66), .ZN(new_n237));
  INV_X1    g0037(.A(KEYINPUT66), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n238), .A2(G20), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g0040(.A1(new_n236), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n231), .A2(new_n241), .ZN(new_n242));
  NOR2_X1   g0042(.A1(new_n224), .A2(G13), .ZN(new_n243));
  OAI211_X1 g0043(.A(new_n243), .B(G250), .C1(G257), .C2(G264), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT0), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n226), .A2(new_n242), .A3(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(G361));
  XNOR2_X1  g0047(.A(G250), .B(G257), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G264), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n249), .B(G270), .Z(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT2), .B(G226), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(G232), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G238), .B(G244), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n250), .B(new_n254), .ZN(G358));
  XNOR2_X1  g0055(.A(G68), .B(G77), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n256), .B(new_n217), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n257), .B(G58), .ZN(new_n258));
  XOR2_X1   g0058(.A(G107), .B(G116), .Z(new_n259));
  XNOR2_X1  g0059(.A(G87), .B(G97), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n259), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n258), .B(new_n261), .ZN(G351));
  OAI21_X1  g0062(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n263));
  INV_X1    g0063(.A(G150), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT66), .B(G20), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  XOR2_X1   g0070(.A(KEYINPUT8), .B(G58), .Z(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  OAI221_X1 g0072(.A(new_n263), .B1(new_n264), .B2(new_n266), .C1(new_n270), .C2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n274));
  AND3_X1   g0074(.A1(new_n233), .A2(new_n235), .A3(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n221), .A2(G13), .A3(G20), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n273), .A2(new_n276), .B1(new_n217), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n275), .B1(G1), .B2(new_n222), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G50), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  OR2_X1    g0083(.A1(new_n283), .A2(KEYINPUT9), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(KEYINPUT9), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G41), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n268), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n236), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT3), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n268), .ZN(new_n291));
  NAND2_X1  g0091(.A1(KEYINPUT3), .A2(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G1698), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G222), .ZN(new_n295));
  INV_X1    g0095(.A(G223), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n293), .B(new_n295), .C1(new_n296), .C2(new_n294), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n289), .B(new_n297), .C1(G77), .C2(new_n293), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n221), .B1(G41), .B2(G45), .ZN(new_n299));
  INV_X1    g0099(.A(G274), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  OAI211_X1 g0102(.A(G1), .B(G13), .C1(new_n268), .C2(new_n287), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n299), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G226), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n298), .A2(new_n302), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G200), .ZN(new_n308));
  INV_X1    g0108(.A(new_n307), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G190), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n286), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT70), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT10), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n312), .A2(KEYINPUT10), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n284), .A2(new_n285), .B1(G190), .B2(new_n309), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n316), .A2(new_n312), .A3(KEYINPUT10), .A4(new_n308), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n307), .A2(G179), .ZN(new_n319));
  INV_X1    g0119(.A(new_n283), .ZN(new_n320));
  INV_X1    g0120(.A(G169), .ZN(new_n321));
  AOI211_X1 g0121(.A(new_n319), .B(new_n320), .C1(new_n321), .C2(new_n307), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n271), .A2(new_n278), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n324), .B1(new_n280), .B2(new_n271), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n301), .B1(new_n305), .B2(G232), .ZN(new_n327));
  NAND2_X1  g0127(.A1(G33), .A2(G87), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n328), .B(KEYINPUT75), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT72), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n290), .ZN(new_n331));
  NAND2_X1  g0131(.A1(KEYINPUT72), .A2(KEYINPUT3), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n331), .A2(G33), .A3(new_n332), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n333), .A2(new_n291), .B1(new_n218), .B2(G1698), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n296), .A2(new_n294), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n329), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n289), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n327), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G200), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  XOR2_X1   g0140(.A(KEYINPUT77), .B(G190), .Z(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n342), .B(new_n327), .C1(new_n336), .C2(new_n337), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT73), .ZN(new_n345));
  AND2_X1   g0145(.A1(KEYINPUT3), .A2(G33), .ZN(new_n346));
  NOR2_X1   g0146(.A1(KEYINPUT3), .A2(G33), .ZN(new_n347));
  NOR3_X1   g0147(.A1(new_n346), .A2(new_n347), .A3(G20), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n345), .B1(new_n348), .B2(KEYINPUT7), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT7), .ZN(new_n350));
  OAI211_X1 g0150(.A(KEYINPUT73), .B(new_n350), .C1(new_n293), .C2(G20), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT74), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n331), .A2(new_n332), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n350), .B1(new_n354), .B2(new_n268), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n346), .B1(new_n237), .B2(new_n239), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n353), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AND2_X1   g0157(.A1(KEYINPUT72), .A2(KEYINPUT3), .ZN(new_n358));
  NOR2_X1   g0158(.A1(KEYINPUT72), .A2(KEYINPUT3), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n268), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n356), .A2(new_n360), .A3(new_n353), .A4(KEYINPUT7), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n352), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(G68), .ZN(new_n364));
  NAND2_X1  g0164(.A1(G58), .A2(G68), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n206), .A2(new_n365), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n366), .A2(G20), .B1(G159), .B2(new_n265), .ZN(new_n367));
  AOI21_X1  g0167(.A(KEYINPUT16), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n333), .A2(new_n222), .A3(new_n291), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT7), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n333), .A2(new_n240), .A3(new_n350), .A4(new_n291), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(G68), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n372), .A2(KEYINPUT16), .A3(new_n367), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n276), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n326), .B(new_n344), .C1(new_n368), .C2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n375), .A2(KEYINPUT78), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT78), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT16), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n360), .A2(new_n240), .A3(KEYINPUT7), .A4(new_n292), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT74), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n361), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n202), .B1(new_n381), .B2(new_n352), .ZN(new_n382));
  INV_X1    g0182(.A(new_n367), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n378), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AND2_X1   g0184(.A1(new_n373), .A2(new_n276), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n325), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n377), .B1(new_n386), .B2(new_n344), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT17), .B1(new_n376), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n375), .A2(KEYINPUT17), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n338), .A2(G169), .ZN(new_n392));
  OAI211_X1 g0192(.A(G179), .B(new_n327), .C1(new_n336), .C2(new_n337), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n380), .A2(new_n361), .B1(new_n349), .B2(new_n351), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n367), .B1(new_n395), .B2(new_n202), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n374), .B1(new_n378), .B2(new_n396), .ZN(new_n397));
  OAI211_X1 g0197(.A(KEYINPUT18), .B(new_n394), .C1(new_n397), .C2(new_n325), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT76), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n326), .B1(new_n368), .B2(new_n374), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n394), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT18), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n401), .A2(KEYINPUT76), .A3(KEYINPUT18), .A4(new_n394), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n400), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n271), .A2(new_n265), .B1(new_n267), .B2(G77), .ZN(new_n407));
  XNOR2_X1  g0207(.A(KEYINPUT15), .B(G87), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n407), .B1(new_n270), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n276), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n278), .A2(new_n209), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n281), .A2(G77), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT69), .ZN(new_n414));
  OR2_X1    g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n294), .A2(G232), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n293), .B(new_n416), .C1(new_n214), .C2(new_n294), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n289), .B(new_n417), .C1(G107), .C2(new_n293), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n418), .B(new_n302), .C1(new_n210), .C2(new_n304), .ZN(new_n419));
  INV_X1    g0219(.A(G190), .ZN(new_n420));
  OR2_X1    g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(G200), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n413), .A2(new_n414), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n415), .A2(new_n421), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n323), .A2(new_n391), .A3(new_n406), .A4(new_n424), .ZN(new_n425));
  OR2_X1    g0225(.A1(new_n304), .A2(KEYINPUT71), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n304), .A2(KEYINPUT71), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n426), .A2(G238), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n219), .A2(G1698), .ZN(new_n429));
  OAI221_X1 g0229(.A(new_n429), .B1(G226), .B2(G1698), .C1(new_n346), .C2(new_n347), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G33), .A2(G97), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n301), .B1(new_n432), .B2(new_n289), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT13), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n428), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n434), .B1(new_n428), .B2(new_n433), .ZN(new_n436));
  OAI21_X1  g0236(.A(G200), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n428), .A2(new_n433), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT13), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n428), .A2(new_n433), .A3(new_n434), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n439), .A2(G190), .A3(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n221), .A2(new_n202), .A3(G13), .A4(G20), .ZN(new_n442));
  XNOR2_X1  g0242(.A(new_n442), .B(KEYINPUT12), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n280), .B2(new_n202), .ZN(new_n444));
  OAI22_X1  g0244(.A1(new_n266), .A2(new_n217), .B1(new_n222), .B2(G68), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n445), .B1(new_n269), .B2(G77), .ZN(new_n446));
  OR3_X1    g0246(.A1(new_n446), .A2(KEYINPUT11), .A3(new_n275), .ZN(new_n447));
  OAI21_X1  g0247(.A(KEYINPUT11), .B1(new_n446), .B2(new_n275), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n444), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n437), .A2(new_n441), .A3(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(G169), .B1(new_n435), .B2(new_n436), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT14), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n439), .A2(G179), .A3(new_n440), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT14), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n454), .B(G169), .C1(new_n435), .C2(new_n436), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n452), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n449), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n450), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n419), .A2(G179), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n459), .B1(new_n415), .B2(new_n423), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n419), .A2(new_n321), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n425), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n277), .B1(G1), .B2(new_n268), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n276), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G116), .ZN(new_n468));
  XNOR2_X1  g0268(.A(KEYINPUT82), .B(G116), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(new_n277), .ZN(new_n470));
  XNOR2_X1  g0270(.A(new_n470), .B(KEYINPUT85), .ZN(new_n471));
  INV_X1    g0271(.A(G116), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT82), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT82), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G116), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n275), .B1(G20), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G283), .ZN(new_n478));
  INV_X1    g0278(.A(G97), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n240), .B(new_n478), .C1(G33), .C2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(KEYINPUT20), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n476), .A2(G20), .ZN(new_n482));
  AND4_X1   g0282(.A1(KEYINPUT20), .A2(new_n276), .A3(new_n480), .A4(new_n482), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n468), .B(new_n471), .C1(new_n481), .C2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT86), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n232), .B1(G33), .B2(G41), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n221), .A2(G45), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT5), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n287), .ZN(new_n491));
  NAND2_X1  g0291(.A1(KEYINPUT5), .A2(G41), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n487), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n488), .B1(new_n491), .B2(new_n492), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n494), .A2(G270), .B1(G274), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n294), .A2(G264), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n497), .B1(new_n333), .B2(new_n291), .ZN(new_n498));
  INV_X1    g0298(.A(G257), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n294), .ZN(new_n500));
  INV_X1    g0300(.A(new_n293), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n498), .A2(new_n500), .B1(G303), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n496), .B1(new_n502), .B2(new_n337), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G200), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n485), .A2(new_n486), .A3(new_n504), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n503), .A2(G200), .ZN(new_n506));
  OAI21_X1  g0306(.A(KEYINPUT86), .B1(new_n506), .B2(new_n484), .ZN(new_n507));
  OR2_X1    g0307(.A1(new_n503), .A2(new_n342), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n484), .A2(G169), .A3(new_n503), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT21), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n496), .B(G179), .C1(new_n502), .C2(new_n337), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n484), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n484), .A2(new_n503), .A3(KEYINPUT21), .A4(G169), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n512), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n509), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n467), .A2(G97), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n278), .A2(new_n479), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT6), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n521), .A2(new_n479), .A3(G107), .ZN(new_n522));
  XNOR2_X1  g0322(.A(G97), .B(G107), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n522), .B1(new_n523), .B2(new_n521), .ZN(new_n524));
  OAI22_X1  g0324(.A1(new_n524), .A2(new_n240), .B1(new_n209), .B2(new_n266), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n525), .B1(new_n363), .B2(G107), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n519), .B(new_n520), .C1(new_n526), .C2(new_n275), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n493), .A2(new_n489), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n528), .A2(G257), .A3(new_n303), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT79), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n494), .A2(KEYINPUT79), .A3(G257), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n495), .A2(G274), .ZN(new_n534));
  OAI211_X1 g0334(.A(G250), .B(G1698), .C1(new_n346), .C2(new_n347), .ZN(new_n535));
  OAI211_X1 g0335(.A(KEYINPUT4), .B(new_n294), .C1(new_n346), .C2(new_n347), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n478), .B(new_n535), .C1(new_n536), .C2(new_n210), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n333), .A2(new_n291), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n538), .A2(G244), .A3(new_n294), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT4), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n533), .B(new_n534), .C1(new_n541), .C2(new_n337), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(G179), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n542), .A2(new_n321), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n527), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n525), .ZN(new_n548));
  INV_X1    g0348(.A(G107), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n548), .B1(new_n395), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n550), .A2(new_n276), .B1(new_n479), .B2(new_n278), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n539), .A2(new_n540), .ZN(new_n552));
  INV_X1    g0352(.A(new_n537), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n337), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n555), .A2(G190), .A3(new_n534), .A4(new_n533), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n542), .A2(G200), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n551), .A2(new_n556), .A3(new_n519), .A4(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT80), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n547), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n559), .B1(new_n547), .B2(new_n558), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n518), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT83), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n240), .A2(G33), .A3(G97), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT19), .ZN(new_n565));
  NAND3_X1  g0365(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n240), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(G87), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(new_n479), .A3(new_n549), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n564), .A2(new_n565), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n538), .A2(G68), .A3(new_n240), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n275), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n408), .A2(new_n278), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n563), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n566), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n569), .B1(new_n267), .B2(new_n576), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n267), .A2(new_n268), .A3(new_n479), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n577), .B1(new_n578), .B2(KEYINPUT19), .ZN(new_n579));
  AOI211_X1 g0379(.A(new_n202), .B(new_n267), .C1(new_n291), .C2(new_n333), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n276), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n581), .A2(KEYINPUT83), .A3(new_n573), .ZN(new_n582));
  XNOR2_X1  g0382(.A(new_n408), .B(KEYINPUT84), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n575), .A2(new_n582), .B1(new_n467), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(G250), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n300), .B1(new_n585), .B2(KEYINPUT81), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n489), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n488), .A2(KEYINPUT81), .A3(G250), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n487), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n473), .A2(new_n475), .A3(G33), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n333), .A2(new_n291), .B1(new_n210), .B2(G1698), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n214), .A2(new_n294), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n590), .B1(new_n595), .B2(new_n337), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n597), .A2(G169), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n596), .A2(G179), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n584), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n575), .A2(new_n582), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n596), .A2(G200), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n467), .A2(G87), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n597), .A2(G190), .ZN(new_n604));
  AND4_X1   g0404(.A1(new_n601), .A2(new_n602), .A3(new_n603), .A4(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  NOR3_X1   g0406(.A1(new_n501), .A2(new_n267), .A3(new_n568), .ZN(new_n607));
  OR2_X1    g0407(.A1(new_n607), .A2(KEYINPUT22), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n538), .A2(KEYINPUT22), .A3(G87), .A4(new_n240), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT23), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n610), .A2(new_n549), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n591), .A2(new_n610), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n611), .B1(new_n612), .B2(new_n222), .ZN(new_n613));
  NOR2_X1   g0413(.A1(KEYINPUT23), .A2(G107), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n237), .A2(new_n239), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(KEYINPUT87), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(G20), .B1(new_n591), .B2(new_n610), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT87), .ZN(new_n619));
  NOR4_X1   g0419(.A1(new_n618), .A2(new_n619), .A3(new_n615), .A4(new_n611), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n608), .B(new_n609), .C1(new_n617), .C2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT24), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n611), .ZN(new_n624));
  AOI21_X1  g0424(.A(KEYINPUT23), .B1(new_n469), .B2(G33), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n616), .B(new_n624), .C1(new_n625), .C2(G20), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n619), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n613), .A2(KEYINPUT87), .A3(new_n616), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n629), .A2(KEYINPUT24), .A3(new_n608), .A4(new_n609), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n623), .A2(new_n276), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n467), .A2(G107), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n277), .A2(G107), .ZN(new_n633));
  XNOR2_X1  g0433(.A(new_n633), .B(KEYINPUT25), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n631), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n494), .A2(G264), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n333), .A2(new_n291), .B1(new_n499), .B2(G1698), .ZN(new_n637));
  OR2_X1    g0437(.A1(G250), .A2(G1698), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n637), .A2(new_n638), .B1(G33), .B2(G294), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n534), .B(new_n636), .C1(new_n639), .C2(new_n337), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(G179), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n641), .B1(new_n321), .B2(new_n640), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n635), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n640), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n644), .A2(new_n339), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(G190), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n631), .A2(new_n632), .A3(new_n634), .A4(new_n646), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n606), .B(new_n643), .C1(new_n645), .C2(new_n647), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n465), .A2(new_n562), .A3(new_n648), .ZN(G372));
  INV_X1    g0449(.A(new_n322), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n404), .A2(new_n398), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n456), .A2(new_n457), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n450), .B2(new_n462), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n651), .B1(new_n391), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n650), .B1(new_n654), .B2(new_n318), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n527), .A2(new_n545), .A3(new_n546), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n467), .A2(new_n583), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n601), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT88), .ZN(new_n660));
  OR3_X1    g0460(.A1(new_n595), .A2(new_n660), .A3(new_n337), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n660), .B1(new_n595), .B2(new_n337), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(new_n590), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n321), .ZN(new_n664));
  INV_X1    g0464(.A(new_n599), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n659), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n663), .A2(G200), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n667), .A2(new_n601), .A3(new_n603), .A4(new_n604), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n657), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT26), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT89), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n600), .A2(new_n547), .A3(new_n605), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(KEYINPUT26), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT89), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n669), .A2(new_n675), .A3(new_n670), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n672), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n666), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n512), .A2(new_n515), .A3(new_n516), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n601), .A2(new_n603), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n680), .B1(G190), .B2(new_n597), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n643), .A2(new_n679), .B1(new_n681), .B2(new_n667), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n547), .A2(new_n558), .ZN(new_n683));
  INV_X1    g0483(.A(new_n647), .ZN(new_n684));
  INV_X1    g0484(.A(new_n645), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n678), .B1(new_n682), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n677), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n656), .B1(new_n465), .B2(new_n689), .ZN(G369));
  INV_X1    g0490(.A(G13), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n267), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n221), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT27), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n692), .A2(new_n695), .A3(new_n221), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n694), .A2(G213), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G343), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT90), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n484), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n518), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n679), .B2(new_n701), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G330), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n684), .A2(new_n685), .B1(new_n635), .B2(new_n642), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n635), .A2(new_n700), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n635), .A2(new_n642), .A3(new_n700), .ZN(new_n709));
  OR2_X1    g0509(.A1(new_n709), .A2(KEYINPUT91), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(KEYINPUT91), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n708), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n705), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n643), .A2(new_n700), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n679), .A2(new_n700), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n715), .B1(new_n712), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n714), .A2(new_n717), .ZN(G399));
  INV_X1    g0518(.A(new_n243), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G41), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n569), .A2(G116), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(G1), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n231), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(new_n721), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT92), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT28), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n700), .B1(new_n677), .B2(new_n687), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT29), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT95), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n657), .A2(new_n668), .A3(new_n666), .A4(KEYINPUT26), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n731), .B(new_n732), .C1(new_n673), .C2(KEYINPUT26), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n732), .A2(new_n731), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n700), .B1(new_n735), .B2(new_n687), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n730), .B1(new_n736), .B2(new_n729), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n679), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n561), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n547), .A2(new_n558), .A3(new_n559), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n698), .B(KEYINPUT90), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n742), .A2(new_n706), .A3(new_n606), .A4(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT31), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT30), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n636), .B1(new_n639), .B2(new_n337), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n747), .B1(new_n513), .B2(KEYINPUT93), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n543), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n597), .B1(KEYINPUT93), .B2(new_n513), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n746), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n750), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n752), .A2(KEYINPUT30), .A3(new_n543), .A4(new_n748), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n542), .A2(new_n640), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(KEYINPUT94), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n755), .A2(new_n503), .A3(new_n663), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n544), .B1(new_n754), .B2(KEYINPUT94), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n751), .B(new_n753), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n745), .B1(new_n758), .B2(new_n700), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n758), .A2(new_n745), .A3(new_n700), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n744), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n737), .B1(G330), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n727), .B1(new_n764), .B2(G1), .ZN(G364));
  NAND2_X1  g0565(.A1(new_n692), .A2(G45), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n721), .A2(G1), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n703), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n236), .B1(G20), .B2(new_n321), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G179), .A2(G200), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G190), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n267), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n479), .ZN(new_n778));
  OAI21_X1  g0578(.A(KEYINPUT97), .B1(new_n240), .B2(new_n544), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT97), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n267), .A2(new_n780), .A3(G179), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n339), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G190), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n782), .A2(new_n420), .A3(G200), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n785), .A2(new_n209), .B1(new_n202), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n267), .A2(new_n420), .A3(new_n774), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G159), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n778), .B(new_n787), .C1(KEYINPUT32), .C2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n339), .A2(G179), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n267), .A2(new_n420), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n549), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n782), .A2(G200), .A3(new_n341), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n794), .B1(new_n796), .B2(G50), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n783), .A2(new_n342), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n797), .B1(new_n201), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n792), .A2(G20), .A3(G190), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n800), .B1(G87), .B2(new_n802), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n790), .A2(KEYINPUT32), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n791), .A2(new_n293), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n798), .A2(G322), .ZN(new_n806));
  INV_X1    g0606(.A(G303), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n801), .B(KEYINPUT98), .ZN(new_n808));
  INV_X1    g0608(.A(G311), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n501), .B1(new_n807), .B2(new_n808), .C1(new_n785), .C2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(G294), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n777), .A2(new_n811), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n789), .A2(G329), .ZN(new_n813));
  NOR4_X1   g0613(.A1(new_n806), .A2(new_n810), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(G283), .ZN(new_n815));
  XOR2_X1   g0615(.A(KEYINPUT33), .B(G317), .Z(new_n816));
  OAI221_X1 g0616(.A(new_n814), .B1(new_n815), .B2(new_n793), .C1(new_n786), .C2(new_n816), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n796), .A2(G326), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n805), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n767), .B(new_n772), .C1(new_n773), .C2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n243), .A2(new_n293), .ZN(new_n821));
  INV_X1    g0621(.A(G355), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n821), .A2(new_n822), .B1(G116), .B2(new_n243), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT96), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n724), .A2(G45), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n719), .A2(new_n538), .ZN(new_n826));
  INV_X1    g0626(.A(G45), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n826), .B1(new_n258), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n824), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n773), .A2(new_n770), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n820), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n767), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n705), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(G330), .B2(new_n703), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G396));
  INV_X1    g0637(.A(new_n538), .ZN(new_n838));
  INV_X1    g0638(.A(new_n786), .ZN(new_n839));
  AOI22_X1  g0639(.A1(G143), .A2(new_n798), .B1(new_n839), .B2(G150), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n796), .A2(G137), .ZN(new_n841));
  INV_X1    g0641(.A(G159), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n840), .B(new_n841), .C1(new_n842), .C2(new_n785), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT34), .Z(new_n844));
  INV_X1    g0644(.A(new_n808), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n838), .B(new_n844), .C1(G50), .C2(new_n845), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n846), .B1(new_n201), .B2(new_n777), .C1(new_n202), .C2(new_n793), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(G132), .B2(new_n789), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n778), .B1(new_n839), .B2(G283), .ZN(new_n849));
  INV_X1    g0649(.A(new_n793), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(G87), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n849), .A2(new_n501), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(G107), .B2(new_n845), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n784), .A2(new_n469), .B1(G311), .B2(new_n789), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n853), .B(new_n854), .C1(new_n811), .C2(new_n799), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(G303), .B2(new_n796), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n773), .B1(new_n848), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n773), .A2(new_n768), .ZN(new_n858));
  XOR2_X1   g0658(.A(new_n858), .B(KEYINPUT99), .Z(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n209), .ZN(new_n860));
  INV_X1    g0660(.A(new_n423), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n413), .A2(new_n414), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n424), .B1(new_n863), .B2(new_n743), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n462), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n462), .B2(new_n700), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n768), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n857), .A2(new_n833), .A3(new_n860), .A4(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n460), .A2(new_n461), .A3(new_n743), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n728), .B(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n763), .A2(G330), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n871), .B(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n868), .B1(new_n873), .B2(new_n833), .ZN(G384));
  XNOR2_X1  g0674(.A(new_n869), .B(KEYINPUT101), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n728), .B2(new_n870), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT102), .ZN(new_n877));
  INV_X1    g0677(.A(new_n450), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n700), .A2(new_n457), .ZN(new_n879));
  AND4_X1   g0679(.A1(new_n877), .A2(new_n652), .A3(new_n878), .A4(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n879), .B1(new_n458), .B2(new_n877), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n876), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  INV_X1    g0684(.A(new_n697), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT16), .B1(new_n372), .B2(new_n367), .ZN(new_n886));
  OR2_X1    g0686(.A1(new_n374), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n885), .B1(new_n887), .B2(new_n326), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n391), .B2(new_n406), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n375), .A2(KEYINPUT78), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n386), .A2(new_n377), .A3(new_n344), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n394), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n887), .B2(new_n326), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n893), .A2(new_n889), .A3(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT103), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n386), .B2(new_n885), .ZN(new_n899));
  OAI211_X1 g0699(.A(KEYINPUT103), .B(new_n697), .C1(new_n397), .C2(new_n325), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT37), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n891), .A2(new_n892), .B1(new_n401), .B2(new_n394), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n897), .A2(KEYINPUT37), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n884), .B1(new_n890), .B2(new_n903), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n400), .A2(new_n404), .A3(new_n405), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n389), .B1(new_n893), .B2(KEYINPUT17), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n888), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n902), .A2(new_n901), .ZN(new_n908));
  AOI211_X1 g0708(.A(new_n888), .B(new_n895), .C1(new_n891), .C2(new_n892), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT37), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n907), .A2(new_n911), .A3(KEYINPUT38), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n904), .A2(new_n912), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n883), .A2(new_n913), .B1(new_n651), .B2(new_n885), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n890), .A2(new_n903), .A3(new_n884), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT38), .B1(new_n907), .B2(new_n911), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT39), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT104), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n913), .A2(KEYINPUT104), .A3(KEYINPUT39), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n899), .A2(new_n900), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n404), .A2(new_n398), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n921), .B1(new_n391), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n921), .A2(new_n375), .A3(new_n402), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n924), .A2(KEYINPUT37), .B1(new_n901), .B2(new_n902), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n884), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT39), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n926), .A2(new_n927), .A3(new_n912), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(KEYINPUT105), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT105), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n926), .A2(new_n912), .A3(new_n930), .A4(new_n927), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n919), .A2(new_n920), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n652), .A2(new_n700), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n914), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n655), .B1(new_n737), .B2(new_n464), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n935), .B(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n870), .B1(new_n880), .B2(new_n881), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n744), .B2(new_n762), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n913), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT40), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n899), .B(new_n900), .C1(new_n906), .C2(new_n651), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n375), .B1(new_n386), .B2(new_n894), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n899), .B2(new_n900), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n908), .B1(new_n910), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(KEYINPUT38), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n939), .B(KEYINPUT40), .C1(new_n915), .C2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n942), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n464), .A2(new_n763), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n949), .B(new_n950), .Z(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(G330), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n937), .B(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n221), .B2(new_n692), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n231), .A2(G77), .A3(new_n365), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(G50), .B2(new_n202), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n956), .A2(G1), .A3(new_n691), .ZN(new_n957));
  INV_X1    g0757(.A(new_n524), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n472), .B1(new_n958), .B2(KEYINPUT35), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n959), .B(new_n241), .C1(KEYINPUT35), .C2(new_n958), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT100), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT36), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n954), .A2(new_n957), .A3(new_n962), .ZN(G367));
  NAND2_X1  g0763(.A1(new_n700), .A2(new_n527), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n964), .A2(new_n547), .A3(new_n558), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n657), .A2(new_n700), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n712), .A2(new_n716), .A3(new_n967), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n968), .A2(KEYINPUT42), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n547), .B1(new_n965), .B2(new_n643), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n743), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n968), .A2(KEYINPUT42), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n969), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n700), .A2(new_n680), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT106), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n678), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n668), .A2(new_n666), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n976), .B1(new_n977), .B2(new_n975), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n973), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n967), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n714), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n980), .B(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n983), .B(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n720), .B(KEYINPUT41), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(KEYINPUT44), .B1(new_n717), .B2(new_n967), .ZN(new_n988));
  OR3_X1    g0788(.A1(new_n717), .A2(KEYINPUT44), .A3(new_n967), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n717), .A2(new_n967), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT45), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(KEYINPUT45), .B1(new_n717), .B2(new_n967), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n988), .B(new_n989), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n994), .A2(new_n713), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n713), .ZN(new_n996));
  INV_X1    g0796(.A(new_n737), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n872), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n712), .B(new_n716), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(new_n704), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n995), .A2(new_n996), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n987), .B1(new_n1002), .B2(new_n764), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n766), .A2(G1), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n985), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n785), .A2(new_n815), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT46), .ZN(new_n1007));
  NOR3_X1   g0807(.A1(new_n808), .A2(new_n1007), .A3(new_n472), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n538), .B(new_n1008), .C1(G107), .C2(new_n776), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1007), .B1(new_n801), .B2(new_n476), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n850), .A2(G97), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n839), .A2(G294), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1006), .B(new_n1013), .C1(G317), .C2(new_n789), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n807), .B2(new_n799), .C1(new_n809), .C2(new_n795), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n793), .A2(new_n209), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n777), .A2(new_n202), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n796), .B2(G143), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n264), .B2(new_n799), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT108), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n789), .A2(G137), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n293), .B1(new_n786), .B2(new_n842), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G58), .B2(new_n802), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n784), .A2(G50), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1020), .A2(new_n1021), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1015), .B1(new_n1016), .B2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT47), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n773), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n978), .A2(new_n771), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n826), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n830), .B1(new_n243), .B2(new_n408), .C1(new_n250), .C2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT107), .Z(new_n1032));
  NAND4_X1  g0832(.A1(new_n1028), .A2(new_n833), .A3(new_n1029), .A4(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1005), .A2(new_n1033), .ZN(G387));
  OAI21_X1  g0834(.A(new_n538), .B1(new_n786), .B2(new_n272), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n795), .A2(new_n842), .B1(new_n209), .B2(new_n801), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1035), .B(new_n1036), .C1(G150), .C2(new_n789), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n784), .A2(G68), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n583), .A2(new_n776), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n798), .A2(G50), .B1(G97), .B2(new_n850), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  XOR2_X1   g0841(.A(KEYINPUT110), .B(G322), .Z(new_n1042));
  AOI22_X1  g0842(.A1(G317), .A2(new_n798), .B1(new_n796), .B2(new_n1042), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n807), .B2(new_n785), .C1(new_n809), .C2(new_n786), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT48), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n815), .B2(new_n777), .C1(new_n811), .C2(new_n801), .ZN(new_n1046));
  XOR2_X1   g0846(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n1047));
  AOI22_X1  g0847(.A1(new_n1046), .A2(new_n1047), .B1(G326), .B2(new_n789), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1048), .B(new_n838), .C1(new_n476), .C2(new_n793), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1041), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n1051), .A2(new_n773), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n712), .A2(new_n771), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n722), .B(new_n827), .C1(new_n202), .C2(new_n209), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT109), .Z(new_n1055));
  NAND2_X1  g0855(.A1(new_n271), .A2(new_n217), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT50), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n826), .B1(new_n254), .B2(new_n827), .C1(new_n1055), .C2(new_n1057), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(G107), .B2(new_n243), .C1(new_n722), .C2(new_n821), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n1059), .A2(new_n830), .ZN(new_n1060));
  NOR4_X1   g0860(.A1(new_n1052), .A2(new_n767), .A3(new_n1053), .A4(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n999), .B(new_n705), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1061), .B1(new_n1062), .B2(new_n1004), .ZN(new_n1063));
  OAI21_X1  g0863(.A(KEYINPUT112), .B1(new_n1001), .B2(new_n721), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n998), .A2(new_n1000), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n764), .A2(new_n1062), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT112), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1066), .A2(new_n1067), .A3(new_n720), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1064), .A2(new_n1065), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1063), .A2(new_n1069), .ZN(G393));
  AOI22_X1  g0870(.A1(G311), .A2(new_n798), .B1(new_n796), .B2(G317), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT52), .Z(new_n1072));
  NAND2_X1  g0872(.A1(new_n789), .A2(new_n1042), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1072), .B(new_n1073), .C1(new_n811), .C2(new_n785), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n786), .A2(new_n807), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n501), .B1(new_n815), .B2(new_n801), .C1(new_n777), .C2(new_n476), .ZN(new_n1076));
  NOR4_X1   g0876(.A1(new_n1074), .A2(new_n794), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n799), .A2(new_n842), .B1(new_n264), .B2(new_n795), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT51), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n538), .B1(new_n202), .B2(new_n801), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(G77), .B2(new_n776), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n784), .A2(new_n271), .B1(G143), .B2(new_n789), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1079), .A2(new_n851), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G50), .B2(new_n839), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n773), .B1(new_n1077), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n981), .A2(new_n770), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n830), .B1(new_n479), .B2(new_n243), .C1(new_n1030), .C2(new_n261), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1085), .A2(new_n833), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n995), .A2(new_n996), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1004), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n721), .B1(new_n1089), .B2(new_n1066), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1091), .B1(new_n1002), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(G390));
  NAND3_X1  g0894(.A1(new_n464), .A2(G330), .A3(new_n763), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n882), .B1(new_n872), .B2(new_n866), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n462), .A2(new_n700), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n736), .B2(new_n865), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n882), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n763), .A2(new_n1099), .A3(G330), .A4(new_n870), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n1096), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n876), .B1(new_n1096), .B2(new_n1100), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n936), .B(new_n1095), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n929), .A2(new_n931), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n934), .B1(new_n876), .B2(new_n882), .ZN(new_n1105));
  AOI21_X1  g0905(.A(KEYINPUT104), .B1(new_n913), .B2(KEYINPUT39), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n918), .B(new_n927), .C1(new_n904), .C2(new_n912), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1104), .B(new_n1105), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n934), .B1(new_n915), .B2(new_n947), .C1(new_n1098), .C2(new_n882), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n1108), .A2(new_n1109), .A3(new_n1100), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1100), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1103), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1100), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1103), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1108), .A2(new_n1109), .A3(new_n1100), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1112), .A2(new_n1118), .A3(new_n720), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1115), .A2(new_n1004), .A3(new_n1117), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n932), .A2(new_n768), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n859), .A2(new_n272), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n793), .A2(new_n217), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(G132), .A2(new_n798), .B1(new_n796), .B2(G128), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT113), .ZN(new_n1125));
  XOR2_X1   g0925(.A(KEYINPUT54), .B(G143), .Z(new_n1126));
  AOI21_X1  g0926(.A(new_n501), .B1(new_n784), .B2(new_n1126), .ZN(new_n1127));
  OR3_X1    g0927(.A1(new_n801), .A2(KEYINPUT53), .A3(new_n264), .ZN(new_n1128));
  OAI21_X1  g0928(.A(KEYINPUT53), .B1(new_n801), .B2(new_n264), .ZN(new_n1129));
  INV_X1    g0929(.A(G125), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1128), .B(new_n1129), .C1(new_n1130), .C2(new_n788), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n839), .B2(G137), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1125), .A2(new_n1127), .A3(new_n1132), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1123), .B(new_n1133), .C1(G159), .C2(new_n776), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n293), .B1(new_n839), .B2(G107), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n850), .A2(G68), .B1(G77), .B2(new_n776), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1135), .B(new_n1136), .C1(new_n568), .C2(new_n808), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n785), .A2(new_n479), .B1(new_n811), .B2(new_n788), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n799), .A2(new_n472), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n795), .A2(new_n815), .ZN(new_n1140));
  NOR4_X1   g0940(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .A4(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n773), .B1(new_n1134), .B2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1121), .A2(new_n833), .A3(new_n1122), .A4(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1119), .A2(new_n1120), .A3(new_n1143), .ZN(G378));
  AOI22_X1  g0944(.A1(new_n583), .A2(new_n784), .B1(new_n839), .B2(G97), .ZN(new_n1145));
  XOR2_X1   g0945(.A(new_n1145), .B(KEYINPUT114), .Z(new_n1146));
  AOI22_X1  g0946(.A1(new_n796), .A2(G116), .B1(G77), .B2(new_n802), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n850), .A2(G58), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  NOR4_X1   g0949(.A1(new_n1149), .A2(G41), .A3(new_n538), .A4(new_n1017), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1150), .B1(new_n549), .B2(new_n799), .C1(new_n815), .C2(new_n788), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT115), .ZN(new_n1152));
  OR2_X1    g0952(.A1(new_n1152), .A2(KEYINPUT58), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(KEYINPUT58), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n333), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n217), .B1(new_n1155), .B2(G41), .ZN(new_n1156));
  INV_X1    g0956(.A(G124), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n287), .B1(new_n788), .B2(new_n1157), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n839), .A2(G132), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n795), .A2(new_n1130), .B1(new_n264), .B2(new_n777), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT116), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n802), .A2(new_n1126), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n798), .A2(G128), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1159), .B(new_n1164), .C1(G137), .C2(new_n784), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT59), .ZN(new_n1166));
  AOI211_X1 g0966(.A(G33), .B(new_n1158), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1167), .B1(new_n1166), .B2(new_n1165), .C1(new_n842), .C2(new_n793), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1153), .A2(new_n1154), .A3(new_n1156), .A4(new_n1168), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n1169), .A2(new_n773), .B1(new_n217), .B2(new_n858), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n315), .A2(new_n317), .A3(new_n650), .ZN(new_n1171));
  XOR2_X1   g0971(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1172));
  OR2_X1    g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n320), .A2(new_n885), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1173), .A2(new_n1176), .A3(new_n1174), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n768), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1170), .A2(new_n833), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n928), .A2(KEYINPUT105), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n931), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n1184), .A2(new_n1185), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(new_n933), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n942), .A2(new_n1180), .A3(G330), .A4(new_n948), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n458), .A2(new_n877), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n879), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n458), .A2(new_n877), .A3(new_n879), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n866), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n562), .A2(new_n648), .A3(new_n700), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n758), .A2(new_n745), .A3(new_n700), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1195), .A2(new_n759), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1193), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n904), .B2(new_n912), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n948), .B(G330), .C1(new_n1198), .C2(KEYINPUT40), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1187), .A2(new_n914), .A3(new_n1188), .A4(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1188), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n935), .A2(new_n1203), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n1110), .A2(new_n1111), .A3(new_n1103), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n936), .A2(new_n1095), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1205), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT57), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n721), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1183), .B1(new_n1208), .B2(new_n1210), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1201), .A2(new_n1188), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT117), .ZN(new_n1213));
  OAI21_X1  g1013(.A(KEYINPUT118), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT118), .ZN(new_n1215));
  OAI21_X1  g1015(.A(KEYINPUT117), .B1(new_n935), .B2(new_n1215), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1214), .A2(new_n935), .B1(new_n1216), .B2(new_n1212), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n720), .A2(new_n1209), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1207), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1218), .B1(new_n1118), .B2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1217), .B1(new_n1220), .B2(new_n1004), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1211), .A2(new_n1221), .ZN(G375));
  NOR2_X1   g1022(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1223), .A2(new_n1090), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G107), .A2(new_n784), .B1(new_n839), .B2(new_n469), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1225), .A2(KEYINPUT119), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n501), .B1(new_n807), .B2(new_n788), .C1(new_n799), .C2(new_n815), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1225), .A2(KEYINPUT119), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n808), .A2(new_n479), .ZN(new_n1229));
  NOR4_X1   g1029(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1016), .B1(new_n583), .B2(new_n776), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1230), .B(new_n1231), .C1(new_n811), .C2(new_n795), .ZN(new_n1232));
  XOR2_X1   g1032(.A(new_n1232), .B(KEYINPUT120), .Z(new_n1233));
  AOI21_X1  g1033(.A(new_n838), .B1(new_n789), .B2(G128), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1148), .B(new_n1234), .C1(new_n785), .C2(new_n264), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G159), .B2(new_n845), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n798), .A2(G137), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n839), .A2(new_n1126), .B1(G50), .B2(new_n776), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(G132), .B2(new_n796), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n773), .B1(new_n1233), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n859), .A2(new_n202), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n882), .A2(new_n768), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1224), .B1(new_n833), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1223), .A2(new_n1207), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1246), .A2(new_n986), .A3(new_n1103), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1245), .A2(new_n1247), .ZN(G381));
  XOR2_X1   g1048(.A(G375), .B(KEYINPUT121), .Z(new_n1249));
  INV_X1    g1049(.A(G378), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1005), .A2(new_n1093), .A3(new_n1033), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1063), .A2(new_n1069), .A3(new_n836), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(G381), .A2(G384), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1249), .A2(new_n1250), .A3(new_n1253), .A4(new_n1254), .ZN(G407));
  INV_X1    g1055(.A(G213), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1256), .A2(G343), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1249), .A2(new_n1250), .A3(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1256), .B1(new_n1258), .B2(KEYINPUT122), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1259), .B(G407), .C1(KEYINPUT122), .C2(new_n1258), .ZN(G409));
  NAND2_X1  g1060(.A1(G387), .A2(G390), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1063), .A2(new_n1069), .A3(new_n836), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n836), .B1(new_n1063), .B2(new_n1069), .ZN(new_n1263));
  OAI21_X1  g1063(.A(KEYINPUT124), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(G393), .A2(G396), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT124), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1265), .A2(new_n1266), .A3(new_n1252), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1261), .A2(new_n1251), .A3(new_n1264), .A4(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1264), .A2(new_n1267), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1005), .A2(new_n1093), .A3(new_n1033), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1093), .B1(new_n1005), .B2(new_n1033), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1269), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n1268), .A2(new_n1272), .A3(KEYINPUT127), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT127), .B1(new_n1268), .B2(new_n1272), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  XOR2_X1   g1075(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1276));
  AOI21_X1  g1076(.A(new_n987), .B1(new_n1118), .B2(new_n1219), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1217), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1205), .A2(new_n1004), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1278), .A2(new_n1182), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1250), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1211), .A2(G378), .A3(new_n1221), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1257), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT60), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1246), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1223), .A2(KEYINPUT60), .A3(new_n1207), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1285), .A2(new_n720), .A3(new_n1103), .A4(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1287), .A2(G384), .A3(new_n1245), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(G384), .B1(new_n1287), .B2(new_n1245), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1276), .B1(new_n1283), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1257), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1211), .A2(G378), .A3(new_n1221), .ZN(new_n1294));
  AOI22_X1  g1094(.A1(new_n1277), .A2(new_n1217), .B1(new_n1004), .B2(new_n1205), .ZN(new_n1295));
  AOI21_X1  g1095(.A(G378), .B1(new_n1295), .B2(new_n1182), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1293), .B1(new_n1294), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT125), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1283), .A2(KEYINPUT125), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1291), .A2(KEYINPUT62), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1292), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1257), .A2(G2897), .ZN(new_n1304));
  XOR2_X1   g1104(.A(new_n1291), .B(new_n1304), .Z(new_n1305));
  NAND3_X1  g1105(.A1(new_n1299), .A2(new_n1305), .A3(new_n1300), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT61), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1275), .B1(new_n1303), .B2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1291), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT63), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(KEYINPUT61), .B1(new_n1301), .B2(new_n1312), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1291), .B(new_n1293), .C1(new_n1294), .C2(new_n1296), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1314), .A2(KEYINPUT123), .A3(new_n1311), .ZN(new_n1315));
  AOI21_X1  g1115(.A(KEYINPUT123), .B1(new_n1314), .B2(new_n1311), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1268), .A2(new_n1272), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1318), .B1(new_n1305), .B2(new_n1297), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1313), .A2(new_n1317), .A3(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1309), .A2(new_n1320), .ZN(G405));
  OAI21_X1  g1121(.A(new_n1291), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT127), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1318), .A2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1268), .A2(new_n1272), .A3(KEYINPUT127), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1324), .A2(new_n1310), .A3(new_n1325), .ZN(new_n1326));
  XNOR2_X1  g1126(.A(G375), .B(G378), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1322), .A2(new_n1326), .A3(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1327), .B1(new_n1322), .B2(new_n1326), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1328), .A2(new_n1329), .ZN(G402));
endmodule


