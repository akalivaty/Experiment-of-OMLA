

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809;

  AND2_X1 U380 ( .A1(n414), .A2(n413), .ZN(n412) );
  OR2_X1 U381 ( .A1(n455), .A2(n454), .ZN(n735) );
  INV_X1 U382 ( .A(G902), .ZN(n572) );
  XNOR2_X1 U383 ( .A(n366), .B(G469), .ZN(n556) );
  NAND2_X2 U384 ( .A1(n452), .A2(n450), .ZN(n449) );
  AND2_X2 U385 ( .A1(n436), .A2(n435), .ZN(n434) );
  XNOR2_X2 U386 ( .A(n498), .B(n497), .ZN(n570) );
  XNOR2_X2 U387 ( .A(G143), .B(KEYINPUT64), .ZN(n498) );
  INV_X1 U388 ( .A(KEYINPUT65), .ZN(n356) );
  NOR2_X1 U389 ( .A1(n698), .A2(n715), .ZN(n562) );
  AND2_X1 U390 ( .A1(n477), .A2(n374), .ZN(n475) );
  AND2_X1 U391 ( .A1(n363), .A2(n364), .ZN(n403) );
  AND2_X1 U392 ( .A1(n468), .A2(n467), .ZN(n466) );
  XNOR2_X1 U393 ( .A(n460), .B(n634), .ZN(n809) );
  AND2_X1 U394 ( .A1(n399), .A2(n395), .ZN(n638) );
  NAND2_X1 U395 ( .A1(n417), .A2(n369), .ZN(n410) );
  XNOR2_X1 U396 ( .A(n735), .B(KEYINPUT6), .ZN(n656) );
  NOR2_X1 U397 ( .A1(n434), .A2(n512), .ZN(n424) );
  AND2_X1 U398 ( .A1(n430), .A2(n429), .ZN(n371) );
  XNOR2_X1 U399 ( .A(n587), .B(n586), .ZN(n607) );
  OR2_X1 U400 ( .A1(n686), .A2(n431), .ZN(n430) );
  BUF_X1 U401 ( .A(n783), .Z(n361) );
  XNOR2_X1 U402 ( .A(n421), .B(n541), .ZN(n796) );
  AND2_X1 U403 ( .A1(n669), .A2(n482), .ZN(n448) );
  XNOR2_X1 U404 ( .A(n441), .B(G140), .ZN(n540) );
  XNOR2_X1 U405 ( .A(n483), .B(G116), .ZN(n484) );
  XNOR2_X1 U406 ( .A(G107), .B(G122), .ZN(n384) );
  XNOR2_X1 U407 ( .A(G116), .B(G134), .ZN(n563) );
  XNOR2_X1 U408 ( .A(KEYINPUT103), .B(KEYINPUT102), .ZN(n564) );
  XNOR2_X1 U409 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n380) );
  XNOR2_X1 U410 ( .A(KEYINPUT8), .B(KEYINPUT71), .ZN(n525) );
  OR2_X2 U411 ( .A1(n453), .A2(n356), .ZN(n452) );
  NAND2_X1 U412 ( .A1(n670), .A2(n668), .ZN(n357) );
  NAND2_X1 U413 ( .A1(n670), .A2(n668), .ZN(n616) );
  XNOR2_X1 U414 ( .A(n400), .B(n609), .ZN(n471) );
  XNOR2_X1 U415 ( .A(n357), .B(KEYINPUT85), .ZN(n358) );
  XNOR2_X1 U416 ( .A(n616), .B(KEYINPUT85), .ZN(n437) );
  INV_X1 U417 ( .A(n660), .ZN(n359) );
  XNOR2_X1 U418 ( .A(n556), .B(KEYINPUT1), .ZN(n591) );
  BUF_X1 U419 ( .A(n796), .Z(n360) );
  INV_X1 U420 ( .A(n474), .ZN(n362) );
  NAND2_X1 U421 ( .A1(n759), .A2(KEYINPUT34), .ZN(n363) );
  AND2_X1 U422 ( .A1(n420), .A2(n639), .ZN(n364) );
  XNOR2_X2 U423 ( .A(n480), .B(n494), .ZN(n783) );
  BUF_X1 U424 ( .A(n538), .Z(n365) );
  NOR2_X1 U425 ( .A1(n770), .A2(G902), .ZN(n366) );
  XNOR2_X1 U426 ( .A(KEYINPUT91), .B(KEYINPUT15), .ZN(n505) );
  INV_X1 U427 ( .A(n529), .ZN(n668) );
  INV_X1 U428 ( .A(G137), .ZN(n441) );
  XNOR2_X1 U429 ( .A(n783), .B(n546), .ZN(n418) );
  NOR2_X1 U430 ( .A1(n673), .A2(n457), .ZN(n454) );
  NAND2_X1 U431 ( .A1(n456), .A2(n459), .ZN(n455) );
  NAND2_X1 U432 ( .A1(n458), .A2(n572), .ZN(n457) );
  XNOR2_X1 U433 ( .A(n391), .B(n445), .ZN(n444) );
  INV_X1 U434 ( .A(KEYINPUT48), .ZN(n445) );
  NOR2_X1 U435 ( .A1(G953), .A2(G237), .ZN(n574) );
  INV_X1 U436 ( .A(KEYINPUT96), .ZN(n469) );
  XNOR2_X1 U437 ( .A(KEYINPUT5), .B(G137), .ZN(n549) );
  INV_X1 U438 ( .A(G146), .ZN(n548) );
  XNOR2_X1 U439 ( .A(G134), .B(G131), .ZN(n537) );
  NAND2_X1 U440 ( .A1(n508), .A2(n668), .ZN(n435) );
  INV_X1 U441 ( .A(KEYINPUT97), .ZN(n558) );
  INV_X1 U442 ( .A(KEYINPUT30), .ZN(n397) );
  NAND2_X2 U443 ( .A1(n728), .A2(n631), .ZN(n617) );
  NOR2_X1 U444 ( .A1(n617), .A2(n469), .ZN(n464) );
  XNOR2_X1 U445 ( .A(G128), .B(KEYINPUT83), .ZN(n521) );
  XNOR2_X1 U446 ( .A(G119), .B(G110), .ZN(n520) );
  NAND2_X1 U447 ( .A1(n388), .A2(n671), .ZN(n481) );
  XNOR2_X1 U448 ( .A(n390), .B(n389), .ZN(n388) );
  INV_X1 U449 ( .A(KEYINPUT86), .ZN(n389) );
  XNOR2_X1 U450 ( .A(n630), .B(n443), .ZN(n442) );
  INV_X1 U451 ( .A(KEYINPUT28), .ZN(n443) );
  XNOR2_X1 U452 ( .A(n633), .B(n632), .ZN(n760) );
  OR2_X1 U453 ( .A1(n359), .A2(KEYINPUT105), .ZN(n476) );
  XNOR2_X1 U454 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n500) );
  NAND2_X1 U455 ( .A1(n433), .A2(n432), .ZN(n431) );
  INV_X1 U456 ( .A(n668), .ZN(n432) );
  INV_X1 U457 ( .A(G237), .ZN(n506) );
  NOR2_X1 U458 ( .A1(n731), .A2(n732), .ZN(n536) );
  INV_X1 U459 ( .A(G472), .ZN(n458) );
  NAND2_X1 U460 ( .A1(G902), .A2(G472), .ZN(n459) );
  XNOR2_X1 U461 ( .A(KEYINPUT101), .B(KEYINPUT12), .ZN(n580) );
  XNOR2_X1 U462 ( .A(G131), .B(KEYINPUT99), .ZN(n581) );
  XNOR2_X1 U463 ( .A(n422), .B(n575), .ZN(n577) );
  XNOR2_X1 U464 ( .A(n576), .B(KEYINPUT11), .ZN(n422) );
  XNOR2_X1 U465 ( .A(G140), .B(KEYINPUT100), .ZN(n576) );
  XNOR2_X1 U466 ( .A(G143), .B(G113), .ZN(n578) );
  NAND2_X1 U467 ( .A1(G234), .A2(G237), .ZN(n513) );
  INV_X1 U468 ( .A(n760), .ZN(n741) );
  INV_X1 U469 ( .A(KEYINPUT104), .ZN(n406) );
  XNOR2_X1 U470 ( .A(n549), .B(n548), .ZN(n553) );
  XNOR2_X1 U471 ( .A(G107), .B(G104), .ZN(n496) );
  NAND2_X1 U472 ( .A1(n451), .A2(KEYINPUT65), .ZN(n450) );
  INV_X1 U473 ( .A(n669), .ZN(n451) );
  NOR2_X1 U474 ( .A1(n385), .A2(KEYINPUT34), .ZN(n419) );
  INV_X1 U475 ( .A(KEYINPUT31), .ZN(n560) );
  AND2_X1 U476 ( .A1(n396), .A2(n625), .ZN(n395) );
  XNOR2_X1 U477 ( .A(n617), .B(KEYINPUT107), .ZN(n399) );
  XNOR2_X1 U478 ( .A(n398), .B(n397), .ZN(n396) );
  NAND2_X1 U479 ( .A1(n367), .A2(n370), .ZN(n643) );
  AND2_X1 U480 ( .A1(n462), .A2(n470), .ZN(n698) );
  NAND2_X1 U481 ( .A1(n466), .A2(n463), .ZN(n462) );
  NAND2_X1 U482 ( .A1(n465), .A2(n464), .ZN(n463) );
  XOR2_X1 U483 ( .A(KEYINPUT62), .B(n673), .Z(n674) );
  INV_X2 U484 ( .A(G953), .ZN(n797) );
  XNOR2_X1 U485 ( .A(KEYINPUT16), .B(G122), .ZN(n494) );
  XNOR2_X1 U486 ( .A(n439), .B(n440), .ZN(n778) );
  XNOR2_X1 U487 ( .A(n528), .B(n527), .ZN(n439) );
  XNOR2_X1 U488 ( .A(n523), .B(n368), .ZN(n440) );
  XNOR2_X1 U489 ( .A(n686), .B(n689), .ZN(n690) );
  INV_X1 U490 ( .A(n481), .ZN(n726) );
  INV_X1 U491 ( .A(KEYINPUT42), .ZN(n634) );
  INV_X1 U492 ( .A(n643), .ZN(n712) );
  NAND2_X1 U493 ( .A1(n474), .A2(n473), .ZN(n472) );
  INV_X1 U494 ( .A(KEYINPUT105), .ZN(n473) );
  INV_X1 U495 ( .A(KEYINPUT60), .ZN(n489) );
  AND2_X1 U496 ( .A1(n417), .A2(n416), .ZN(n367) );
  XOR2_X1 U497 ( .A(n522), .B(n521), .Z(n368) );
  NOR2_X1 U498 ( .A1(n424), .A2(n411), .ZN(n369) );
  INV_X1 U499 ( .A(n557), .ZN(n728) );
  XNOR2_X1 U500 ( .A(n536), .B(KEYINPUT69), .ZN(n557) );
  AND2_X1 U501 ( .A1(n442), .A2(n631), .ZN(n370) );
  NAND2_X1 U502 ( .A1(n444), .A2(n667), .ZN(n723) );
  INV_X1 U503 ( .A(n735), .ZN(n470) );
  AND2_X1 U504 ( .A1(n392), .A2(n806), .ZN(n372) );
  AND2_X1 U505 ( .A1(n426), .A2(n425), .ZN(n373) );
  AND2_X1 U506 ( .A1(n476), .A2(n598), .ZN(n374) );
  XOR2_X1 U507 ( .A(KEYINPUT75), .B(KEYINPUT22), .Z(n375) );
  XOR2_X1 U508 ( .A(KEYINPUT108), .B(KEYINPUT40), .Z(n376) );
  XNOR2_X1 U509 ( .A(KEYINPUT59), .B(n684), .ZN(n377) );
  INV_X1 U510 ( .A(KEYINPUT65), .ZN(n482) );
  NOR2_X1 U511 ( .A1(n449), .A2(n446), .ZN(n378) );
  NOR2_X1 U512 ( .A1(n449), .A2(n446), .ZN(n379) );
  NOR2_X1 U513 ( .A1(n449), .A2(n446), .ZN(n777) );
  XNOR2_X1 U514 ( .A(n407), .B(n406), .ZN(n405) );
  INV_X1 U515 ( .A(G122), .ZN(n683) );
  NOR2_X1 U516 ( .A1(n408), .A2(n385), .ZN(n561) );
  XNOR2_X1 U517 ( .A(n559), .B(n558), .ZN(n408) );
  XOR2_X1 U518 ( .A(n380), .B(n564), .Z(n565) );
  NOR2_X1 U519 ( .A1(n434), .A2(n383), .ZN(n381) );
  NOR2_X1 U520 ( .A1(n381), .A2(n382), .ZN(n413) );
  AND2_X1 U521 ( .A1(KEYINPUT0), .A2(n518), .ZN(n382) );
  OR2_X1 U522 ( .A1(n512), .A2(n519), .ZN(n383) );
  XNOR2_X1 U523 ( .A(n623), .B(KEYINPUT38), .ZN(n744) );
  XOR2_X1 U524 ( .A(n384), .B(n563), .Z(n566) );
  NAND2_X1 U525 ( .A1(n412), .A2(n410), .ZN(n385) );
  NAND2_X1 U526 ( .A1(n412), .A2(n410), .ZN(n589) );
  NAND2_X1 U527 ( .A1(n403), .A2(n401), .ZN(n400) );
  NAND2_X1 U528 ( .A1(n735), .A2(n743), .ZN(n398) );
  NOR2_X1 U529 ( .A1(n748), .A2(n745), .ZN(n633) );
  XNOR2_X1 U530 ( .A(n418), .B(n504), .ZN(n686) );
  XNOR2_X1 U531 ( .A(n605), .B(KEYINPUT33), .ZN(n386) );
  NOR2_X1 U532 ( .A1(n591), .A2(n557), .ZN(n387) );
  XNOR2_X1 U533 ( .A(n605), .B(KEYINPUT33), .ZN(n759) );
  NAND2_X1 U534 ( .A1(n491), .A2(n692), .ZN(n490) );
  XNOR2_X1 U535 ( .A(n492), .B(n377), .ZN(n491) );
  INV_X1 U536 ( .A(n415), .ZN(n417) );
  NAND2_X1 U537 ( .A1(n415), .A2(KEYINPUT0), .ZN(n414) );
  NAND2_X1 U538 ( .A1(n409), .A2(n373), .ZN(n415) );
  OR2_X1 U539 ( .A1(n686), .A2(n427), .ZN(n426) );
  OR2_X2 U540 ( .A1(n606), .A2(n590), .ZN(n745) );
  INV_X1 U541 ( .A(n556), .ZN(n631) );
  NAND2_X1 U542 ( .A1(n402), .A2(n419), .ZN(n401) );
  NAND2_X1 U543 ( .A1(n447), .A2(n481), .ZN(n446) );
  NAND2_X1 U544 ( .A1(n453), .A2(n448), .ZN(n447) );
  NAND2_X1 U545 ( .A1(n672), .A2(KEYINPUT2), .ZN(n390) );
  NAND2_X1 U546 ( .A1(n393), .A2(n372), .ZN(n391) );
  XNOR2_X1 U547 ( .A(n652), .B(KEYINPUT76), .ZN(n392) );
  XNOR2_X1 U548 ( .A(n394), .B(KEYINPUT46), .ZN(n393) );
  NOR2_X2 U549 ( .A1(n805), .A2(n809), .ZN(n394) );
  INV_X1 U550 ( .A(n795), .ZN(n528) );
  XNOR2_X2 U551 ( .A(n524), .B(KEYINPUT10), .ZN(n795) );
  XNOR2_X2 U552 ( .A(G125), .B(G146), .ZN(n524) );
  INV_X1 U553 ( .A(n386), .ZN(n402) );
  XNOR2_X2 U554 ( .A(n404), .B(n375), .ZN(n601) );
  NOR2_X2 U555 ( .A1(n589), .A2(n405), .ZN(n404) );
  NOR2_X2 U556 ( .A1(n745), .A2(n732), .ZN(n407) );
  NAND2_X1 U557 ( .A1(n739), .A2(n408), .ZN(n740) );
  NAND2_X1 U558 ( .A1(n371), .A2(n434), .ZN(n409) );
  INV_X1 U559 ( .A(n424), .ZN(n416) );
  OR2_X1 U560 ( .A1(n518), .A2(KEYINPUT0), .ZN(n411) );
  NAND2_X1 U561 ( .A1(n385), .A2(KEYINPUT34), .ZN(n420) );
  XNOR2_X1 U562 ( .A(n421), .B(n555), .ZN(n673) );
  XNOR2_X2 U563 ( .A(n538), .B(n537), .ZN(n421) );
  XNOR2_X1 U564 ( .A(n796), .B(n547), .ZN(n770) );
  XNOR2_X1 U565 ( .A(n423), .B(n612), .ZN(n613) );
  NOR2_X2 U566 ( .A1(n471), .A2(n610), .ZN(n423) );
  NAND2_X1 U567 ( .A1(n510), .A2(n511), .ZN(n425) );
  NAND2_X1 U568 ( .A1(n428), .A2(n511), .ZN(n427) );
  INV_X1 U569 ( .A(n431), .ZN(n428) );
  NAND2_X1 U570 ( .A1(n434), .A2(n430), .ZN(n623) );
  NOR2_X1 U571 ( .A1(n510), .A2(n511), .ZN(n429) );
  INV_X1 U572 ( .A(n508), .ZN(n433) );
  NAND2_X1 U573 ( .A1(n686), .A2(n508), .ZN(n436) );
  NAND2_X1 U574 ( .A1(n437), .A2(n672), .ZN(n488) );
  NAND2_X1 U575 ( .A1(n358), .A2(n486), .ZN(n485) );
  XNOR2_X2 U576 ( .A(n438), .B(n533), .ZN(n731) );
  NAND2_X1 U577 ( .A1(n778), .A2(n572), .ZN(n438) );
  NAND2_X1 U578 ( .A1(n487), .A2(n485), .ZN(n453) );
  NAND2_X1 U579 ( .A1(n379), .A2(G475), .ZN(n492) );
  NAND2_X1 U580 ( .A1(n613), .A2(n614), .ZN(n615) );
  NAND2_X2 U581 ( .A1(n475), .A2(n472), .ZN(n685) );
  NAND2_X1 U582 ( .A1(n673), .A2(G472), .ZN(n456) );
  NAND2_X1 U583 ( .A1(n760), .A2(n370), .ZN(n460) );
  XNOR2_X2 U584 ( .A(n461), .B(n376), .ZN(n805) );
  NAND2_X1 U585 ( .A1(n663), .A2(n711), .ZN(n461) );
  XNOR2_X2 U586 ( .A(n624), .B(KEYINPUT39), .ZN(n663) );
  INV_X1 U587 ( .A(n385), .ZN(n465) );
  NAND2_X1 U588 ( .A1(n617), .A2(n469), .ZN(n467) );
  NAND2_X1 U589 ( .A1(n385), .A2(n469), .ZN(n468) );
  XNOR2_X1 U590 ( .A(n471), .B(n683), .ZN(G24) );
  INV_X1 U591 ( .A(n601), .ZN(n474) );
  NAND2_X1 U592 ( .A1(n601), .A2(n478), .ZN(n477) );
  AND2_X1 U593 ( .A1(n359), .A2(KEYINPUT105), .ZN(n478) );
  NAND2_X1 U594 ( .A1(n681), .A2(n685), .ZN(n610) );
  XNOR2_X2 U595 ( .A(n479), .B(n602), .ZN(n681) );
  NAND2_X1 U596 ( .A1(n601), .A2(n600), .ZN(n479) );
  XNOR2_X1 U597 ( .A(n480), .B(n554), .ZN(n555) );
  XNOR2_X2 U598 ( .A(n484), .B(n493), .ZN(n480) );
  XNOR2_X2 U599 ( .A(G113), .B(KEYINPUT73), .ZN(n483) );
  NOR2_X1 U600 ( .A1(n723), .A2(KEYINPUT84), .ZN(n486) );
  NAND2_X1 U601 ( .A1(n488), .A2(KEYINPUT84), .ZN(n487) );
  XNOR2_X1 U602 ( .A(n490), .B(n489), .ZN(G60) );
  XNOR2_X1 U603 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U604 ( .A(n553), .B(n552), .ZN(n554) );
  INV_X1 U605 ( .A(n511), .ZN(n512) );
  XNOR2_X1 U606 ( .A(n561), .B(n560), .ZN(n715) );
  XOR2_X1 U607 ( .A(KEYINPUT3), .B(G119), .Z(n493) );
  XNOR2_X1 U608 ( .A(KEYINPUT77), .B(G110), .ZN(n495) );
  XNOR2_X1 U609 ( .A(n496), .B(n495), .ZN(n784) );
  XNOR2_X1 U610 ( .A(KEYINPUT68), .B(G101), .ZN(n550) );
  XNOR2_X1 U611 ( .A(n784), .B(n550), .ZN(n546) );
  INV_X1 U612 ( .A(G128), .ZN(n497) );
  XNOR2_X2 U613 ( .A(n570), .B(KEYINPUT4), .ZN(n538) );
  NAND2_X1 U614 ( .A1(n797), .A2(G224), .ZN(n499) );
  XNOR2_X1 U615 ( .A(n499), .B(KEYINPUT92), .ZN(n502) );
  XNOR2_X1 U616 ( .A(n524), .B(n500), .ZN(n501) );
  XNOR2_X1 U617 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U618 ( .A(n365), .B(n503), .ZN(n504) );
  XNOR2_X1 U619 ( .A(n505), .B(n572), .ZN(n529) );
  NAND2_X1 U620 ( .A1(n572), .A2(n506), .ZN(n509) );
  NAND2_X1 U621 ( .A1(n509), .A2(G210), .ZN(n507) );
  XNOR2_X1 U622 ( .A(n507), .B(KEYINPUT80), .ZN(n508) );
  NAND2_X1 U623 ( .A1(n509), .A2(G214), .ZN(n743) );
  INV_X1 U624 ( .A(n743), .ZN(n510) );
  XNOR2_X1 U625 ( .A(KEYINPUT67), .B(KEYINPUT19), .ZN(n511) );
  XNOR2_X1 U626 ( .A(KEYINPUT14), .B(n513), .ZN(n515) );
  NAND2_X1 U627 ( .A1(G952), .A2(n515), .ZN(n757) );
  NOR2_X1 U628 ( .A1(n757), .A2(G953), .ZN(n514) );
  XNOR2_X1 U629 ( .A(n514), .B(KEYINPUT93), .ZN(n622) );
  NAND2_X1 U630 ( .A1(G902), .A2(n515), .ZN(n618) );
  INV_X1 U631 ( .A(n618), .ZN(n516) );
  NOR2_X1 U632 ( .A1(G898), .A2(n797), .ZN(n786) );
  NAND2_X1 U633 ( .A1(n516), .A2(n786), .ZN(n517) );
  AND2_X1 U634 ( .A1(n622), .A2(n517), .ZN(n518) );
  INV_X1 U635 ( .A(KEYINPUT0), .ZN(n519) );
  XNOR2_X1 U636 ( .A(n540), .B(n520), .ZN(n523) );
  XOR2_X1 U637 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n522) );
  NAND2_X1 U638 ( .A1(n797), .A2(G234), .ZN(n526) );
  XNOR2_X1 U639 ( .A(n526), .B(n525), .ZN(n567) );
  NAND2_X1 U640 ( .A1(G221), .A2(n567), .ZN(n527) );
  XOR2_X1 U641 ( .A(KEYINPUT95), .B(KEYINPUT25), .Z(n532) );
  NAND2_X1 U642 ( .A1(n529), .A2(G234), .ZN(n530) );
  XNOR2_X1 U643 ( .A(n530), .B(KEYINPUT20), .ZN(n534) );
  NAND2_X1 U644 ( .A1(n534), .A2(G217), .ZN(n531) );
  XNOR2_X1 U645 ( .A(n532), .B(n531), .ZN(n533) );
  AND2_X1 U646 ( .A1(n534), .A2(G221), .ZN(n535) );
  XNOR2_X1 U647 ( .A(n535), .B(KEYINPUT21), .ZN(n626) );
  INV_X1 U648 ( .A(n626), .ZN(n732) );
  INV_X1 U649 ( .A(KEYINPUT94), .ZN(n539) );
  XNOR2_X1 U650 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U651 ( .A(KEYINPUT78), .B(KEYINPUT79), .ZN(n544) );
  NAND2_X1 U652 ( .A1(G227), .A2(n797), .ZN(n542) );
  XNOR2_X1 U653 ( .A(G146), .B(n542), .ZN(n543) );
  XNOR2_X1 U654 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U655 ( .A(n546), .B(n545), .ZN(n547) );
  NAND2_X1 U656 ( .A1(n574), .A2(G210), .ZN(n551) );
  NOR2_X1 U657 ( .A1(n591), .A2(n557), .ZN(n604) );
  NAND2_X1 U658 ( .A1(n387), .A2(n735), .ZN(n559) );
  XNOR2_X1 U659 ( .A(n562), .B(KEYINPUT98), .ZN(n588) );
  XOR2_X1 U660 ( .A(n566), .B(n565), .Z(n569) );
  NAND2_X1 U661 ( .A1(G217), .A2(n567), .ZN(n568) );
  XNOR2_X1 U662 ( .A(n569), .B(n568), .ZN(n571) );
  XNOR2_X1 U663 ( .A(n570), .B(n571), .ZN(n775) );
  NAND2_X1 U664 ( .A1(n775), .A2(n572), .ZN(n573) );
  XNOR2_X1 U665 ( .A(n573), .B(G478), .ZN(n606) );
  NAND2_X1 U666 ( .A1(n574), .A2(G214), .ZN(n575) );
  XNOR2_X1 U667 ( .A(n577), .B(n795), .ZN(n585) );
  XNOR2_X1 U668 ( .A(n683), .B(G104), .ZN(n579) );
  XNOR2_X1 U669 ( .A(n579), .B(n578), .ZN(n583) );
  XNOR2_X1 U670 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U671 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U672 ( .A(n585), .B(n584), .ZN(n684) );
  OR2_X1 U673 ( .A1(n684), .A2(G902), .ZN(n587) );
  XNOR2_X1 U674 ( .A(G475), .B(KEYINPUT13), .ZN(n586) );
  AND2_X1 U675 ( .A1(n606), .A2(n607), .ZN(n706) );
  INV_X1 U676 ( .A(n706), .ZN(n718) );
  OR2_X1 U677 ( .A1(n606), .A2(n607), .ZN(n716) );
  AND2_X1 U678 ( .A1(n718), .A2(n716), .ZN(n749) );
  NOR2_X1 U679 ( .A1(n588), .A2(n749), .ZN(n597) );
  INV_X1 U680 ( .A(n607), .ZN(n590) );
  INV_X1 U681 ( .A(n591), .ZN(n660) );
  INV_X1 U682 ( .A(n731), .ZN(n628) );
  NAND2_X1 U683 ( .A1(n656), .A2(n628), .ZN(n592) );
  NOR2_X1 U684 ( .A1(n660), .A2(n592), .ZN(n593) );
  NAND2_X1 U685 ( .A1(n362), .A2(n593), .ZN(n696) );
  INV_X1 U686 ( .A(KEYINPUT74), .ZN(n594) );
  NAND2_X1 U687 ( .A1(n594), .A2(KEYINPUT44), .ZN(n595) );
  NAND2_X1 U688 ( .A1(n696), .A2(n595), .ZN(n596) );
  NOR2_X1 U689 ( .A1(n597), .A2(n596), .ZN(n614) );
  NOR2_X1 U690 ( .A1(n628), .A2(n735), .ZN(n598) );
  NAND2_X1 U691 ( .A1(n656), .A2(n731), .ZN(n599) );
  NOR2_X1 U692 ( .A1(n359), .A2(n599), .ZN(n600) );
  XNOR2_X1 U693 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n602) );
  INV_X1 U694 ( .A(n656), .ZN(n603) );
  AND2_X2 U695 ( .A1(n604), .A2(n603), .ZN(n605) );
  INV_X1 U696 ( .A(n606), .ZN(n608) );
  NOR2_X1 U697 ( .A1(n608), .A2(n607), .ZN(n639) );
  XOR2_X1 U698 ( .A(KEYINPUT87), .B(KEYINPUT35), .Z(n609) );
  INV_X1 U699 ( .A(KEYINPUT44), .ZN(n611) );
  NAND2_X1 U700 ( .A1(n611), .A2(KEYINPUT74), .ZN(n612) );
  XNOR2_X2 U701 ( .A(n615), .B(KEYINPUT45), .ZN(n670) );
  NOR2_X1 U702 ( .A1(G900), .A2(n618), .ZN(n619) );
  NAND2_X1 U703 ( .A1(G953), .A2(n619), .ZN(n620) );
  XNOR2_X1 U704 ( .A(KEYINPUT106), .B(n620), .ZN(n621) );
  NAND2_X1 U705 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n638), .A2(n744), .ZN(n624) );
  INV_X1 U707 ( .A(n716), .ZN(n711) );
  AND2_X1 U708 ( .A1(n626), .A2(n625), .ZN(n627) );
  XOR2_X1 U709 ( .A(KEYINPUT72), .B(n627), .Z(n654) );
  NOR2_X1 U710 ( .A1(n654), .A2(n628), .ZN(n629) );
  NAND2_X1 U711 ( .A1(n629), .A2(n735), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n744), .A2(n743), .ZN(n748) );
  XNOR2_X1 U713 ( .A(KEYINPUT41), .B(KEYINPUT109), .ZN(n632) );
  INV_X1 U714 ( .A(KEYINPUT82), .ZN(n644) );
  INV_X1 U715 ( .A(KEYINPUT70), .ZN(n635) );
  OR2_X1 U716 ( .A1(n749), .A2(n635), .ZN(n645) );
  NOR2_X1 U717 ( .A1(n643), .A2(n645), .ZN(n636) );
  NOR2_X1 U718 ( .A1(n644), .A2(n636), .ZN(n637) );
  NOR2_X1 U719 ( .A1(KEYINPUT47), .A2(n637), .ZN(n651) );
  INV_X1 U720 ( .A(n638), .ZN(n641) );
  INV_X1 U721 ( .A(n623), .ZN(n658) );
  NAND2_X1 U722 ( .A1(n639), .A2(n658), .ZN(n640) );
  NOR2_X1 U723 ( .A1(n641), .A2(n640), .ZN(n710) );
  NOR2_X1 U724 ( .A1(n749), .A2(KEYINPUT82), .ZN(n642) );
  NOR2_X1 U725 ( .A1(n710), .A2(n642), .ZN(n649) );
  NAND2_X1 U726 ( .A1(KEYINPUT82), .A2(n645), .ZN(n646) );
  NAND2_X1 U727 ( .A1(n712), .A2(n646), .ZN(n647) );
  NAND2_X1 U728 ( .A1(KEYINPUT47), .A2(n647), .ZN(n648) );
  NAND2_X1 U729 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U730 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U731 ( .A1(n731), .A2(n743), .ZN(n653) );
  NOR2_X1 U732 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U733 ( .A1(n655), .A2(n711), .ZN(n657) );
  NOR2_X1 U734 ( .A1(n657), .A2(n656), .ZN(n664) );
  NAND2_X1 U735 ( .A1(n664), .A2(n658), .ZN(n659) );
  XOR2_X1 U736 ( .A(n659), .B(KEYINPUT36), .Z(n661) );
  NAND2_X1 U737 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U738 ( .A(n662), .B(KEYINPUT110), .ZN(n806) );
  NAND2_X1 U739 ( .A1(n663), .A2(n706), .ZN(n722) );
  NAND2_X1 U740 ( .A1(n664), .A2(n359), .ZN(n665) );
  XNOR2_X1 U741 ( .A(n665), .B(KEYINPUT43), .ZN(n666) );
  NAND2_X1 U742 ( .A1(n666), .A2(n623), .ZN(n682) );
  AND2_X1 U743 ( .A1(n722), .A2(n682), .ZN(n667) );
  NAND2_X1 U744 ( .A1(n668), .A2(KEYINPUT2), .ZN(n669) );
  BUF_X1 U745 ( .A(n670), .Z(n671) );
  INV_X1 U746 ( .A(n671), .ZN(n724) );
  INV_X1 U747 ( .A(n723), .ZN(n672) );
  NAND2_X1 U748 ( .A1(n777), .A2(G472), .ZN(n675) );
  XNOR2_X1 U749 ( .A(n675), .B(n674), .ZN(n678) );
  INV_X1 U750 ( .A(G952), .ZN(n676) );
  NAND2_X1 U751 ( .A1(n676), .A2(G953), .ZN(n677) );
  XNOR2_X1 U752 ( .A(n677), .B(KEYINPUT90), .ZN(n692) );
  NAND2_X1 U753 ( .A1(n678), .A2(n692), .ZN(n680) );
  XOR2_X1 U754 ( .A(KEYINPUT63), .B(KEYINPUT111), .Z(n679) );
  XNOR2_X1 U755 ( .A(n680), .B(n679), .ZN(G57) );
  XNOR2_X1 U756 ( .A(n681), .B(G119), .ZN(G21) );
  XNOR2_X1 U757 ( .A(n682), .B(G140), .ZN(G42) );
  INV_X1 U758 ( .A(n692), .ZN(n782) );
  XNOR2_X1 U759 ( .A(n685), .B(G110), .ZN(G12) );
  NAND2_X1 U760 ( .A1(n777), .A2(G210), .ZN(n691) );
  XNOR2_X1 U761 ( .A(KEYINPUT89), .B(KEYINPUT54), .ZN(n688) );
  XNOR2_X1 U762 ( .A(KEYINPUT55), .B(KEYINPUT81), .ZN(n687) );
  XNOR2_X1 U763 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U764 ( .A(n691), .B(n690), .ZN(n693) );
  NAND2_X1 U765 ( .A1(n693), .A2(n692), .ZN(n695) );
  XOR2_X1 U766 ( .A(KEYINPUT88), .B(KEYINPUT56), .Z(n694) );
  XNOR2_X1 U767 ( .A(n695), .B(n694), .ZN(G51) );
  XNOR2_X1 U768 ( .A(n696), .B(G101), .ZN(n697) );
  XNOR2_X1 U769 ( .A(KEYINPUT112), .B(n697), .ZN(G3) );
  INV_X1 U770 ( .A(n698), .ZN(n703) );
  NOR2_X1 U771 ( .A1(n703), .A2(n716), .ZN(n700) );
  XNOR2_X1 U772 ( .A(G104), .B(KEYINPUT113), .ZN(n699) );
  XNOR2_X1 U773 ( .A(n700), .B(n699), .ZN(G6) );
  XOR2_X1 U774 ( .A(KEYINPUT26), .B(KEYINPUT114), .Z(n702) );
  XNOR2_X1 U775 ( .A(G107), .B(KEYINPUT27), .ZN(n701) );
  XNOR2_X1 U776 ( .A(n702), .B(n701), .ZN(n705) );
  NOR2_X1 U777 ( .A1(n703), .A2(n718), .ZN(n704) );
  XOR2_X1 U778 ( .A(n705), .B(n704), .Z(G9) );
  XOR2_X1 U779 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n708) );
  NAND2_X1 U780 ( .A1(n712), .A2(n706), .ZN(n707) );
  XNOR2_X1 U781 ( .A(n708), .B(n707), .ZN(n709) );
  XOR2_X1 U782 ( .A(G128), .B(n709), .Z(G30) );
  XOR2_X1 U783 ( .A(G143), .B(n710), .Z(G45) );
  NAND2_X1 U784 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U785 ( .A(n713), .B(KEYINPUT116), .ZN(n714) );
  XNOR2_X1 U786 ( .A(G146), .B(n714), .ZN(G48) );
  INV_X1 U787 ( .A(n715), .ZN(n719) );
  NOR2_X1 U788 ( .A1(n719), .A2(n716), .ZN(n717) );
  XOR2_X1 U789 ( .A(G113), .B(n717), .Z(G15) );
  NOR2_X1 U790 ( .A1(n719), .A2(n718), .ZN(n721) );
  XNOR2_X1 U791 ( .A(G116), .B(KEYINPUT117), .ZN(n720) );
  XNOR2_X1 U792 ( .A(n721), .B(n720), .ZN(G18) );
  XNOR2_X1 U793 ( .A(G134), .B(n722), .ZN(G36) );
  NOR2_X1 U794 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U795 ( .A1(n725), .A2(KEYINPUT2), .ZN(n727) );
  NOR2_X1 U796 ( .A1(n727), .A2(n726), .ZN(n764) );
  NAND2_X1 U797 ( .A1(n359), .A2(n557), .ZN(n730) );
  XNOR2_X1 U798 ( .A(KEYINPUT50), .B(KEYINPUT120), .ZN(n729) );
  XNOR2_X1 U799 ( .A(n730), .B(n729), .ZN(n738) );
  NAND2_X1 U800 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U801 ( .A(n733), .B(KEYINPUT119), .ZN(n734) );
  XNOR2_X1 U802 ( .A(KEYINPUT49), .B(n734), .ZN(n736) );
  AND2_X1 U803 ( .A1(n736), .A2(n470), .ZN(n737) );
  NAND2_X1 U804 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U805 ( .A(KEYINPUT51), .B(n740), .ZN(n742) );
  NOR2_X1 U806 ( .A1(n742), .A2(n741), .ZN(n754) );
  NOR2_X1 U807 ( .A1(n744), .A2(n743), .ZN(n746) );
  NOR2_X1 U808 ( .A1(n746), .A2(n745), .ZN(n747) );
  XOR2_X1 U809 ( .A(KEYINPUT121), .B(n747), .Z(n751) );
  NOR2_X1 U810 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U811 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U812 ( .A1(n386), .A2(n752), .ZN(n753) );
  NOR2_X1 U813 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U814 ( .A(n755), .B(KEYINPUT52), .ZN(n756) );
  NOR2_X1 U815 ( .A1(n757), .A2(n756), .ZN(n758) );
  XOR2_X1 U816 ( .A(KEYINPUT122), .B(n758), .Z(n762) );
  NAND2_X1 U817 ( .A1(n402), .A2(n760), .ZN(n761) );
  NAND2_X1 U818 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U819 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U820 ( .A(n765), .B(KEYINPUT123), .ZN(n766) );
  NOR2_X1 U821 ( .A1(G953), .A2(n766), .ZN(n767) );
  XNOR2_X1 U822 ( .A(KEYINPUT53), .B(n767), .ZN(G75) );
  NAND2_X1 U823 ( .A1(n379), .A2(G469), .ZN(n772) );
  XOR2_X1 U824 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n768) );
  XNOR2_X1 U825 ( .A(n768), .B(KEYINPUT124), .ZN(n769) );
  XNOR2_X1 U826 ( .A(n770), .B(n769), .ZN(n771) );
  XNOR2_X1 U827 ( .A(n772), .B(n771), .ZN(n773) );
  NOR2_X1 U828 ( .A1(n782), .A2(n773), .ZN(G54) );
  NAND2_X1 U829 ( .A1(n378), .A2(G478), .ZN(n774) );
  XOR2_X1 U830 ( .A(n775), .B(n774), .Z(n776) );
  NOR2_X1 U831 ( .A1(n782), .A2(n776), .ZN(G63) );
  NAND2_X1 U832 ( .A1(n378), .A2(G217), .ZN(n780) );
  XNOR2_X1 U833 ( .A(n778), .B(KEYINPUT125), .ZN(n779) );
  XNOR2_X1 U834 ( .A(n780), .B(n779), .ZN(n781) );
  NOR2_X1 U835 ( .A1(n782), .A2(n781), .ZN(G66) );
  XOR2_X1 U836 ( .A(G101), .B(n784), .Z(n785) );
  XNOR2_X1 U837 ( .A(n361), .B(n785), .ZN(n787) );
  NOR2_X1 U838 ( .A1(n787), .A2(n786), .ZN(n794) );
  NAND2_X1 U839 ( .A1(n671), .A2(n797), .ZN(n791) );
  NAND2_X1 U840 ( .A1(G953), .A2(G224), .ZN(n788) );
  XNOR2_X1 U841 ( .A(KEYINPUT61), .B(n788), .ZN(n789) );
  NAND2_X1 U842 ( .A1(n789), .A2(G898), .ZN(n790) );
  NAND2_X1 U843 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U844 ( .A(n792), .B(KEYINPUT126), .ZN(n793) );
  XNOR2_X1 U845 ( .A(n794), .B(n793), .ZN(G69) );
  XNOR2_X1 U846 ( .A(n360), .B(n795), .ZN(n799) );
  XNOR2_X1 U847 ( .A(n723), .B(n799), .ZN(n798) );
  NAND2_X1 U848 ( .A1(n798), .A2(n797), .ZN(n803) );
  XNOR2_X1 U849 ( .A(n799), .B(G227), .ZN(n800) );
  NAND2_X1 U850 ( .A1(n800), .A2(G900), .ZN(n801) );
  NAND2_X1 U851 ( .A1(n801), .A2(G953), .ZN(n802) );
  NAND2_X1 U852 ( .A1(n803), .A2(n802), .ZN(n804) );
  XOR2_X1 U853 ( .A(KEYINPUT127), .B(n804), .Z(G72) );
  XOR2_X1 U854 ( .A(G131), .B(n805), .Z(G33) );
  XOR2_X1 U855 ( .A(KEYINPUT37), .B(KEYINPUT118), .Z(n808) );
  XNOR2_X1 U856 ( .A(G125), .B(n806), .ZN(n807) );
  XNOR2_X1 U857 ( .A(n808), .B(n807), .ZN(G27) );
  XOR2_X1 U858 ( .A(G137), .B(n809), .Z(G39) );
endmodule

