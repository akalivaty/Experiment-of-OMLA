//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0 1 0 0 1 0 0 0 0 0 0 1 1 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n826, new_n827, new_n828,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(G1gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT91), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n202), .B1(new_n206), .B2(G1gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n205), .A2(new_n208), .A3(G8gat), .ZN(new_n209));
  INV_X1    g008(.A(G8gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n203), .B(new_n207), .C1(new_n204), .C2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  XOR2_X1   g012(.A(G43gat), .B(G50gat), .Z(new_n214));
  INV_X1    g013(.A(G36gat), .ZN(new_n215));
  AND2_X1   g014(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G29gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n219), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n214), .B1(new_n221), .B2(KEYINPUT15), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n222), .B1(KEYINPUT15), .B2(new_n221), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(KEYINPUT15), .A3(new_n214), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT17), .B1(new_n225), .B2(KEYINPUT90), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT90), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT17), .ZN(new_n228));
  AOI211_X1 g027(.A(new_n227), .B(new_n228), .C1(new_n223), .C2(new_n224), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n213), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G229gat), .A2(G233gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n225), .A2(new_n212), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT18), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n230), .A2(KEYINPUT18), .A3(new_n231), .A4(new_n232), .ZN(new_n236));
  OR3_X1    g035(.A1(new_n225), .A2(new_n212), .A3(KEYINPUT92), .ZN(new_n237));
  OAI21_X1  g036(.A(KEYINPUT92), .B1(new_n225), .B2(new_n212), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(new_n232), .A3(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n231), .B(KEYINPUT13), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n235), .A2(new_n236), .A3(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G113gat), .B(G141gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(G197gat), .ZN(new_n244));
  XOR2_X1   g043(.A(KEYINPUT11), .B(G169gat), .Z(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(KEYINPUT12), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n242), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n235), .A2(new_n247), .A3(new_n236), .A4(new_n241), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT22), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT76), .B(G218gat), .ZN(new_n254));
  INV_X1    g053(.A(G211gat), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G197gat), .B(G204gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G211gat), .B(G218gat), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n256), .A2(new_n257), .A3(new_n259), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G148gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(G141gat), .ZN(new_n265));
  XOR2_X1   g064(.A(KEYINPUT80), .B(G141gat), .Z(new_n266));
  OAI21_X1  g065(.A(new_n265), .B1(new_n266), .B2(new_n264), .ZN(new_n267));
  XOR2_X1   g066(.A(G155gat), .B(G162gat), .Z(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G155gat), .A2(G162gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT2), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n267), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G141gat), .B(G148gat), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT79), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n271), .B1(new_n273), .B2(new_n274), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n268), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AND2_X1   g076(.A1(new_n272), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT3), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT29), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n263), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n263), .A2(new_n281), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n278), .B1(new_n283), .B2(new_n279), .ZN(new_n284));
  INV_X1    g083(.A(G228gat), .ZN(new_n285));
  INV_X1    g084(.A(G233gat), .ZN(new_n286));
  OAI22_X1  g085(.A1(new_n282), .A2(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(KEYINPUT86), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n263), .B(KEYINPUT77), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT29), .B1(new_n278), .B2(new_n279), .ZN(new_n290));
  OR2_X1    g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n285), .A2(new_n286), .ZN(new_n292));
  INV_X1    g091(.A(new_n284), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n291), .A2(KEYINPUT87), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT87), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n292), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n289), .A2(new_n290), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G22gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n288), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n300), .B1(new_n288), .B2(new_n299), .ZN(new_n303));
  OAI21_X1  g102(.A(G78gat), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n303), .ZN(new_n305));
  INV_X1    g104(.A(G78gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(new_n306), .A3(new_n301), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT31), .B(G50gat), .ZN(new_n308));
  INV_X1    g107(.A(G106gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n304), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n310), .B1(new_n304), .B2(new_n307), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(G169gat), .A2(G176gat), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n314), .B1(KEYINPUT23), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT25), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G183gat), .ZN(new_n321));
  INV_X1    g120(.A(G190gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n320), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT23), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n314), .B(KEYINPUT66), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n318), .B(new_n325), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(KEYINPUT67), .ZN(new_n329));
  INV_X1    g128(.A(new_n314), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n330), .A2(new_n326), .ZN(new_n331));
  OR2_X1    g130(.A1(new_n331), .A2(new_n316), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT64), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n319), .B(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n334), .A2(new_n323), .A3(new_n324), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n332), .B1(new_n335), .B2(KEYINPUT65), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT65), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n334), .A2(new_n337), .A3(new_n323), .A4(new_n324), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT25), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT27), .B(G183gat), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT28), .B1(new_n340), .B2(new_n322), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n341), .B(KEYINPUT69), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n340), .B(KEYINPUT70), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n343), .A2(KEYINPUT28), .A3(new_n322), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT26), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n315), .B(new_n346), .C1(new_n327), .C2(KEYINPUT26), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n347), .B1(new_n321), .B2(new_n322), .ZN(new_n348));
  OAI22_X1  g147(.A1(new_n329), .A2(new_n339), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(G226gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n350), .A2(new_n286), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n351), .A2(KEYINPUT29), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n317), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT67), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n328), .B(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n355), .A2(new_n357), .A3(KEYINPUT68), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT68), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n359), .B1(new_n329), .B2(new_n339), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n345), .A2(new_n348), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n351), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n353), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n263), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n349), .A2(new_n365), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n368), .B1(new_n364), .B2(new_n352), .ZN(new_n369));
  INV_X1    g168(.A(new_n289), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  XOR2_X1   g170(.A(G8gat), .B(G36gat), .Z(new_n372));
  XNOR2_X1  g171(.A(new_n372), .B(KEYINPUT78), .ZN(new_n373));
  XNOR2_X1  g172(.A(G64gat), .B(G92gat), .ZN(new_n374));
  XOR2_X1   g173(.A(new_n373), .B(new_n374), .Z(new_n375));
  NAND3_X1  g174(.A1(new_n367), .A2(new_n371), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT30), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n367), .A2(new_n371), .A3(KEYINPUT30), .A4(new_n375), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n367), .A2(new_n371), .ZN(new_n380));
  INV_X1    g179(.A(new_n375), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n378), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G113gat), .B(G120gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n384), .A2(KEYINPUT1), .ZN(new_n385));
  XOR2_X1   g184(.A(G127gat), .B(G134gat), .Z(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n278), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n388), .A2(KEYINPUT4), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT4), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n390), .B1(new_n278), .B2(new_n387), .ZN(new_n391));
  OR3_X1    g190(.A1(new_n389), .A2(KEYINPUT83), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(G225gat), .A2(G233gat), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n272), .A2(new_n277), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n387), .B1(new_n395), .B2(KEYINPUT3), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n394), .B1(new_n280), .B2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT81), .B(KEYINPUT5), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n389), .A2(KEYINPUT83), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n392), .A2(new_n397), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n397), .B1(new_n389), .B2(new_n391), .ZN(new_n401));
  INV_X1    g200(.A(new_n387), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n395), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n398), .B1(new_n404), .B2(new_n394), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n401), .A2(KEYINPUT82), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT82), .B1(new_n401), .B2(new_n405), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n400), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G1gat), .B(G29gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(KEYINPUT0), .ZN(new_n410));
  XNOR2_X1  g209(.A(G57gat), .B(G85gat), .ZN(new_n411));
  XOR2_X1   g210(.A(new_n410), .B(new_n411), .Z(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n408), .A2(KEYINPUT6), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT85), .ZN(new_n415));
  OR2_X1    g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n415), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n400), .B(new_n412), .C1(new_n406), .C2(new_n407), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT6), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OR2_X1    g220(.A1(new_n421), .A2(KEYINPUT84), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n408), .A2(new_n413), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(KEYINPUT84), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n383), .B1(new_n418), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n362), .B1(new_n358), .B2(new_n360), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n427), .A2(new_n387), .ZN(new_n428));
  AOI211_X1 g227(.A(new_n402), .B(new_n362), .C1(new_n358), .C2(new_n360), .ZN(new_n429));
  OAI211_X1 g228(.A(G227gat), .B(G233gat), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT32), .ZN(new_n431));
  XOR2_X1   g230(.A(KEYINPUT71), .B(KEYINPUT33), .Z(new_n432));
  NAND2_X1  g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(G15gat), .B(G43gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n434), .B(G99gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(KEYINPUT72), .B(G71gat), .ZN(new_n436));
  XOR2_X1   g235(.A(new_n435), .B(new_n436), .Z(new_n437));
  NAND3_X1  g236(.A1(new_n431), .A2(new_n433), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT75), .ZN(new_n439));
  INV_X1    g238(.A(new_n437), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n430), .B(KEYINPUT32), .C1(new_n432), .C2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n438), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n439), .B1(new_n438), .B2(new_n441), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n364), .A2(new_n402), .ZN(new_n445));
  NAND2_X1  g244(.A1(G227gat), .A2(G233gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n427), .A2(new_n387), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  XOR2_X1   g247(.A(KEYINPUT73), .B(KEYINPUT34), .Z(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT74), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT74), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n448), .A2(new_n452), .A3(new_n449), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n448), .A2(KEYINPUT34), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n443), .A2(new_n444), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n438), .A2(new_n441), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n455), .B1(new_n451), .B2(new_n453), .ZN(new_n460));
  NOR3_X1   g259(.A1(new_n459), .A2(new_n460), .A3(KEYINPUT75), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n313), .B(new_n426), .C1(new_n458), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT35), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n459), .A2(KEYINPUT75), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n464), .A2(new_n442), .A3(new_n460), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n457), .A2(new_n439), .A3(new_n438), .A4(new_n441), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n423), .A2(new_n420), .A3(new_n419), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n416), .A2(new_n417), .A3(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n469), .A2(KEYINPUT35), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT88), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n383), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n378), .A2(new_n382), .A3(KEYINPUT88), .A4(new_n379), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n467), .A2(new_n313), .A3(new_n470), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n463), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n376), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT37), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n375), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n479), .B1(new_n380), .B2(new_n381), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  OAI22_X1  g280(.A1(new_n263), .A2(new_n366), .B1(new_n369), .B2(new_n370), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT38), .B1(new_n482), .B2(KEYINPUT37), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n477), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n478), .B1(new_n367), .B2(new_n371), .ZN(new_n485));
  OAI211_X1 g284(.A(KEYINPUT89), .B(KEYINPUT38), .C1(new_n480), .C2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n380), .A2(KEYINPUT37), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n375), .B1(new_n367), .B2(new_n371), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n488), .B1(new_n489), .B2(new_n479), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT89), .B1(new_n490), .B2(KEYINPUT38), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n469), .B(new_n484), .C1(new_n487), .C2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT40), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n280), .A2(new_n396), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n392), .A2(new_n494), .A3(new_n399), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n394), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n388), .A2(new_n393), .A3(new_n403), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n496), .A2(KEYINPUT39), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n412), .B1(new_n496), .B2(KEYINPUT39), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n493), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n423), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n498), .A2(new_n499), .A3(new_n493), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n503), .A2(new_n472), .A3(new_n473), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n492), .A2(new_n313), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n304), .A2(new_n307), .ZN(new_n506));
  INV_X1    g305(.A(new_n310), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n304), .A2(new_n307), .A3(new_n310), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n418), .A2(new_n425), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n510), .B1(new_n512), .B2(new_n383), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n465), .A2(KEYINPUT36), .A3(new_n466), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT36), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n467), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n505), .A2(new_n513), .A3(new_n514), .A4(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n252), .B1(new_n476), .B2(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(G120gat), .B(G148gat), .Z(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(KEYINPUT102), .ZN(new_n520));
  XNOR2_X1  g319(.A(G176gat), .B(G204gat), .ZN(new_n521));
  XOR2_X1   g320(.A(new_n520), .B(new_n521), .Z(new_n522));
  INV_X1    g321(.A(G230gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n523), .A2(new_n286), .ZN(new_n524));
  XOR2_X1   g323(.A(KEYINPUT100), .B(KEYINPUT10), .Z(new_n525));
  XNOR2_X1  g324(.A(G57gat), .B(G64gat), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(G71gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(new_n306), .ZN(new_n529));
  NAND2_X1  g328(.A1(G71gat), .A2(G78gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT9), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n527), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n530), .B(new_n529), .C1(new_n526), .C2(new_n532), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(G99gat), .A2(G106gat), .ZN(new_n538));
  INV_X1    g337(.A(G85gat), .ZN(new_n539));
  INV_X1    g338(.A(G92gat), .ZN(new_n540));
  AOI22_X1  g339(.A1(KEYINPUT8), .A2(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT7), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT95), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT95), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT7), .ZN(new_n545));
  AND2_X1   g344(.A1(G85gat), .A2(G92gat), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n543), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n546), .B1(new_n543), .B2(new_n545), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n541), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g348(.A1(G99gat), .A2(G106gat), .ZN(new_n550));
  NOR2_X1   g349(.A1(G99gat), .A2(G106gat), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT96), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(G99gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(new_n309), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT96), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n554), .A2(new_n555), .A3(new_n538), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n549), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G85gat), .A2(G92gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n544), .A2(KEYINPUT7), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n542), .A2(KEYINPUT95), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n543), .A2(new_n545), .A3(new_n546), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI22_X1  g363(.A1(new_n564), .A2(new_n541), .B1(new_n552), .B2(new_n556), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n537), .B1(new_n558), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n557), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n552), .A2(new_n556), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n568), .A2(new_n564), .A3(new_n541), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n567), .A2(new_n569), .A3(new_n536), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n566), .A2(KEYINPUT99), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n567), .A2(new_n569), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT99), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(new_n573), .A3(new_n537), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n525), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT101), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n536), .B1(new_n567), .B2(new_n569), .ZN(new_n577));
  AOI22_X1  g376(.A1(new_n575), .A2(new_n576), .B1(KEYINPUT10), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n525), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n570), .A2(KEYINPUT99), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n580), .A2(new_n577), .ZN(new_n581));
  INV_X1    g380(.A(new_n574), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n579), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT101), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n524), .B1(new_n578), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n571), .A2(new_n524), .A3(new_n574), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n522), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n524), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n576), .B(new_n579), .C1(new_n581), .C2(new_n582), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n577), .A2(KEYINPUT10), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n575), .A2(new_n576), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n589), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n522), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n594), .A2(new_n586), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n588), .A2(new_n596), .A3(KEYINPUT103), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT103), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n598), .B(new_n522), .C1(new_n585), .C2(new_n587), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G232gat), .A2(G233gat), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT41), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n604), .B1(new_n225), .B2(new_n572), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT97), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n569), .B(new_n567), .C1(new_n226), .C2(new_n229), .ZN(new_n607));
  XNOR2_X1  g406(.A(G134gat), .B(G162gat), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  AND3_X1   g408(.A1(new_n606), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n609), .B1(new_n606), .B2(new_n607), .ZN(new_n611));
  XOR2_X1   g410(.A(G190gat), .B(G218gat), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT98), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n602), .A2(new_n603), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT94), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n613), .B(new_n615), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  OR3_X1    g416(.A1(new_n610), .A2(new_n611), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n617), .B1(new_n610), .B2(new_n611), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT21), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n536), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G127gat), .B(G155gat), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n622), .B(new_n623), .Z(new_n624));
  AOI21_X1  g423(.A(new_n212), .B1(KEYINPUT21), .B2(new_n537), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G231gat), .A2(G233gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT93), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G183gat), .B(G211gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n626), .A2(new_n632), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n601), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n518), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(new_n511), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT104), .B(G1gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(G1324gat));
  INV_X1    g440(.A(KEYINPUT105), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n476), .A2(new_n517), .ZN(new_n643));
  INV_X1    g442(.A(new_n474), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n643), .A2(new_n644), .A3(new_n251), .A4(new_n637), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(G8gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT16), .B(G8gat), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n518), .A2(new_n644), .A3(new_n637), .A4(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(KEYINPUT42), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT42), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n642), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n652), .B1(new_n646), .B2(new_n649), .ZN(new_n655));
  INV_X1    g454(.A(new_n653), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n655), .A2(new_n656), .A3(KEYINPUT105), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n654), .A2(new_n657), .ZN(G1325gat));
  AND2_X1   g457(.A1(new_n518), .A2(new_n637), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT106), .ZN(new_n660));
  INV_X1    g459(.A(new_n514), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT36), .B1(new_n465), .B2(new_n466), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n516), .A2(KEYINPUT106), .A3(new_n514), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n659), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n467), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(G15gat), .ZN(new_n669));
  AOI22_X1  g468(.A1(new_n667), .A2(G15gat), .B1(new_n659), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT107), .ZN(G1326gat));
  NOR2_X1   g470(.A1(new_n638), .A2(new_n313), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT43), .B(G22gat), .Z(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(G1327gat));
  AOI21_X1  g473(.A(new_n620), .B1(new_n476), .B2(new_n517), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n601), .A2(new_n635), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n251), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n675), .A2(new_n219), .A3(new_n512), .A4(new_n678), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n426), .A2(new_n313), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n504), .A2(new_n313), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n683), .B1(new_n684), .B2(new_n492), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n661), .A2(new_n662), .ZN(new_n686));
  AOI22_X1  g485(.A1(new_n685), .A2(new_n686), .B1(new_n463), .B2(new_n475), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n682), .B1(new_n687), .B2(new_n620), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n675), .A2(KEYINPUT44), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n690), .A2(new_n512), .A3(new_n678), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n681), .B1(new_n691), .B2(new_n219), .ZN(G1328gat));
  NOR2_X1   g491(.A1(new_n474), .A2(G36gat), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n675), .A2(new_n678), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n675), .A2(new_n678), .A3(new_n697), .A4(new_n693), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n688), .A2(new_n689), .A3(new_n644), .A4(new_n678), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(G36gat), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(KEYINPUT110), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT110), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n699), .A2(new_n701), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(G1329gat));
  NOR2_X1   g505(.A1(new_n620), .A2(G43gat), .ZN(new_n707));
  AND4_X1   g506(.A1(new_n467), .A2(new_n518), .A3(new_n676), .A4(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT47), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n708), .B1(KEYINPUT111), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n686), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n688), .A2(new_n689), .A3(new_n711), .A4(new_n678), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n712), .A2(KEYINPUT47), .A3(G43gat), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n688), .A2(new_n689), .A3(new_n666), .A4(new_n678), .ZN(new_n715));
  AOI22_X1  g514(.A1(new_n715), .A2(G43gat), .B1(new_n708), .B2(KEYINPUT111), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n714), .B1(KEYINPUT47), .B2(new_n716), .ZN(G1330gat));
  NAND3_X1  g516(.A1(new_n675), .A2(new_n510), .A3(new_n678), .ZN(new_n718));
  INV_X1    g517(.A(G50gat), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT112), .ZN(new_n720));
  AOI22_X1  g519(.A1(new_n718), .A2(new_n719), .B1(new_n720), .B2(KEYINPUT48), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n313), .A2(new_n719), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n688), .A2(new_n689), .A3(new_n678), .A4(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  OR2_X1    g523(.A1(new_n720), .A2(KEYINPUT48), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1331gat));
  NOR2_X1   g525(.A1(new_n636), .A2(new_n251), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n643), .A2(new_n601), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n512), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n644), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n732));
  XOR2_X1   g531(.A(KEYINPUT49), .B(G64gat), .Z(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n731), .B2(new_n733), .ZN(G1333gat));
  NAND2_X1  g533(.A1(new_n728), .A2(new_n467), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n528), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n665), .A2(new_n528), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n728), .A2(KEYINPUT113), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT113), .B1(new_n728), .B2(new_n737), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n736), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT50), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT50), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n736), .B(new_n742), .C1(new_n738), .C2(new_n739), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(G1334gat));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n510), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g545(.A1(new_n251), .A2(new_n635), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n601), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT114), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n690), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G85gat), .B1(new_n750), .B2(new_n511), .ZN(new_n751));
  INV_X1    g550(.A(new_n620), .ZN(new_n752));
  AND4_X1   g551(.A1(KEYINPUT51), .A2(new_n643), .A3(new_n752), .A4(new_n747), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT51), .B1(new_n675), .B2(new_n747), .ZN(new_n754));
  OR2_X1    g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n755), .A2(new_n539), .A3(new_n512), .A4(new_n601), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n751), .A2(new_n756), .ZN(G1336gat));
  NAND4_X1  g556(.A1(new_n688), .A2(new_n689), .A3(new_n644), .A4(new_n749), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(G92gat), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n474), .A2(G92gat), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n601), .B(new_n760), .C1(new_n753), .C2(new_n754), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n759), .A2(new_n761), .A3(KEYINPUT115), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(KEYINPUT52), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n759), .A2(new_n761), .A3(KEYINPUT115), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(G1337gat));
  OAI21_X1  g565(.A(G99gat), .B1(new_n750), .B2(new_n665), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n668), .A2(new_n600), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n755), .A2(new_n553), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(G1338gat));
  NAND4_X1  g569(.A1(new_n688), .A2(new_n689), .A3(new_n510), .A4(new_n749), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G106gat), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n313), .A2(G106gat), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n601), .B(new_n773), .C1(new_n753), .C2(new_n754), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT53), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n772), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(G1339gat));
  NAND2_X1  g578(.A1(new_n727), .A2(new_n600), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n239), .A2(new_n240), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n231), .B1(new_n230), .B2(new_n232), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n246), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n250), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n597), .A2(new_n599), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT116), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n578), .A2(new_n584), .A3(new_n524), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n594), .A2(KEYINPUT54), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n522), .B1(new_n594), .B2(KEYINPUT54), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n788), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n595), .B1(new_n585), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n594), .A2(KEYINPUT54), .A3(new_n789), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n794), .A2(new_n795), .A3(KEYINPUT55), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n792), .A2(new_n251), .A3(new_n596), .A4(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n597), .A2(new_n798), .A3(new_n785), .A4(new_n599), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n787), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n620), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n796), .A2(new_n596), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n785), .A2(new_n618), .A3(new_n619), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT55), .B1(new_n794), .B2(new_n795), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n801), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n635), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n781), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(new_n511), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n467), .A2(new_n313), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(new_n644), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(G113gat), .B1(new_n814), .B2(new_n251), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n809), .A2(new_n510), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n644), .A2(new_n511), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n818), .A2(new_n668), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n251), .A2(G113gat), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n815), .B1(new_n819), .B2(new_n820), .ZN(G1340gat));
  NOR2_X1   g620(.A1(new_n813), .A2(new_n600), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n768), .A2(G120gat), .ZN(new_n823));
  OAI22_X1  g622(.A1(new_n822), .A2(G120gat), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(KEYINPUT117), .ZN(G1341gat));
  INV_X1    g624(.A(new_n819), .ZN(new_n826));
  OAI21_X1  g625(.A(G127gat), .B1(new_n826), .B2(new_n808), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n808), .A2(G127gat), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n827), .B1(new_n813), .B2(new_n828), .ZN(G1342gat));
  NAND2_X1  g628(.A1(new_n474), .A2(new_n752), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(KEYINPUT118), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n831), .A2(G134gat), .A3(new_n811), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n810), .ZN(new_n833));
  XOR2_X1   g632(.A(new_n833), .B(KEYINPUT56), .Z(new_n834));
  OAI21_X1  g633(.A(G134gat), .B1(new_n826), .B2(new_n620), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(G1343gat));
  AND2_X1   g635(.A1(new_n686), .A2(new_n817), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n838));
  OAI211_X1 g637(.A(KEYINPUT119), .B(new_n838), .C1(new_n809), .C2(new_n313), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n797), .A2(new_n786), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n805), .B1(new_n840), .B2(new_n620), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n780), .B1(new_n841), .B2(new_n635), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n313), .A2(new_n838), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n839), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n805), .B1(new_n800), .B2(new_n620), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n780), .B1(new_n846), .B2(new_n635), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n510), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT119), .B1(new_n848), .B2(new_n838), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n837), .B1(new_n845), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n266), .B1(new_n850), .B2(new_n252), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n313), .B1(new_n663), .B2(new_n664), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(new_n474), .A3(new_n810), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n252), .A2(G141gat), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(KEYINPUT121), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(new_n854), .B2(new_n856), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n851), .A2(new_n852), .A3(new_n858), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n850), .A2(KEYINPUT120), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n863), .B(new_n837), .C1(new_n845), .C2(new_n849), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n862), .A2(new_n251), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n857), .B1(new_n865), .B2(new_n266), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n861), .B1(new_n866), .B2(new_n852), .ZN(G1344gat));
  NAND2_X1  g666(.A1(new_n264), .A2(KEYINPUT59), .ZN(new_n868));
  INV_X1    g667(.A(new_n854), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n868), .B1(new_n869), .B2(new_n601), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n862), .A2(new_n864), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n600), .A2(KEYINPUT59), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n847), .A2(new_n843), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n842), .A2(new_n510), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n876), .B2(KEYINPUT57), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n601), .A3(new_n837), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n264), .B1(new_n878), .B2(KEYINPUT59), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n870), .B1(new_n874), .B2(new_n879), .ZN(G1345gat));
  AOI21_X1  g679(.A(G155gat), .B1(new_n869), .B2(new_n635), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n635), .A2(G155gat), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT122), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n881), .B1(new_n872), .B2(new_n883), .ZN(G1346gat));
  OAI21_X1  g683(.A(G162gat), .B1(new_n871), .B2(new_n620), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n831), .A2(G162gat), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n853), .A2(new_n810), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(G1347gat));
  NOR2_X1   g687(.A1(new_n512), .A2(new_n474), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n816), .A2(new_n467), .A3(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(G169gat), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n890), .A2(new_n891), .A3(new_n252), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n811), .A2(new_n474), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT123), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n809), .A2(new_n512), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n251), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n892), .B1(new_n898), .B2(new_n891), .ZN(G1348gat));
  INV_X1    g698(.A(G176gat), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n890), .A2(new_n900), .A3(new_n600), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n897), .A2(new_n601), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n902), .B2(new_n900), .ZN(G1349gat));
  NAND3_X1  g702(.A1(new_n897), .A2(new_n343), .A3(new_n635), .ZN(new_n904));
  OAI21_X1  g703(.A(G183gat), .B1(new_n890), .B2(new_n808), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g706(.A(G190gat), .B1(new_n890), .B2(new_n620), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT61), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n897), .A2(new_n322), .A3(new_n752), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(G1351gat));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n853), .A2(new_n644), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n912), .B1(new_n913), .B2(new_n896), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n853), .A2(KEYINPUT124), .A3(new_n644), .A4(new_n895), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n914), .A2(new_n251), .A3(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(G197gat), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n877), .A2(new_n665), .A3(new_n889), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n252), .A2(new_n917), .ZN(new_n919));
  AOI22_X1  g718(.A1(new_n916), .A2(new_n917), .B1(new_n918), .B2(new_n919), .ZN(G1352gat));
  NOR4_X1   g719(.A1(new_n913), .A2(G204gat), .A3(new_n896), .A4(new_n600), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n918), .A2(new_n601), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G204gat), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n921), .A2(new_n922), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n923), .A2(new_n925), .A3(new_n926), .ZN(G1353gat));
  NAND4_X1  g726(.A1(new_n877), .A2(new_n635), .A3(new_n665), .A4(new_n889), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT126), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(KEYINPUT63), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n928), .A2(G211gat), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n928), .B2(G211gat), .ZN(new_n932));
  OAI22_X1  g731(.A1(new_n931), .A2(new_n932), .B1(new_n929), .B2(KEYINPUT63), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n914), .A2(new_n255), .A3(new_n635), .A4(new_n915), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n934), .A2(KEYINPUT125), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n934), .A2(KEYINPUT125), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(G1354gat));
  AOI211_X1 g736(.A(new_n254), .B(new_n620), .C1(new_n918), .C2(KEYINPUT127), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n918), .A2(KEYINPUT127), .ZN(new_n939));
  INV_X1    g738(.A(G218gat), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n914), .A2(new_n752), .A3(new_n915), .ZN(new_n941));
  AOI22_X1  g740(.A1(new_n938), .A2(new_n939), .B1(new_n940), .B2(new_n941), .ZN(G1355gat));
endmodule


