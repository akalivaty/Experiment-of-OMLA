//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 0 0 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  OAI211_X1 g003(.A(KEYINPUT72), .B(new_n188), .C1(new_n189), .C2(KEYINPUT71), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT72), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT71), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G125), .ZN(new_n193));
  OAI21_X1  g007(.A(G140), .B1(new_n189), .B2(KEYINPUT72), .ZN(new_n194));
  OAI211_X1 g008(.A(KEYINPUT16), .B(new_n190), .C1(new_n193), .C2(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n189), .A2(G140), .ZN(new_n196));
  OR2_X1    g010(.A1(new_n196), .A2(KEYINPUT16), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n187), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n188), .A2(G125), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n189), .A2(G140), .ZN(new_n201));
  AND3_X1   g015(.A1(new_n200), .A2(new_n201), .A3(KEYINPUT74), .ZN(new_n202));
  AOI21_X1  g016(.A(KEYINPUT74), .B1(new_n200), .B2(new_n201), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n187), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT69), .ZN(new_n205));
  INV_X1    g019(.A(G119), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(G128), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(G128), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(KEYINPUT69), .A3(G119), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT24), .B(G110), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT73), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT23), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n215), .B1(new_n206), .B2(G128), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n209), .A2(KEYINPUT23), .A3(G119), .ZN(new_n217));
  INV_X1    g031(.A(G110), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n208), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n213), .A2(new_n214), .A3(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n214), .B1(new_n213), .B2(new_n219), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n199), .B(new_n204), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n210), .A2(new_n208), .ZN(new_n223));
  INV_X1    g037(.A(new_n212), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT70), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n223), .A2(new_n224), .A3(new_n225), .A4(new_n207), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT70), .B1(new_n211), .B2(new_n212), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n216), .A2(new_n217), .A3(new_n208), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G110), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n195), .A2(new_n187), .A3(new_n197), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n228), .B(new_n230), .C1(new_n232), .C2(new_n198), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n222), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G953), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(G221), .A3(G234), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n236), .B(KEYINPUT75), .ZN(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT22), .B(G137), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n234), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G902), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n222), .A2(new_n233), .A3(new_n239), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT76), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT25), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G217), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n249), .B1(G234), .B2(new_n242), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n244), .A2(new_n245), .A3(KEYINPUT25), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n248), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n250), .A2(G902), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n253), .B(KEYINPUT78), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT77), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n241), .A2(new_n256), .A3(new_n243), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n256), .B1(new_n241), .B2(new_n243), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n255), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n252), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n206), .A2(G116), .ZN(new_n261));
  INV_X1    g075(.A(G116), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G119), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT2), .B(G113), .ZN(new_n265));
  OR2_X1    g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n265), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n269));
  INV_X1    g083(.A(G134), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n269), .B1(new_n270), .B2(G137), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(G137), .ZN(new_n272));
  INV_X1    g086(.A(G137), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(KEYINPUT65), .A3(G134), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n271), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G131), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT11), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n277), .B1(new_n270), .B2(G137), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n273), .A2(KEYINPUT11), .A3(G134), .ZN(new_n279));
  INV_X1    g093(.A(G131), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n278), .A2(new_n279), .A3(new_n280), .A4(new_n272), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n276), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n209), .A2(KEYINPUT1), .ZN(new_n283));
  INV_X1    g097(.A(G143), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G146), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n187), .A2(G143), .ZN(new_n286));
  OAI22_X1  g100(.A1(new_n283), .A2(new_n285), .B1(new_n286), .B2(G128), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(G143), .B(G146), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT66), .B1(new_n289), .B2(new_n283), .ZN(new_n290));
  AND4_X1   g104(.A1(KEYINPUT66), .A2(new_n283), .A3(new_n286), .A4(new_n285), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n288), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n278), .A2(new_n279), .A3(new_n272), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G131), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n281), .ZN(new_n295));
  AND2_X1   g109(.A1(KEYINPUT0), .A2(G128), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n286), .A2(new_n285), .A3(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT0), .B(G128), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n297), .B1(new_n289), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n282), .A2(new_n292), .B1(new_n295), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT30), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n283), .A2(new_n286), .A3(new_n285), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT66), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n289), .A2(KEYINPUT66), .A3(new_n283), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n287), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n276), .A2(new_n281), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n295), .A2(new_n300), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT64), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n299), .B1(new_n281), .B2(new_n294), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT64), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n309), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n268), .B(new_n302), .C1(new_n315), .C2(KEYINPUT30), .ZN(new_n316));
  NOR2_X1   g130(.A1(G237), .A2(G953), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G210), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n318), .B(KEYINPUT27), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT26), .B(G101), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n319), .B(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT67), .ZN(new_n322));
  INV_X1    g136(.A(new_n268), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n322), .B1(new_n301), .B2(new_n323), .ZN(new_n324));
  NOR4_X1   g138(.A1(new_n309), .A2(new_n313), .A3(KEYINPUT67), .A4(new_n268), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n316), .A2(new_n321), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT31), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT31), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n316), .A2(new_n326), .A3(new_n329), .A4(new_n321), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT28), .B1(new_n301), .B2(new_n323), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n310), .B(new_n323), .C1(new_n307), .C2(new_n308), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT67), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n301), .A2(new_n322), .A3(new_n323), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n333), .B(new_n334), .C1(new_n315), .C2(new_n323), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n331), .B1(new_n335), .B2(KEYINPUT28), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n328), .B(new_n330), .C1(new_n321), .C2(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(G472), .A2(G902), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n337), .A2(KEYINPUT32), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT32), .B1(new_n337), .B2(new_n338), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n333), .B(new_n334), .C1(new_n323), .C2(new_n301), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n331), .B1(new_n342), .B2(KEYINPUT28), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n321), .A2(KEYINPUT29), .ZN(new_n344));
  AOI21_X1  g158(.A(G902), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n336), .A2(KEYINPUT68), .A3(new_n321), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n316), .A2(new_n326), .ZN(new_n347));
  INV_X1    g161(.A(new_n321), .ZN(new_n348));
  AOI21_X1  g162(.A(KEYINPUT29), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT68), .B1(new_n336), .B2(new_n321), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n345), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G472), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n260), .B1(new_n341), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT9), .B(G234), .ZN(new_n355));
  OAI21_X1  g169(.A(G221), .B1(new_n355), .B2(G902), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G104), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT3), .B1(new_n358), .B2(G107), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT3), .ZN(new_n360));
  INV_X1    g174(.A(G107), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n361), .A3(G104), .ZN(new_n362));
  INV_X1    g176(.A(G101), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n358), .A2(G107), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n359), .A2(new_n362), .A3(new_n363), .A4(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n358), .A2(G107), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n361), .A2(G104), .ZN(new_n367));
  OAI21_X1  g181(.A(G101), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT80), .B1(new_n292), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n292), .A2(new_n370), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT80), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n307), .A2(new_n373), .A3(new_n369), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n371), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(KEYINPUT12), .A3(new_n295), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(KEYINPUT12), .B1(new_n375), .B2(new_n295), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT81), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n374), .A2(new_n372), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n373), .B1(new_n307), .B2(new_n369), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n295), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT12), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT81), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(new_n376), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n295), .B(KEYINPUT79), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT10), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n372), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n359), .A2(new_n362), .A3(new_n364), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G101), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(KEYINPUT4), .A3(new_n365), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n390), .A2(new_n393), .A3(G101), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n300), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n292), .A2(KEYINPUT10), .A3(new_n370), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n387), .A2(new_n389), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(G110), .B(G140), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n235), .A2(G227), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n398), .B(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n379), .A2(new_n386), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n389), .A2(new_n395), .A3(new_n396), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n295), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n401), .B1(new_n406), .B2(new_n397), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G469), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n410), .A3(new_n242), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n397), .B1(new_n377), .B2(new_n378), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n412), .A2(new_n400), .B1(new_n406), .B2(new_n403), .ZN(new_n413));
  OAI21_X1  g227(.A(G469), .B1(new_n413), .B2(G902), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n357), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(G113), .B(G122), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT91), .B(G104), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n416), .B(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT89), .ZN(new_n419));
  NOR3_X1   g233(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT19), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT19), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n188), .B1(new_n191), .B2(G125), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT72), .B1(new_n189), .B2(KEYINPUT71), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n421), .B1(new_n424), .B2(new_n190), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n419), .B(new_n187), .C1(new_n420), .C2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n199), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n190), .B1(new_n193), .B2(new_n194), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(KEYINPUT19), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT74), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n188), .A2(G125), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n430), .B1(new_n196), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n200), .A2(new_n201), .A3(KEYINPUT74), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n421), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(G146), .B1(new_n429), .B2(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(new_n419), .ZN(new_n436));
  OAI21_X1  g250(.A(KEYINPUT90), .B1(new_n427), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(G237), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n235), .A3(G214), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT86), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n440), .A3(new_n284), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n317), .B(G214), .C1(KEYINPUT86), .C2(G143), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G131), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n441), .A2(new_n280), .A3(new_n442), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n198), .B1(new_n435), .B2(new_n419), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n187), .B1(new_n420), .B2(new_n425), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT89), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT90), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n447), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n437), .A2(new_n446), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT18), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n453), .A2(new_n280), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT88), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT88), .B1(new_n453), .B2(new_n280), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n441), .A2(new_n456), .A3(new_n442), .A4(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n424), .A2(G146), .A3(new_n190), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n204), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT87), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n443), .A2(new_n461), .A3(new_n454), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n461), .B1(new_n443), .B2(new_n454), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n458), .B(new_n460), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n418), .B1(new_n452), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT17), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n444), .A2(new_n466), .A3(new_n445), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n443), .A2(KEYINPUT17), .A3(G131), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n467), .A2(new_n199), .A3(new_n231), .A4(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(new_n464), .A3(new_n418), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT92), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(G475), .A2(G902), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(KEYINPUT20), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT20), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n476), .B(new_n473), .C1(new_n465), .C2(new_n471), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(G214), .B1(G237), .B2(G902), .ZN(new_n479));
  XOR2_X1   g293(.A(new_n479), .B(KEYINPUT82), .Z(new_n480));
  NAND2_X1  g294(.A1(G234), .A2(G237), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(G952), .A3(new_n235), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n481), .A2(G902), .A3(G953), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT21), .B(G898), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(G210), .B1(G237), .B2(G902), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n300), .A2(G125), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n490), .B1(G125), .B2(new_n307), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n235), .A2(G224), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(KEYINPUT85), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n491), .B(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n392), .A2(new_n268), .A3(new_n394), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT5), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT83), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT83), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT5), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n497), .A2(new_n499), .A3(G116), .A4(new_n206), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n497), .A2(new_n499), .ZN(new_n501));
  OAI211_X1 g315(.A(G113), .B(new_n500), .C1(new_n501), .C2(new_n264), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n370), .A2(new_n266), .A3(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(G110), .B(G122), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n495), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT6), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n495), .A2(new_n503), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n504), .A2(KEYINPUT84), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n507), .A2(KEYINPUT6), .A3(new_n508), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n494), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n504), .B(KEYINPUT8), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n370), .B1(new_n266), .B2(new_n502), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n261), .A2(new_n263), .A3(KEYINPUT5), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n500), .A2(G113), .A3(new_n515), .ZN(new_n516));
  AND4_X1   g330(.A1(new_n266), .A2(new_n516), .A3(new_n365), .A4(new_n368), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n513), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n492), .A2(KEYINPUT7), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n491), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n490), .B(new_n519), .C1(G125), .C2(new_n307), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n518), .A2(new_n521), .A3(new_n505), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n242), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n489), .B1(new_n512), .B2(new_n524), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n523), .A2(new_n242), .ZN(new_n526));
  INV_X1    g340(.A(new_n493), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n491), .B(new_n527), .ZN(new_n528));
  AOI22_X1  g342(.A1(new_n505), .A2(KEYINPUT6), .B1(new_n507), .B2(new_n508), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n507), .A2(KEYINPUT6), .A3(new_n508), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n526), .A2(new_n531), .A3(new_n488), .ZN(new_n532));
  AOI211_X1 g346(.A(new_n480), .B(new_n487), .C1(new_n525), .C2(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(G128), .B(G143), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT13), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n209), .A2(KEYINPUT13), .A3(G143), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n536), .A2(new_n270), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n534), .A2(new_n270), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n535), .A2(new_n537), .B1(new_n538), .B2(KEYINPUT94), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n539), .B1(KEYINPUT94), .B2(new_n538), .ZN(new_n540));
  AND2_X1   g354(.A1(KEYINPUT93), .A2(G122), .ZN(new_n541));
  NOR2_X1   g355(.A1(KEYINPUT93), .A2(G122), .ZN(new_n542));
  OAI21_X1  g356(.A(G116), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n262), .A2(G122), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(new_n361), .ZN(new_n546));
  OR2_X1    g360(.A1(new_n540), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n544), .B(KEYINPUT14), .ZN(new_n548));
  INV_X1    g362(.A(new_n543), .ZN(new_n549));
  OAI21_X1  g363(.A(G107), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n534), .B(new_n270), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n550), .B(new_n551), .C1(G107), .C2(new_n545), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n355), .A2(new_n249), .A3(G953), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n547), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n552), .B1(new_n540), .B2(new_n546), .ZN(new_n555));
  INV_X1    g369(.A(new_n553), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(G478), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(KEYINPUT15), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n558), .A2(new_n242), .A3(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n561), .B1(new_n558), .B2(new_n242), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(G475), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT92), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n470), .B(new_n567), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n469), .A2(new_n464), .ZN(new_n569));
  OR2_X1    g383(.A1(new_n569), .A2(new_n418), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n566), .B1(new_n571), .B2(new_n242), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n478), .A2(new_n533), .A3(new_n565), .A4(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n354), .A2(new_n415), .A3(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(G101), .ZN(G3));
  AOI21_X1  g391(.A(new_n572), .B1(new_n475), .B2(new_n477), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n558), .A2(new_n559), .A3(new_n242), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n559), .A2(new_n242), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  XOR2_X1   g396(.A(new_n558), .B(KEYINPUT33), .Z(new_n583));
  AOI21_X1  g397(.A(new_n582), .B1(new_n583), .B2(G478), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n479), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n488), .B1(new_n526), .B2(new_n531), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n586), .B1(new_n587), .B2(KEYINPUT96), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT96), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n525), .A2(new_n589), .A3(new_n532), .ZN(new_n590));
  INV_X1    g404(.A(new_n487), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n578), .A2(new_n585), .A3(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n250), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n594), .B1(new_n246), .B2(new_n247), .ZN(new_n595));
  OR2_X1    g409(.A1(new_n257), .A2(new_n258), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n251), .A2(new_n595), .B1(new_n596), .B2(new_n255), .ZN(new_n597));
  AOI211_X1 g411(.A(G469), .B(G902), .C1(new_n404), .C2(new_n408), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n403), .A2(new_n406), .ZN(new_n599));
  INV_X1    g413(.A(new_n397), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n384), .B2(new_n376), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n599), .B1(new_n601), .B2(new_n401), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n410), .B1(new_n602), .B2(new_n242), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n597), .B(new_n356), .C1(new_n598), .C2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n337), .A2(new_n242), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT95), .ZN(new_n607));
  INV_X1    g421(.A(G472), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n337), .B(new_n242), .C1(new_n607), .C2(new_n608), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n593), .A2(new_n605), .A3(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT34), .B(G104), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G6));
  INV_X1    g429(.A(new_n464), .ZN(new_n616));
  INV_X1    g430(.A(new_n446), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n447), .A2(new_n449), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n617), .B1(new_n618), .B2(KEYINPUT90), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n616), .B1(new_n619), .B2(new_n451), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n568), .B1(new_n620), .B2(new_n418), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n476), .B1(new_n621), .B2(new_n473), .ZN(new_n622));
  INV_X1    g436(.A(new_n477), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n573), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n624), .A2(new_n565), .A3(new_n592), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n625), .A2(new_n605), .A3(new_n612), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT35), .B(G107), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G9));
  NOR2_X1   g442(.A1(new_n240), .A2(KEYINPUT36), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n234), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n255), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n252), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n610), .A2(new_n611), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n356), .B1(new_n598), .B2(new_n603), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n633), .A2(new_n574), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT37), .B(G110), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(KEYINPUT97), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n635), .B(new_n637), .ZN(G12));
  AOI21_X1  g452(.A(new_n634), .B1(new_n341), .B2(new_n353), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n640));
  INV_X1    g454(.A(new_n565), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n482), .B1(new_n484), .B2(G900), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n578), .A2(new_n640), .A3(new_n641), .A4(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n578), .A2(new_n641), .A3(new_n642), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(KEYINPUT98), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n588), .A2(new_n590), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n646), .A2(new_n632), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n639), .A2(new_n643), .A3(new_n645), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G128), .ZN(G30));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n337), .A2(new_n338), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT32), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n337), .A2(KEYINPUT32), .A3(new_n338), .ZN(new_n654));
  INV_X1    g468(.A(new_n347), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n348), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n242), .B1(new_n342), .B2(new_n321), .ZN(new_n657));
  OAI21_X1  g471(.A(G472), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n653), .A2(new_n654), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(KEYINPUT99), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT99), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n653), .A2(new_n661), .A3(new_n654), .A4(new_n658), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT100), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n525), .A2(new_n532), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n665), .B(KEYINPUT38), .Z(new_n666));
  NOR2_X1   g480(.A1(new_n578), .A2(new_n565), .ZN(new_n667));
  INV_X1    g481(.A(new_n632), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n666), .A2(new_n479), .A3(new_n667), .A4(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n642), .B(KEYINPUT39), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g486(.A(KEYINPUT101), .B1(new_n634), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT101), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n415), .A2(new_n674), .A3(new_n671), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n673), .A2(KEYINPUT40), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(KEYINPUT40), .B1(new_n673), .B2(new_n675), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n670), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n650), .B1(new_n664), .B2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT100), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n663), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n673), .A2(new_n675), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT40), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n673), .A2(KEYINPUT40), .A3(new_n675), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n669), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n681), .A2(new_n686), .A3(KEYINPUT102), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n679), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(new_n284), .ZN(G45));
  NAND3_X1  g503(.A1(new_n624), .A2(new_n584), .A3(new_n642), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n624), .A2(KEYINPUT103), .A3(new_n584), .A4(new_n642), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n639), .A2(new_n692), .A3(new_n647), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  NAND2_X1  g509(.A1(new_n384), .A2(new_n376), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n402), .B1(new_n696), .B2(KEYINPUT81), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n407), .B1(new_n697), .B2(new_n386), .ZN(new_n698));
  OAI21_X1  g512(.A(G469), .B1(new_n698), .B2(G902), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n699), .A2(new_n356), .A3(new_n411), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n354), .A2(new_n593), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT41), .B(G113), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G15));
  NAND3_X1  g517(.A1(new_n354), .A2(new_n625), .A3(new_n700), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  NAND3_X1  g519(.A1(new_n353), .A2(new_n653), .A3(new_n654), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n624), .A2(new_n641), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n668), .A2(new_n592), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n706), .A2(new_n707), .A3(new_n700), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G119), .ZN(G21));
  NAND2_X1  g524(.A1(new_n700), .A2(new_n591), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n624), .A2(new_n646), .A3(new_n712), .A4(new_n641), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n624), .A2(new_n646), .A3(new_n641), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(KEYINPUT108), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n711), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n343), .A2(KEYINPUT104), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n348), .B1(new_n343), .B2(KEYINPUT104), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n328), .B(new_n330), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n338), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT105), .B(G472), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n606), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n252), .A2(KEYINPUT106), .A3(new_n259), .ZN(new_n724));
  AOI21_X1  g538(.A(KEYINPUT106), .B1(new_n252), .B2(new_n259), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g540(.A(KEYINPUT107), .B1(new_n723), .B2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n725), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n597), .A2(KEYINPUT106), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n731));
  AOI22_X1  g545(.A1(new_n338), .A2(new_n719), .B1(new_n606), .B2(new_n721), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n727), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n716), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  NAND3_X1  g550(.A1(new_n720), .A2(new_n722), .A3(new_n632), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n646), .A2(new_n699), .A3(new_n356), .A4(new_n411), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n692), .A2(new_n738), .A3(new_n740), .A4(new_n693), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G125), .ZN(G27));
  NAND3_X1  g556(.A1(new_n525), .A2(new_n532), .A3(new_n479), .ZN(new_n743));
  NAND2_X1  g557(.A1(G469), .A2(G902), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT109), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n746), .B1(new_n413), .B2(G469), .ZN(new_n747));
  AOI211_X1 g561(.A(new_n357), .B(new_n743), .C1(new_n411), .C2(new_n747), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n748), .A2(KEYINPUT42), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n726), .B1(new_n353), .B2(new_n341), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n692), .A2(new_n693), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT42), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n706), .A2(new_n597), .A3(new_n748), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n755), .B(new_n756), .C1(new_n752), .C2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n354), .A2(new_n692), .A3(new_n693), .A4(new_n748), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n755), .B1(new_n760), .B2(new_n756), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n754), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G131), .ZN(G33));
  NAND2_X1  g577(.A1(new_n645), .A2(new_n643), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n757), .ZN(new_n765));
  XNOR2_X1  g579(.A(KEYINPUT111), .B(G134), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(G36));
  NOR2_X1   g581(.A1(new_n612), .A2(new_n668), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT43), .B1(new_n624), .B2(new_n585), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n624), .A2(new_n585), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT43), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n768), .A2(new_n769), .A3(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT44), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n743), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n768), .A2(KEYINPUT44), .A3(new_n769), .A4(new_n772), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT46), .ZN(new_n780));
  OAI21_X1  g594(.A(G469), .B1(new_n413), .B2(KEYINPUT45), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT45), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n602), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n780), .B1(new_n784), .B2(new_n746), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n411), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n784), .A2(new_n780), .A3(new_n746), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n356), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n672), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n773), .A2(new_n774), .ZN(new_n790));
  INV_X1    g604(.A(new_n743), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n790), .A2(KEYINPUT112), .A3(new_n791), .A4(new_n776), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n779), .A2(new_n789), .A3(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G137), .ZN(G39));
  INV_X1    g608(.A(KEYINPUT47), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n788), .A2(new_n795), .ZN(new_n796));
  OAI211_X1 g610(.A(KEYINPUT47), .B(new_n356), .C1(new_n786), .C2(new_n787), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR4_X1   g612(.A1(new_n752), .A2(new_n706), .A3(new_n597), .A4(new_n743), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G140), .ZN(G42));
  NOR3_X1   g615(.A1(new_n666), .A2(new_n357), .A3(new_n480), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n802), .A2(new_n730), .A3(new_n770), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n699), .A2(new_n411), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT49), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n664), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT51), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n798), .B1(new_n357), .B2(new_n804), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n772), .A2(new_n769), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n809), .A2(new_n734), .A3(new_n483), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n791), .ZN(new_n811));
  INV_X1    g625(.A(new_n700), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n812), .A2(new_n666), .A3(new_n479), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n810), .A2(KEYINPUT50), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT50), .B1(new_n810), .B2(new_n813), .ZN(new_n815));
  OAI22_X1  g629(.A1(new_n808), .A2(new_n811), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n812), .A2(new_n482), .A3(new_n743), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n597), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n681), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n578), .A3(new_n585), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n809), .A2(new_n817), .A3(new_n738), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n807), .B1(new_n816), .B2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(G952), .ZN(new_n824));
  AOI211_X1 g638(.A(new_n824), .B(G953), .C1(new_n810), .C2(new_n740), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n809), .A2(new_n817), .A3(new_n750), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT48), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n578), .A2(new_n585), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n828), .B1(new_n829), .B2(new_n819), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n823), .A2(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n816), .A2(new_n822), .A3(new_n807), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n692), .A2(new_n693), .A3(new_n732), .A4(new_n748), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n835), .B1(new_n563), .B2(new_n564), .ZN(new_n836));
  INV_X1    g650(.A(new_n564), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(KEYINPUT113), .A3(new_n562), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  AND4_X1   g654(.A1(new_n578), .A2(new_n840), .A3(new_n642), .A4(new_n791), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n639), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n834), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n765), .B1(new_n843), .B2(new_n632), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n648), .A2(new_n694), .A3(new_n741), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n715), .A2(new_n713), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n668), .A2(new_n356), .A3(new_n642), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n847), .B1(new_n411), .B2(new_n747), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n846), .A2(new_n663), .A3(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT52), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n844), .B1(new_n845), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n756), .B1(new_n752), .B2(new_n757), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT110), .ZN(new_n854));
  AOI22_X1  g668(.A1(new_n854), .A2(new_n758), .B1(new_n753), .B2(new_n751), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n846), .A2(new_n663), .A3(new_n848), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT52), .B1(new_n845), .B2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n415), .A2(new_n597), .A3(new_n610), .A4(new_n611), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n829), .A2(new_n533), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n576), .B(new_n709), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n701), .A2(new_n704), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n578), .A2(new_n533), .A3(new_n839), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT114), .B1(new_n865), .B2(new_n635), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n575), .A2(new_n612), .A3(new_n415), .A4(new_n632), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n624), .A2(new_n840), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n605), .A2(new_n612), .A3(new_n533), .A4(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT114), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n867), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n735), .A2(new_n866), .A3(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n858), .A2(new_n863), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n856), .A2(new_n873), .A3(KEYINPUT53), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT53), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n639), .A2(new_n647), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n645), .A2(new_n643), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n876), .B1(new_n753), .B2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n878), .A2(new_n850), .A3(new_n741), .A4(new_n849), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n762), .A2(new_n879), .A3(new_n844), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n858), .A2(new_n872), .A3(new_n863), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n875), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n874), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT115), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n883), .B1(new_n874), .B2(new_n882), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT53), .B1(new_n856), .B2(new_n873), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n880), .A2(new_n881), .A3(new_n875), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n890), .A2(KEYINPUT115), .A3(new_n883), .ZN(new_n891));
  OAI211_X1 g705(.A(KEYINPUT116), .B(new_n833), .C1(new_n887), .C2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n824), .A2(new_n235), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n885), .A2(new_n886), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n874), .A2(new_n882), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(KEYINPUT54), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(KEYINPUT115), .A3(new_n884), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT116), .B1(new_n899), .B2(new_n833), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n806), .B1(new_n894), .B2(new_n900), .ZN(G75));
  NAND2_X1  g715(.A1(new_n896), .A2(G902), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(G210), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n510), .A2(new_n511), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT117), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT55), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(new_n494), .ZN(new_n908));
  NOR2_X1   g722(.A1(KEYINPUT118), .A2(KEYINPUT56), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n904), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n908), .B1(new_n904), .B2(new_n909), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n235), .A2(G952), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(G51));
  INV_X1    g727(.A(KEYINPUT119), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n897), .A2(new_n914), .A3(new_n884), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n890), .A2(KEYINPUT119), .A3(new_n883), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n745), .B(KEYINPUT57), .Z(new_n917));
  NAND3_X1  g731(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n409), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n903), .A2(new_n784), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n912), .B1(new_n919), .B2(new_n920), .ZN(G54));
  NAND3_X1  g735(.A1(new_n903), .A2(KEYINPUT58), .A3(G475), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n922), .A2(new_n472), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n922), .A2(new_n472), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n923), .A2(new_n924), .A3(new_n912), .ZN(G60));
  XNOR2_X1  g739(.A(new_n580), .B(KEYINPUT59), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n583), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n915), .A2(new_n916), .A3(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n912), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OR2_X1    g744(.A1(new_n899), .A2(new_n926), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n930), .B1(new_n931), .B2(new_n583), .ZN(G63));
  XNOR2_X1  g746(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n249), .A2(new_n242), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n936), .B1(new_n874), .B2(new_n882), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n937), .A2(new_n630), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n929), .B1(new_n937), .B2(new_n596), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT121), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n941));
  OAI22_X1  g755(.A1(new_n938), .A2(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(G66));
  INV_X1    g758(.A(G224), .ZN(new_n945));
  OAI21_X1  g759(.A(G953), .B1(new_n486), .B2(new_n945), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n872), .A2(new_n863), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(G953), .ZN(new_n948));
  INV_X1    g762(.A(new_n906), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(G898), .B2(new_n235), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n948), .B(new_n950), .ZN(G69));
  OAI21_X1  g765(.A(new_n302), .B1(new_n315), .B2(KEYINPUT30), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n429), .A2(new_n434), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n954), .B1(G900), .B2(G953), .ZN(new_n955));
  INV_X1    g769(.A(new_n765), .ZN(new_n956));
  INV_X1    g770(.A(new_n845), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n789), .A2(new_n846), .A3(new_n750), .ZN(new_n958));
  AND4_X1   g772(.A1(new_n956), .A2(new_n800), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n959), .A2(new_n762), .A3(new_n793), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n955), .B1(new_n960), .B2(G953), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n235), .B1(G227), .B2(G900), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n961), .B1(KEYINPUT124), .B2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT123), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n679), .A2(new_n687), .A3(new_n957), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n679), .A2(new_n687), .A3(KEYINPUT62), .A4(new_n957), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n354), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n791), .B1(new_n829), .B2(new_n868), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n971), .A2(new_n682), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(new_n798), .B2(new_n799), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n792), .A2(new_n789), .ZN(new_n975));
  AOI21_X1  g789(.A(KEYINPUT112), .B1(new_n775), .B2(new_n776), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n965), .B1(new_n970), .B2(new_n978), .ZN(new_n979));
  AOI211_X1 g793(.A(KEYINPUT123), .B(new_n977), .C1(new_n968), .C2(new_n969), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n235), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n954), .B(KEYINPUT122), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n964), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT124), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n962), .A2(new_n984), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n983), .B(new_n985), .ZN(G72));
  NAND2_X1  g800(.A1(G472), .A2(G902), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT63), .Z(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n347), .A2(new_n321), .ZN(new_n990));
  OR4_X1    g804(.A1(new_n656), .A2(new_n890), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(KEYINPUT126), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n959), .A2(new_n762), .A3(new_n793), .A4(new_n947), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n993), .B1(new_n994), .B2(new_n988), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n995), .A2(new_n912), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n996), .A2(KEYINPUT127), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT127), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n995), .A2(new_n998), .A3(new_n912), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n991), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT125), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n979), .A2(new_n980), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n989), .B1(new_n1002), .B2(new_n947), .ZN(new_n1003));
  INV_X1    g817(.A(new_n656), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1001), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n872), .A2(new_n863), .ZN(new_n1006));
  NOR3_X1   g820(.A1(new_n979), .A2(new_n980), .A3(new_n1006), .ZN(new_n1007));
  OAI211_X1 g821(.A(KEYINPUT125), .B(new_n656), .C1(new_n1007), .C2(new_n989), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1000), .B1(new_n1005), .B2(new_n1008), .ZN(G57));
endmodule


