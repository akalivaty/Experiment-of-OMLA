//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 1 1 0 0 0 1 1 1 0 1 0 1 0 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n557,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n579, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n623,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n452), .A2(new_n457), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT67), .Z(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G137), .ZN(new_n466));
  NAND2_X1  g041(.A1(G101), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n462), .A2(new_n464), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(KEYINPUT68), .B1(new_n472), .B2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n472), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n468), .B1(new_n474), .B2(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n465), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  INV_X1    g054(.A(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n465), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n480), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n479), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NAND3_X1  g062(.A1(new_n462), .A2(new_n464), .A3(G126), .ZN(new_n488));
  NAND2_X1  g063(.A1(G114), .A2(G2104), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n480), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  OAI22_X1  g067(.A1(new_n490), .A2(new_n491), .B1(new_n481), .B2(new_n492), .ZN(new_n493));
  NOR3_X1   g068(.A1(new_n470), .A2(new_n491), .A3(new_n492), .ZN(new_n494));
  AND2_X1   g069(.A1(G102), .A2(G2104), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n480), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AND3_X1   g071(.A1(new_n493), .A2(KEYINPUT69), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(KEYINPUT69), .B1(new_n493), .B2(new_n496), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(KEYINPUT70), .A3(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n506), .B1(new_n504), .B2(KEYINPUT5), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n502), .A2(KEYINPUT71), .A3(G543), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n503), .A2(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G50), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n509), .A2(new_n513), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n512), .A2(new_n519), .ZN(G166));
  NAND3_X1  g095(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n515), .A2(G51), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n509), .A2(G89), .A3(new_n513), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n523), .A2(KEYINPUT72), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g101(.A(KEYINPUT72), .B1(new_n523), .B2(new_n525), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n521), .B(new_n522), .C1(new_n526), .C2(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  NAND2_X1  g104(.A1(G77), .A2(G543), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n503), .A2(new_n505), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n507), .A2(new_n508), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G64), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n530), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G651), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n531), .A2(new_n532), .A3(G90), .A4(new_n513), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT73), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n513), .A2(G52), .A3(G543), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n538), .B1(new_n537), .B2(new_n539), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n536), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(G171));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  INV_X1    g119(.A(G68), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n533), .A2(new_n544), .B1(new_n545), .B2(new_n504), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(KEYINPUT74), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT74), .ZN(new_n548));
  OAI221_X1 g123(.A(new_n548), .B1(new_n545), .B2(new_n504), .C1(new_n533), .C2(new_n544), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n547), .A2(G651), .A3(new_n549), .ZN(new_n550));
  AND3_X1   g125(.A1(new_n531), .A2(new_n532), .A3(new_n513), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n551), .A2(G81), .B1(G43), .B2(new_n515), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(new_n557));
  XOR2_X1   g132(.A(new_n557), .B(KEYINPUT75), .Z(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(G188));
  XNOR2_X1  g136(.A(KEYINPUT76), .B(KEYINPUT9), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n513), .A2(new_n562), .A3(G53), .A4(G543), .ZN(new_n563));
  AND2_X1   g138(.A1(KEYINPUT6), .A2(G651), .ZN(new_n564));
  NOR2_X1   g139(.A1(KEYINPUT6), .A2(G651), .ZN(new_n565));
  OAI211_X1 g140(.A(G53), .B(G543), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  OR2_X1    g141(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n551), .A2(G91), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n531), .A2(new_n532), .A3(G65), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT77), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(KEYINPUT78), .B1(new_n574), .B2(G651), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n576));
  AOI211_X1 g151(.A(new_n576), .B(new_n511), .C1(new_n571), .C2(new_n573), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n569), .B(new_n570), .C1(new_n575), .C2(new_n577), .ZN(G299));
  INV_X1    g153(.A(KEYINPUT79), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n542), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n536), .B(KEYINPUT79), .C1(new_n540), .C2(new_n541), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(G301));
  INV_X1    g157(.A(G166), .ZN(G303));
  OAI21_X1  g158(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n584));
  INV_X1    g159(.A(G49), .ZN(new_n585));
  INV_X1    g160(.A(G87), .ZN(new_n586));
  OAI221_X1 g161(.A(new_n584), .B1(new_n585), .B2(new_n514), .C1(new_n586), .C2(new_n517), .ZN(G288));
  AND4_X1   g162(.A1(G86), .A2(new_n531), .A3(new_n532), .A4(new_n513), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n533), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n588), .B1(new_n591), .B2(G651), .ZN(new_n592));
  OAI211_X1 g167(.A(G48), .B(G543), .C1(new_n564), .C2(new_n565), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT80), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n592), .A2(new_n595), .ZN(G305));
  XOR2_X1   g171(.A(KEYINPUT81), .B(G85), .Z(new_n597));
  AOI22_X1  g172(.A1(new_n551), .A2(new_n597), .B1(G47), .B2(new_n515), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n511), .B2(new_n599), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n600), .A2(KEYINPUT82), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(KEYINPUT82), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(G290));
  NAND4_X1  g178(.A1(new_n531), .A2(new_n532), .A3(G92), .A4(new_n513), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(KEYINPUT83), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT83), .ZN(new_n606));
  NAND4_X1  g181(.A1(new_n509), .A2(new_n606), .A3(G92), .A4(new_n513), .ZN(new_n607));
  AOI21_X1  g182(.A(KEYINPUT10), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n515), .A2(G54), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n509), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(new_n511), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n605), .A2(new_n607), .A3(KEYINPUT10), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n609), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(G301), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(new_n616), .ZN(G321));
  XOR2_X1   g194(.A(G321), .B(KEYINPUT84), .Z(G284));
  NAND2_X1  g195(.A1(G286), .A2(G868), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT85), .Z(new_n622));
  INV_X1    g197(.A(G299), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(G868), .B2(new_n623), .ZN(G297));
  OAI21_X1  g199(.A(new_n622), .B1(G868), .B2(new_n623), .ZN(G280));
  INV_X1    g200(.A(new_n614), .ZN(new_n626));
  NOR3_X1   g201(.A1(new_n626), .A2(new_n608), .A3(new_n612), .ZN(new_n627));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G860), .ZN(G148));
  NAND2_X1  g204(.A1(new_n553), .A2(new_n616), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n615), .A2(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(new_n616), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g208(.A1(new_n480), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT12), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2100), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n478), .A2(G123), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n482), .A2(G135), .ZN(new_n639));
  NOR2_X1   g214(.A1(G99), .A2(G2105), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(new_n480), .B2(G111), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n638), .B(new_n639), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(KEYINPUT86), .B(G2096), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n637), .A2(new_n644), .ZN(G156));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2435), .ZN(new_n647));
  XOR2_X1   g222(.A(G2427), .B(G2438), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(KEYINPUT14), .ZN(new_n650));
  XOR2_X1   g225(.A(G2451), .B(G2454), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G1341), .B(G1348), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2443), .B(G2446), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(G14), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT87), .Z(G401));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  XOR2_X1   g235(.A(G2067), .B(G2678), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n660), .B1(new_n664), .B2(KEYINPUT18), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2096), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2100), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n662), .A2(new_n663), .ZN(new_n669));
  AOI21_X1  g244(.A(KEYINPUT18), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n667), .B(new_n670), .Z(G227));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n672), .A2(new_n673), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n678), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n675), .A2(new_n677), .A3(new_n679), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n682), .B(new_n683), .C1(new_n681), .C2(new_n680), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT21), .B(G1986), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1991), .B(G1996), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT22), .B(G1981), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n688), .B(new_n689), .Z(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G229));
  INV_X1    g266(.A(KEYINPUT88), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G16), .B2(G23), .ZN(new_n693));
  OR3_X1    g268(.A1(new_n692), .A2(G16), .A3(G23), .ZN(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n693), .B(new_n694), .C1(G288), .C2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT33), .ZN(new_n697));
  INV_X1    g272(.A(G1976), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n695), .A2(G22), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G166), .B2(new_n695), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT89), .B(G1971), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n695), .A2(G6), .ZN(new_n704));
  INV_X1    g279(.A(G305), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(new_n705), .B2(new_n695), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT32), .B(G1981), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n699), .A2(new_n703), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT34), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n695), .A2(G24), .ZN(new_n711));
  INV_X1    g286(.A(G290), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(new_n695), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n713), .A2(G1986), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(G1986), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n478), .A2(G119), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n482), .A2(G131), .ZN(new_n717));
  NOR2_X1   g292(.A1(G95), .A2(G2105), .ZN(new_n718));
  OAI21_X1  g293(.A(G2104), .B1(new_n480), .B2(G107), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n716), .B(new_n717), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  MUX2_X1   g295(.A(G25), .B(new_n720), .S(G29), .Z(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT35), .B(G1991), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n721), .B(new_n723), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n714), .A2(new_n715), .A3(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(KEYINPUT91), .B1(new_n710), .B2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT34), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n709), .B(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT91), .ZN(new_n729));
  INV_X1    g304(.A(new_n725), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n726), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n726), .A2(new_n731), .A3(KEYINPUT90), .A4(KEYINPUT36), .ZN(new_n735));
  NOR2_X1   g310(.A1(G29), .A2(G35), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G162), .B2(G29), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT29), .ZN(new_n738));
  INV_X1    g313(.A(G2090), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G29), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n741), .A2(G26), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n478), .A2(G128), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n482), .A2(G140), .ZN(new_n744));
  NOR2_X1   g319(.A1(G104), .A2(G2105), .ZN(new_n745));
  OAI21_X1  g320(.A(G2104), .B1(new_n480), .B2(G116), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n743), .B(new_n744), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n742), .B1(new_n747), .B2(G29), .ZN(new_n748));
  MUX2_X1   g323(.A(new_n742), .B(new_n748), .S(KEYINPUT28), .Z(new_n749));
  INV_X1    g324(.A(G2067), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  AND2_X1   g326(.A1(KEYINPUT30), .A2(G28), .ZN(new_n752));
  NOR2_X1   g327(.A1(KEYINPUT30), .A2(G28), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n741), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n642), .B2(new_n741), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT93), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n758), .A2(G2105), .B1(G139), .B2(new_n482), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n480), .A2(G103), .A3(G2104), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT92), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT25), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G29), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G29), .B2(G33), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT94), .B(G2072), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT31), .B(G11), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n756), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n766), .B2(new_n767), .ZN(new_n771));
  NOR2_X1   g346(.A1(G29), .A2(G32), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n482), .A2(G141), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT96), .Z(new_n774));
  AND3_X1   g349(.A1(new_n480), .A2(G105), .A3(G2104), .ZN(new_n775));
  NAND3_X1  g350(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT26), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n775), .B(new_n777), .C1(new_n478), .C2(G129), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n772), .B1(new_n779), .B2(G29), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT27), .B(G1996), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n695), .A2(G5), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G171), .B2(new_n695), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(G1961), .Z(new_n785));
  INV_X1    g360(.A(G2078), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n741), .A2(G27), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G164), .B2(new_n741), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n554), .A2(G16), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G16), .B2(G19), .ZN(new_n791));
  INV_X1    g366(.A(G1341), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n786), .A2(new_n789), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n771), .A2(new_n782), .A3(new_n785), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n695), .A2(G21), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G168), .B2(new_n695), .ZN(new_n796));
  INV_X1    g371(.A(G1966), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(G160), .A2(G29), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT24), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(G34), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(G34), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n801), .A2(new_n802), .A3(new_n741), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(G2084), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(KEYINPUT95), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n807), .A2(KEYINPUT95), .B1(new_n788), .B2(G2078), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n627), .A2(G16), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G4), .B2(G16), .ZN(new_n811));
  INV_X1    g386(.A(G1348), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n798), .A2(new_n808), .A3(new_n809), .A4(new_n813), .ZN(new_n814));
  OAI22_X1  g389(.A1(new_n791), .A2(new_n792), .B1(new_n811), .B2(new_n812), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n794), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n734), .A2(new_n735), .A3(new_n740), .A4(new_n816), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n695), .A2(KEYINPUT23), .A3(G20), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT23), .ZN(new_n819));
  INV_X1    g394(.A(G20), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n820), .B2(G16), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n818), .B(new_n821), .C1(new_n623), .C2(new_n695), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G1956), .ZN(new_n823));
  INV_X1    g398(.A(new_n804), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n824), .A2(G2084), .ZN(new_n825));
  NOR3_X1   g400(.A1(new_n817), .A2(new_n823), .A3(new_n825), .ZN(G311));
  AND3_X1   g401(.A1(new_n734), .A2(new_n735), .A3(new_n816), .ZN(new_n827));
  INV_X1    g402(.A(new_n823), .ZN(new_n828));
  INV_X1    g403(.A(new_n825), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n827), .A2(new_n828), .A3(new_n829), .A4(new_n740), .ZN(G150));
  AOI22_X1  g405(.A1(new_n551), .A2(G93), .B1(G55), .B2(new_n515), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n531), .A2(new_n532), .A3(G67), .ZN(new_n832));
  NAND2_X1  g407(.A1(G80), .A2(G543), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(G651), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(G860), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT37), .Z(new_n838));
  NAND2_X1  g413(.A1(new_n627), .A2(G559), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT39), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT97), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n831), .A2(new_n835), .A3(new_n843), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n531), .A2(new_n532), .A3(G93), .A4(new_n513), .ZN(new_n845));
  INV_X1    g420(.A(G55), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n845), .B1(new_n846), .B2(new_n514), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n511), .B1(new_n832), .B2(new_n833), .ZN(new_n848));
  OAI21_X1  g423(.A(KEYINPUT97), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n553), .A2(new_n850), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n552), .A2(new_n550), .B1(new_n844), .B2(new_n849), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n842), .B(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n838), .B1(new_n856), .B2(G860), .ZN(G145));
  XNOR2_X1  g432(.A(new_n486), .B(KEYINPUT99), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n642), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(G160), .Z(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n493), .A2(new_n496), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n747), .B(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n764), .B(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n779), .ZN(new_n865));
  AOI22_X1  g440(.A1(G130), .A2(new_n478), .B1(new_n482), .B2(G142), .ZN(new_n866));
  OAI21_X1  g441(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n480), .A2(G118), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT100), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n866), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n720), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT101), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n872), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n873), .A2(new_n635), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n874), .ZN(new_n876));
  INV_X1    g451(.A(new_n635), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n865), .A2(new_n875), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT102), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n878), .A2(new_n875), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n865), .B(new_n882), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n861), .B(new_n881), .C1(new_n883), .C2(new_n880), .ZN(new_n884));
  INV_X1    g459(.A(G37), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n884), .B(new_n885), .C1(new_n883), .C2(new_n861), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g462(.A(new_n854), .B(new_n631), .Z(new_n888));
  NAND2_X1  g463(.A1(new_n623), .A2(new_n615), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n627), .A2(G299), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n890), .A3(KEYINPUT41), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n890), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT41), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n888), .A2(new_n891), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT103), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n623), .A2(new_n615), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n627), .A2(G299), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n889), .A2(new_n890), .A3(KEYINPUT103), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n895), .B1(new_n902), .B2(new_n888), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n903), .A2(KEYINPUT42), .ZN(new_n904));
  INV_X1    g479(.A(G288), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(G166), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(G290), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n906), .A2(G290), .ZN(new_n909));
  OAI21_X1  g484(.A(G305), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(G166), .B(G288), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n712), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n912), .A2(new_n705), .A3(new_n907), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n903), .A2(KEYINPUT42), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n904), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n915), .B1(new_n904), .B2(new_n916), .ZN(new_n918));
  OAI21_X1  g493(.A(G868), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n836), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n919), .B1(G868), .B2(new_n920), .ZN(G295));
  OAI21_X1  g496(.A(new_n919), .B1(G868), .B2(new_n920), .ZN(G331));
  INV_X1    g497(.A(KEYINPUT108), .ZN(new_n923));
  NAND2_X1  g498(.A1(G301), .A2(G168), .ZN(new_n924));
  NAND2_X1  g499(.A1(G286), .A2(G171), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n924), .A2(new_n851), .A3(new_n853), .A4(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(G286), .B1(new_n580), .B2(new_n581), .ZN(new_n927));
  AND2_X1   g502(.A1(G286), .A2(G171), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n553), .A2(new_n850), .ZN(new_n929));
  OAI22_X1  g504(.A1(new_n927), .A2(new_n928), .B1(new_n929), .B2(new_n852), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n926), .A2(new_n930), .A3(KEYINPUT105), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n894), .A2(new_n891), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT105), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n854), .B(new_n933), .C1(new_n927), .C2(new_n928), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n931), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n926), .A2(new_n930), .A3(new_n892), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n914), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(new_n885), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n931), .A2(new_n934), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n902), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n926), .A2(new_n930), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n932), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n939), .A2(KEYINPUT107), .A3(new_n902), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n942), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n912), .A2(new_n705), .A3(new_n907), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n705), .B1(new_n912), .B2(new_n907), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n910), .A2(KEYINPUT106), .A3(new_n913), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n938), .B1(new_n946), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n923), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n950), .A2(new_n951), .ZN(new_n956));
  AOI211_X1 g531(.A(new_n941), .B(new_n901), .C1(new_n931), .C2(new_n934), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT107), .B1(new_n939), .B2(new_n902), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n956), .B1(new_n959), .B2(new_n944), .ZN(new_n960));
  OAI211_X1 g535(.A(KEYINPUT108), .B(KEYINPUT43), .C1(new_n960), .C2(new_n938), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n935), .A2(new_n936), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n938), .B1(new_n963), .B2(new_n952), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n962), .B1(new_n964), .B2(new_n954), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n955), .A2(new_n961), .A3(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n967));
  AOI211_X1 g542(.A(KEYINPUT43), .B(new_n938), .C1(new_n946), .C2(new_n952), .ZN(new_n968));
  INV_X1    g543(.A(new_n938), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n952), .A2(new_n963), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n954), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n967), .B1(new_n968), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n966), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT109), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n966), .A2(KEYINPUT109), .A3(new_n972), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(G397));
  INV_X1    g552(.A(KEYINPUT62), .ZN(new_n978));
  INV_X1    g553(.A(G8), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT69), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n862), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G1384), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n493), .A2(KEYINPUT69), .A3(new_n496), .ZN(new_n983));
  XOR2_X1   g558(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n984));
  NAND4_X1  g559(.A1(new_n981), .A2(new_n982), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(G1384), .B1(new_n493), .B2(new_n496), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n986), .A2(KEYINPUT45), .ZN(new_n987));
  INV_X1    g562(.A(new_n468), .ZN(new_n988));
  INV_X1    g563(.A(new_n475), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n988), .B(G40), .C1(new_n989), .C2(new_n473), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n985), .A2(new_n987), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n797), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT50), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT50), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n990), .B1(new_n996), .B2(new_n986), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(new_n805), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n979), .B1(new_n993), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(G286), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n993), .A2(G168), .A3(new_n998), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n979), .A2(KEYINPUT122), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n1001), .A2(KEYINPUT51), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT51), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n978), .B(new_n1000), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n984), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n990), .B1(new_n994), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n986), .A2(KEYINPUT45), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(new_n786), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n995), .A2(new_n997), .ZN(new_n1011));
  XNOR2_X1  g586(.A(KEYINPUT123), .B(G1961), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n1009), .A2(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1010), .A2(G2078), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n985), .A2(new_n987), .A3(new_n991), .A4(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n618), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1005), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1981), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n592), .A2(new_n1020), .A3(new_n595), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1020), .B1(new_n592), .B2(new_n595), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT112), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT49), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n979), .B1(new_n991), .B2(new_n986), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT49), .ZN(new_n1026));
  OAI211_X1 g601(.A(KEYINPUT112), .B(new_n1026), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1024), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n991), .A2(new_n986), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1029), .B(G8), .C1(new_n698), .C2(G288), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT52), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT52), .B1(G288), .B2(new_n698), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1025), .B(new_n1032), .C1(new_n698), .C2(G288), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1028), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n497), .A2(new_n498), .A3(G1384), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n991), .B(new_n1008), .C1(new_n1035), .C2(new_n984), .ZN(new_n1036));
  INV_X1    g611(.A(G1971), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n995), .A2(new_n739), .A3(new_n997), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n979), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(G303), .A2(G8), .ZN(new_n1041));
  XOR2_X1   g616(.A(new_n1041), .B(KEYINPUT55), .Z(new_n1042));
  AOI21_X1  g617(.A(new_n1034), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n990), .B1(new_n1035), .B2(new_n996), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n862), .A2(new_n982), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT50), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(new_n739), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n979), .B1(new_n1048), .B2(new_n1038), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1044), .B1(new_n1049), .B2(new_n1042), .ZN(new_n1050));
  AOI21_X1  g625(.A(G1971), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n991), .B(new_n1047), .C1(new_n994), .C2(KEYINPUT50), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1052), .A2(G2090), .ZN(new_n1053));
  OAI21_X1  g628(.A(G8), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1042), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1054), .A2(KEYINPUT114), .A3(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1043), .A2(new_n1050), .A3(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT125), .B1(new_n1019), .B2(new_n1057), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1043), .A2(new_n1050), .A3(new_n1056), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT125), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1059), .A2(new_n1060), .A3(new_n1018), .A4(new_n1005), .ZN(new_n1061));
  OR2_X1    g636(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n1000), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT62), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1058), .A2(new_n1061), .A3(new_n1064), .ZN(new_n1065));
  XOR2_X1   g640(.A(KEYINPUT115), .B(KEYINPUT63), .Z(new_n1066));
  OR2_X1    g641(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1043), .A2(new_n1067), .A3(KEYINPUT63), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n999), .A2(G168), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1066), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1034), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1071), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n1025), .B(KEYINPUT113), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1028), .A2(new_n698), .A3(new_n905), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1073), .B1(new_n1074), .B2(new_n1021), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1070), .A2(new_n1072), .A3(new_n1075), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n1065), .A2(new_n1076), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1068), .A2(G168), .A3(new_n999), .ZN(new_n1078));
  INV_X1    g653(.A(G1956), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1052), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n994), .A2(new_n1006), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT56), .B(G2072), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1081), .A2(new_n991), .A3(new_n1008), .A4(new_n1082), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n563), .A2(new_n568), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1085), .B1(new_n563), .B2(new_n568), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1088), .B(new_n570), .C1(new_n575), .C2(new_n577), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT118), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1089), .A2(new_n1093), .A3(new_n1090), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n623), .A2(KEYINPUT57), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT119), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1089), .A2(new_n1093), .A3(new_n1090), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1093), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1099));
  OAI211_X1 g674(.A(KEYINPUT119), .B(new_n1096), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1084), .B1(new_n1097), .B2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1029), .A2(G2067), .ZN(new_n1103));
  AOI21_X1  g678(.A(G1348), .B1(new_n995), .B2(new_n997), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1102), .B(new_n627), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1096), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(new_n1100), .A3(new_n1109), .ZN(new_n1110));
  XOR2_X1   g685(.A(KEYINPUT58), .B(G1341), .Z(new_n1111));
  NAND2_X1  g686(.A1(new_n1029), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(new_n1036), .B2(G1996), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT120), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT120), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1115), .B(new_n1112), .C1(new_n1036), .C2(G1996), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1114), .A2(new_n554), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n1118));
  OR2_X1    g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1108), .A2(new_n1100), .A3(new_n1109), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1109), .B1(new_n1108), .B2(new_n1100), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1121), .A2(new_n1122), .A3(KEYINPUT61), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT61), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1124), .B1(new_n1102), .B2(new_n1110), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1119), .B(new_n1120), .C1(new_n1123), .C2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT60), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n1104), .B2(new_n1103), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n627), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT121), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1128), .A2(new_n1131), .A3(new_n627), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1104), .A2(new_n1103), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT60), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1130), .A2(KEYINPUT60), .A3(new_n1134), .A4(new_n1132), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1105), .B(new_n1110), .C1(new_n1126), .C2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1016), .A2(new_n618), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n986), .A2(new_n984), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n986), .A2(KEYINPUT45), .B1(G2105), .B2(new_n472), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1014), .B1(new_n468), .B2(KEYINPUT124), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1144), .B1(KEYINPUT124), .B2(new_n468), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1142), .A2(G40), .A3(new_n1143), .A4(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n542), .B1(new_n1013), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(KEYINPUT54), .B1(new_n1140), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT54), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1013), .A2(G301), .A3(new_n1146), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1017), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  AOI22_X1  g726(.A1(new_n1148), .A2(new_n1151), .B1(new_n1062), .B2(new_n1000), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1078), .B1(new_n1139), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1077), .B1(new_n1153), .B2(new_n1057), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n991), .A2(new_n1141), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1155), .A2(G1996), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n779), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1157), .A2(KEYINPUT111), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1157), .A2(KEYINPUT111), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1155), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n747), .B(new_n750), .ZN(new_n1161));
  INV_X1    g736(.A(G1996), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1161), .B1(new_n779), .B2(new_n1162), .ZN(new_n1163));
  AOI211_X1 g738(.A(new_n1158), .B(new_n1159), .C1(new_n1160), .C2(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n720), .B(new_n723), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1164), .B1(new_n1155), .B2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g741(.A(G290), .B(G1986), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1166), .B1(new_n1160), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1154), .A2(new_n1168), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1156), .A2(KEYINPUT46), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1156), .A2(KEYINPUT46), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1155), .B1(new_n779), .B2(new_n1161), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  XOR2_X1   g748(.A(new_n1173), .B(KEYINPUT47), .Z(new_n1174));
  NOR3_X1   g749(.A1(G290), .A2(G1986), .A3(new_n1155), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1175), .B(KEYINPUT127), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT48), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1174), .B1(new_n1166), .B2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n747), .A2(G2067), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n720), .A2(new_n722), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1179), .B1(new_n1164), .B2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(KEYINPUT126), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1178), .B1(new_n1182), .B2(new_n1160), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1169), .A2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g759(.A(G319), .B1(new_n968), .B2(new_n971), .ZN(new_n1186));
  NOR2_X1   g760(.A1(new_n1186), .A2(G229), .ZN(new_n1187));
  AOI21_X1  g761(.A(G227), .B1(new_n657), .B2(G14), .ZN(new_n1188));
  NAND3_X1  g762(.A1(new_n1187), .A2(new_n886), .A3(new_n1188), .ZN(G225));
  INV_X1    g763(.A(G225), .ZN(G308));
endmodule


