//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 1 0 1 0 1 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n562, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT67), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT68), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT69), .Z(G319));
  NAND2_X1  g033(.A1(G113), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n462), .A2(KEYINPUT70), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT3), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n472), .A2(G137), .A3(new_n473), .A4(new_n461), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n471), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n467), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  XOR2_X1   g052(.A(new_n477), .B(KEYINPUT71), .Z(G160));
  NAND3_X1  g053(.A1(new_n472), .A2(G2105), .A3(new_n461), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n472), .A2(new_n473), .A3(new_n461), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n473), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT72), .Z(new_n487));
  NAND3_X1  g062(.A1(new_n481), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR4_X1   g065(.A1(new_n464), .A2(KEYINPUT4), .A3(new_n490), .A4(G2105), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n472), .A2(G138), .A3(new_n473), .A4(new_n461), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(KEYINPUT4), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G114), .C2(new_n473), .ZN(new_n495));
  INV_X1    g070(.A(G126), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n495), .B1(new_n479), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n493), .A2(new_n497), .ZN(G164));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT75), .B1(new_n501), .B2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT75), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(new_n499), .A3(G543), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n500), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT74), .A2(G651), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT73), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT6), .ZN(new_n514));
  AOI21_X1  g089(.A(KEYINPUT73), .B1(KEYINPUT74), .B2(G651), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(G50), .A3(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n505), .A2(new_n516), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n508), .A2(new_n520), .ZN(G166));
  NAND2_X1  g096(.A1(new_n516), .A2(G89), .ZN(new_n522));
  INV_X1    g097(.A(G63), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n522), .B1(new_n523), .B2(new_n507), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(new_n505), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n516), .A2(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT76), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT76), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n516), .A2(new_n528), .A3(G543), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n527), .A2(G51), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  AND3_X1   g107(.A1(new_n525), .A2(new_n530), .A3(new_n532), .ZN(G168));
  AND3_X1   g108(.A1(new_n516), .A2(new_n528), .A3(G543), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n528), .B1(new_n516), .B2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  NOR3_X1   g111(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n505), .A2(new_n516), .A3(G90), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n539), .B2(new_n507), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT77), .ZN(new_n541));
  NOR3_X1   g116(.A1(new_n537), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n500), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n503), .B1(new_n499), .B2(G543), .ZN(new_n544));
  NOR3_X1   g119(.A1(new_n501), .A2(KEYINPUT75), .A3(KEYINPUT5), .ZN(new_n545));
  OAI211_X1 g120(.A(G64), .B(new_n543), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(G77), .A2(G543), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n507), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AND3_X1   g123(.A1(new_n505), .A2(new_n516), .A3(G90), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n527), .A2(G52), .A3(new_n529), .ZN(new_n551));
  AOI21_X1  g126(.A(KEYINPUT77), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n542), .A2(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  INV_X1    g129(.A(G43), .ZN(new_n555));
  NOR3_X1   g130(.A1(new_n534), .A2(new_n535), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n505), .A2(new_n516), .A3(G81), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n558), .B2(new_n507), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(G188));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G651), .ZN(new_n571));
  INV_X1    g146(.A(new_n518), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G91), .ZN(new_n573));
  INV_X1    g148(.A(G53), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT9), .B1(new_n526), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  NOR3_X1   g151(.A1(new_n526), .A2(KEYINPUT9), .A3(new_n574), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n571), .B(new_n573), .C1(new_n576), .C2(new_n577), .ZN(G299));
  NAND3_X1  g153(.A1(new_n525), .A2(new_n530), .A3(new_n532), .ZN(G286));
  OAI221_X1 g154(.A(new_n517), .B1(new_n518), .B2(new_n519), .C1(new_n506), .C2(new_n507), .ZN(G303));
  OAI21_X1  g155(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n505), .A2(new_n516), .A3(G87), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n516), .A2(G49), .A3(G543), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(G288));
  NAND3_X1  g159(.A1(new_n505), .A2(new_n516), .A3(G86), .ZN(new_n585));
  INV_X1    g160(.A(G48), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n505), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n587));
  OAI221_X1 g162(.A(new_n585), .B1(new_n526), .B2(new_n586), .C1(new_n587), .C2(new_n507), .ZN(G305));
  NOR2_X1   g163(.A1(new_n534), .A2(new_n535), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G47), .ZN(new_n590));
  NAND2_X1  g165(.A1(G72), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G60), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n568), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(G651), .A2(new_n593), .B1(new_n572), .B2(G85), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n590), .A2(new_n594), .ZN(G290));
  NAND3_X1  g170(.A1(new_n572), .A2(KEYINPUT10), .A3(G92), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  INV_X1    g172(.A(G92), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n518), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n568), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n596), .A2(new_n599), .B1(G651), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n589), .A2(G54), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G171), .B2(new_n606), .ZN(G284));
  OAI21_X1  g183(.A(new_n607), .B1(G171), .B2(new_n606), .ZN(G321));
  NOR2_X1   g184(.A1(G168), .A2(new_n606), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G299), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(KEYINPUT78), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(KEYINPUT78), .B2(new_n610), .ZN(G297));
  OAI21_X1  g190(.A(new_n614), .B1(KEYINPUT78), .B2(new_n610), .ZN(G280));
  INV_X1    g191(.A(new_n605), .ZN(new_n617));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G860), .ZN(G148));
  INV_X1    g194(.A(KEYINPUT79), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n617), .A2(new_n620), .A3(new_n618), .ZN(new_n621));
  OAI21_X1  g196(.A(KEYINPUT79), .B1(new_n605), .B2(G559), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G868), .B2(new_n560), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g201(.A1(new_n480), .A2(G123), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n483), .A2(G135), .ZN(new_n628));
  OR2_X1    g203(.A1(G99), .A2(G2105), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n629), .B(G2104), .C1(G111), .C2(new_n473), .ZN(new_n630));
  AND3_X1   g205(.A1(new_n627), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2096), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n475), .A2(new_n461), .A3(new_n463), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT12), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT80), .B(G2100), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n634), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n632), .A2(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(KEYINPUT15), .B(G2435), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT82), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2438), .Z(new_n643));
  XOR2_X1   g218(.A(G2427), .B(G2430), .Z(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(new_n646), .A3(KEYINPUT14), .ZN(new_n647));
  XOR2_X1   g222(.A(G2451), .B(G2454), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT81), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT16), .Z(new_n650));
  OR2_X1    g225(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n647), .A2(new_n650), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n651), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n653), .B1(new_n651), .B2(new_n654), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n640), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n659), .A2(new_n639), .A3(new_n655), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n658), .A2(new_n660), .A3(G14), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT83), .Z(G401));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2067), .B(G2678), .Z(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(new_n667), .A3(KEYINPUT17), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT84), .B(KEYINPUT18), .Z(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n666), .B2(new_n669), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n671), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2096), .B(G2100), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  INV_X1    g251(.A(KEYINPUT20), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT85), .ZN(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n677), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n679), .A2(new_n680), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n685), .A2(new_n683), .A3(new_n681), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n679), .A2(KEYINPUT20), .A3(new_n680), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n684), .B(new_n686), .C1(new_n688), .C2(new_n683), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT86), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n691), .B(new_n692), .Z(new_n693));
  AND2_X1   g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n690), .A2(new_n693), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1981), .B(G1986), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n697), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(new_n694), .B2(new_n695), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n698), .A2(new_n700), .ZN(G229));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G25), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n480), .A2(G119), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n483), .A2(G131), .ZN(new_n705));
  OR2_X1    g280(.A1(G95), .A2(G2105), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n706), .B(G2104), .C1(G107), .C2(new_n473), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT87), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n704), .A2(new_n705), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n703), .B1(new_n710), .B2(new_n702), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT35), .B(G1991), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n711), .B(new_n712), .Z(new_n713));
  INV_X1    g288(.A(G1986), .ZN(new_n714));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n715), .A2(G24), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G290), .B2(G16), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n713), .B1(new_n714), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT88), .B(KEYINPUT34), .ZN(new_n719));
  INV_X1    g294(.A(G22), .ZN(new_n720));
  OAI21_X1  g295(.A(KEYINPUT90), .B1(new_n720), .B2(G16), .ZN(new_n721));
  OR3_X1    g296(.A1(new_n720), .A2(KEYINPUT90), .A3(G16), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n721), .B(new_n722), .C1(G166), .C2(new_n715), .ZN(new_n723));
  INV_X1    g298(.A(G1971), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n715), .A2(G6), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n587), .A2(new_n507), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n585), .B1(new_n586), .B2(new_n526), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n726), .B1(new_n729), .B2(new_n715), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT32), .B(G1981), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(KEYINPUT89), .B1(G16), .B2(G23), .ZN(new_n733));
  OR3_X1    g308(.A1(KEYINPUT89), .A2(G16), .A3(G23), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n733), .B(new_n734), .C1(G288), .C2(new_n715), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT33), .B(G1976), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n725), .A2(new_n732), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n718), .B1(new_n719), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n717), .A2(new_n714), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n739), .B(new_n740), .C1(new_n719), .C2(new_n738), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT91), .B(KEYINPUT36), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n741), .B(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT97), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n702), .A2(G33), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT25), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G139), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n749), .B1(new_n482), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT93), .ZN(new_n752));
  INV_X1    g327(.A(new_n464), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n753), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(new_n473), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n746), .B1(new_n757), .B2(new_n702), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(G2072), .Z(new_n759));
  OR2_X1    g334(.A1(KEYINPUT24), .A2(G34), .ZN(new_n760));
  NAND2_X1  g335(.A1(KEYINPUT24), .A2(G34), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n760), .A2(new_n702), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G160), .B2(new_n702), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(G2084), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  OR2_X1    g340(.A1(G29), .A2(G32), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n483), .A2(G141), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT94), .ZN(new_n768));
  NAND3_X1  g343(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT95), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT26), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n480), .A2(G129), .B1(G105), .B2(new_n475), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n768), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n766), .B1(new_n773), .B2(new_n702), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT27), .B(G1996), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT96), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n745), .B1(new_n765), .B2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n777), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n779), .A2(KEYINPUT97), .A3(new_n764), .A4(new_n759), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(G168), .A2(G16), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G16), .B2(G21), .ZN(new_n783));
  INV_X1    g358(.A(G1966), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n631), .A2(G29), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT98), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT30), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n702), .B1(new_n790), .B2(G28), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n790), .B2(G28), .ZN(new_n792));
  NOR4_X1   g367(.A1(new_n785), .A2(new_n786), .A3(new_n789), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n715), .A2(G4), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n617), .B2(new_n715), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(G1348), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT31), .B(G11), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n715), .A2(G19), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n560), .B2(new_n715), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT92), .B(G1341), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n793), .A2(new_n796), .A3(new_n797), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n715), .A2(G5), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G171), .B2(new_n715), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n804), .A2(G1961), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n715), .A2(G20), .ZN(new_n806));
  OAI211_X1 g381(.A(KEYINPUT23), .B(new_n806), .C1(new_n612), .C2(new_n715), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(KEYINPUT23), .B2(new_n806), .ZN(new_n808));
  INV_X1    g383(.A(G1956), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n702), .A2(G26), .ZN(new_n811));
  OR2_X1    g386(.A1(G104), .A2(G2105), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n812), .B(G2104), .C1(G116), .C2(new_n473), .ZN(new_n813));
  INV_X1    g388(.A(G140), .ZN(new_n814));
  INV_X1    g389(.A(G128), .ZN(new_n815));
  OAI221_X1 g390(.A(new_n813), .B1(new_n482), .B2(new_n814), .C1(new_n815), .C2(new_n479), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n811), .B1(new_n817), .B2(new_n702), .ZN(new_n818));
  MUX2_X1   g393(.A(new_n811), .B(new_n818), .S(KEYINPUT28), .Z(new_n819));
  OR2_X1    g394(.A1(new_n819), .A2(G2067), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n702), .A2(G35), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G162), .B2(new_n702), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT29), .B(G2090), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n795), .A2(G1348), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n819), .A2(G2067), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n820), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  NOR4_X1   g402(.A1(new_n802), .A2(new_n805), .A3(new_n810), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n702), .A2(G27), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(G164), .B2(new_n702), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT100), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(G2078), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n763), .A2(G2084), .ZN(new_n833));
  OAI221_X1 g408(.A(new_n833), .B1(new_n774), .B2(new_n775), .C1(G1961), .C2(new_n804), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT99), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n781), .A2(new_n828), .A3(new_n832), .A4(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(KEYINPUT101), .B1(new_n744), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n741), .B(new_n742), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n828), .A2(new_n832), .A3(new_n835), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT101), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n838), .A2(new_n839), .A3(new_n840), .A4(new_n781), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n837), .A2(new_n841), .ZN(G311));
  NAND3_X1  g417(.A1(new_n838), .A2(new_n781), .A3(new_n839), .ZN(G150));
  NOR2_X1   g418(.A1(new_n605), .A2(new_n618), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  AND3_X1   g420(.A1(new_n505), .A2(new_n516), .A3(G81), .ZN(new_n846));
  NAND2_X1  g421(.A1(G68), .A2(G543), .ZN(new_n847));
  INV_X1    g422(.A(G56), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n847), .B1(new_n568), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n846), .B1(new_n849), .B2(G651), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n527), .A2(G43), .A3(new_n529), .ZN(new_n851));
  INV_X1    g426(.A(G55), .ZN(new_n852));
  NOR3_X1   g427(.A1(new_n534), .A2(new_n535), .A3(new_n852), .ZN(new_n853));
  AOI22_X1  g428(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n854));
  INV_X1    g429(.A(G93), .ZN(new_n855));
  OAI22_X1  g430(.A1(new_n854), .A2(new_n507), .B1(new_n855), .B2(new_n518), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n850), .B(new_n851), .C1(new_n853), .C2(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n527), .A2(G55), .A3(new_n529), .ZN(new_n858));
  OAI211_X1 g433(.A(G67), .B(new_n543), .C1(new_n544), .C2(new_n545), .ZN(new_n859));
  NAND2_X1  g434(.A1(G80), .A2(G543), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n507), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AND3_X1   g436(.A1(new_n505), .A2(new_n516), .A3(G93), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g438(.A(new_n858), .B(new_n863), .C1(new_n556), .C2(new_n559), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n857), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT39), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n845), .B(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(G860), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT102), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n853), .A2(new_n856), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n871), .A2(new_n868), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT37), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n870), .A2(new_n873), .ZN(G145));
  XNOR2_X1  g449(.A(G160), .B(new_n488), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(new_n631), .Z(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n756), .A2(G164), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n756), .A2(G164), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(new_n816), .A3(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n816), .B1(new_n878), .B2(new_n879), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n773), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n882), .ZN(new_n884));
  INV_X1    g459(.A(new_n773), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n885), .A3(new_n880), .ZN(new_n886));
  INV_X1    g461(.A(G130), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n479), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT104), .ZN(new_n889));
  OR2_X1    g464(.A1(G106), .A2(G2105), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n890), .B(G2104), .C1(G118), .C2(new_n473), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n483), .A2(G142), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n894), .B(KEYINPUT103), .Z(new_n895));
  AOI21_X1  g470(.A(new_n634), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n893), .A2(new_n895), .A3(new_n634), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(new_n710), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n898), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n709), .B1(new_n900), .B2(new_n896), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n883), .A2(new_n886), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n902), .B1(new_n883), .B2(new_n886), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n903), .B1(new_n904), .B2(KEYINPUT105), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n906));
  AOI211_X1 g481(.A(new_n906), .B(new_n902), .C1(new_n883), .C2(new_n886), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n877), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(G37), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n903), .A2(new_n876), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n910), .A2(new_n904), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n908), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g488(.A(KEYINPUT106), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n590), .A2(new_n594), .A3(G288), .ZN(new_n915));
  AOI21_X1  g490(.A(G288), .B1(new_n590), .B2(new_n594), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(G288), .ZN(new_n918));
  NAND2_X1  g493(.A1(G290), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n590), .A2(new_n594), .A3(G288), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(KEYINPUT106), .A3(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(G303), .B(G305), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n917), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(G166), .B(G305), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n924), .A2(KEYINPUT106), .A3(new_n919), .A4(new_n920), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n923), .A2(KEYINPUT107), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT107), .B1(new_n923), .B2(new_n925), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT42), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT41), .ZN(new_n930));
  NAND3_X1  g505(.A1(G299), .A2(new_n604), .A3(new_n603), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(G299), .B1(new_n604), .B2(new_n603), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n605), .A2(new_n612), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n935), .A2(KEYINPUT41), .A3(new_n931), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n623), .A2(new_n865), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n857), .A2(new_n864), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n938), .B1(new_n621), .B2(new_n622), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n934), .B(new_n936), .C1(new_n937), .C2(new_n939), .ZN(new_n940));
  OR2_X1    g515(.A1(new_n937), .A2(new_n939), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n935), .A2(new_n931), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT42), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n923), .A2(new_n944), .A3(new_n925), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n929), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n943), .B1(new_n929), .B2(new_n945), .ZN(new_n947));
  OAI21_X1  g522(.A(G868), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n871), .A2(G868), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(KEYINPUT108), .ZN(G295));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n951), .B(new_n953), .ZN(G331));
  NOR3_X1   g529(.A1(new_n542), .A2(new_n552), .A3(G286), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n541), .B1(new_n537), .B2(new_n540), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n550), .A2(new_n551), .A3(KEYINPUT77), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n589), .A2(G51), .B1(new_n505), .B2(new_n524), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n956), .A2(new_n957), .B1(new_n958), .B2(new_n532), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n865), .B1(new_n955), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT110), .ZN(new_n961));
  OAI21_X1  g536(.A(G286), .B1(new_n542), .B2(new_n552), .ZN(new_n962));
  NAND3_X1  g537(.A1(G168), .A2(new_n956), .A3(new_n957), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n938), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n960), .A2(new_n961), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n934), .A2(new_n936), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n938), .A2(new_n962), .A3(KEYINPUT110), .A4(new_n963), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT111), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n960), .A2(new_n942), .A3(new_n964), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n965), .A2(new_n966), .A3(new_n971), .A4(new_n967), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n969), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n973), .A2(new_n928), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n926), .A2(new_n927), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n969), .A2(new_n975), .A3(new_n970), .A4(new_n972), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n909), .ZN(new_n977));
  OR3_X1    g552(.A1(new_n974), .A2(new_n977), .A3(KEYINPUT43), .ZN(new_n978));
  AOI22_X1  g553(.A1(new_n934), .A2(new_n936), .B1(new_n960), .B2(new_n964), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n965), .A2(new_n967), .B1(new_n935), .B2(new_n931), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n928), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n981), .A2(new_n976), .A3(new_n909), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT113), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n982), .A2(KEYINPUT113), .A3(KEYINPUT43), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n978), .A2(new_n985), .A3(KEYINPUT44), .A4(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT43), .B1(new_n974), .B2(new_n977), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT43), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n981), .A2(new_n976), .A3(new_n990), .A4(new_n909), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n988), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AOI211_X1 g569(.A(KEYINPUT112), .B(KEYINPUT44), .C1(new_n989), .C2(new_n991), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n987), .B1(new_n994), .B2(new_n995), .ZN(G397));
  INV_X1    g571(.A(G1384), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(new_n493), .B2(new_n497), .ZN(new_n998));
  XNOR2_X1  g573(.A(KEYINPUT114), .B(KEYINPUT45), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n467), .A2(new_n474), .A3(G40), .A4(new_n476), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n773), .B(G1996), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n816), .B(G2067), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1005), .B(KEYINPUT116), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n709), .B(new_n712), .ZN(new_n1008));
  XOR2_X1   g583(.A(new_n1008), .B(KEYINPUT117), .Z(new_n1009));
  OAI21_X1  g584(.A(new_n1003), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  NOR4_X1   g585(.A1(new_n1001), .A2(G290), .A3(G1986), .A4(new_n1002), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1003), .A2(G1986), .A3(G290), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1014), .B(KEYINPUT115), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n1010), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1001), .A2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g595(.A(KEYINPUT45), .B(new_n997), .C1(new_n493), .C2(new_n497), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1002), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n998), .A2(KEYINPUT118), .A3(new_n1000), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1020), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1018), .B1(new_n1025), .B2(G2078), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n998), .A2(KEYINPUT50), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT50), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1028), .B(new_n997), .C1(new_n493), .C2(new_n497), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n1027), .A2(new_n1022), .A3(new_n1029), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n1030), .A2(G1961), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT45), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n998), .A2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1033), .B(new_n1022), .C1(new_n998), .C2(new_n1000), .ZN(new_n1034));
  OR2_X1    g609(.A1(new_n1018), .A2(G2078), .ZN(new_n1035));
  OR2_X1    g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1026), .A2(new_n1031), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1017), .B1(new_n1037), .B2(G301), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n474), .A2(G40), .A3(new_n476), .ZN(new_n1039));
  OR2_X1    g614(.A1(new_n466), .A2(KEYINPUT125), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n473), .B1(new_n466), .B2(KEYINPUT125), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1035), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1001), .A2(new_n1039), .A3(new_n1021), .A4(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1026), .A2(new_n1031), .A3(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1038), .B1(G301), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1037), .A2(G171), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT124), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT124), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1037), .A2(new_n1048), .A3(G171), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1017), .B1(new_n1044), .B2(G171), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1045), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT57), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n576), .A2(new_n577), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1053), .B1(new_n1054), .B2(KEYINPUT122), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n1055), .B(new_n612), .ZN(new_n1056));
  XOR2_X1   g631(.A(KEYINPUT56), .B(G2072), .Z(new_n1057));
  XNOR2_X1  g632(.A(new_n1057), .B(KEYINPUT123), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1020), .A2(new_n1023), .A3(new_n1024), .A4(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1027), .A2(new_n1022), .A3(new_n1029), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n809), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1056), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(G1348), .ZN(new_n1063));
  INV_X1    g638(.A(G2067), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n998), .A2(new_n1002), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n1060), .A2(new_n1063), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1066), .A2(new_n605), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1062), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n1055), .B(G299), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT61), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1071), .A2(new_n1072), .A3(new_n1062), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1072), .B1(new_n1071), .B2(new_n1062), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n998), .A2(G2067), .A3(new_n1002), .ZN(new_n1076));
  AOI211_X1 g651(.A(new_n1076), .B(new_n617), .C1(new_n1060), .C2(new_n1063), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT60), .B1(new_n1067), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT60), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1066), .A2(new_n1079), .A3(new_n617), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT58), .B(G1341), .ZN(new_n1081));
  OAI22_X1  g656(.A1(new_n1025), .A2(G1996), .B1(new_n1065), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1082), .A2(new_n1083), .A3(new_n560), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1083), .B1(new_n1082), .B2(new_n560), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1078), .B(new_n1080), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1068), .B(new_n1071), .C1(new_n1075), .C2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1981), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n729), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(G305), .A2(G1981), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT49), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT49), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1089), .A2(new_n1090), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(G8), .B1(new_n998), .B2(new_n1002), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT121), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT121), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1098), .B(G8), .C1(new_n998), .C2(new_n1002), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1095), .A2(new_n1100), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1097), .A2(new_n1099), .B1(G1976), .B2(new_n918), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT52), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(G1976), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT52), .B1(G288), .B2(new_n1105), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1102), .A2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(G2090), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1025), .A2(new_n724), .B1(new_n1030), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G8), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT119), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n1115));
  NAND4_X1  g690(.A1(G303), .A2(new_n1115), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT120), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(G166), .A2(new_n1111), .ZN(new_n1120));
  OR2_X1    g695(.A1(new_n1120), .A2(KEYINPUT55), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1114), .A2(KEYINPUT120), .A3(new_n1116), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1119), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1112), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1123), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1108), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  OR2_X1    g702(.A1(new_n1060), .A2(G2084), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1034), .A2(new_n784), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(G168), .A2(new_n1111), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT51), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1111), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1131), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1133), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1134), .A2(KEYINPUT51), .A3(new_n1131), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1132), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1052), .A2(new_n1087), .A3(new_n1127), .A4(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1101), .A2(new_n1105), .A3(new_n918), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1141), .A2(new_n1089), .B1(new_n1099), .B2(new_n1097), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1127), .A2(KEYINPUT63), .A3(G168), .A4(new_n1134), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT63), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1108), .A2(new_n1124), .A3(new_n1126), .A4(new_n1134), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1144), .B1(new_n1145), .B2(G286), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1142), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1140), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1108), .A2(new_n1126), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1139), .A2(KEYINPUT62), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT62), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1151), .B(new_n1132), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1150), .A2(new_n1050), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1149), .B1(new_n1153), .B2(new_n1124), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1016), .B1(new_n1148), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1003), .B1(new_n1006), .B2(new_n773), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1001), .A2(G1996), .A3(new_n1002), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n1157), .A2(KEYINPUT46), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(KEYINPUT46), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1156), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT47), .ZN(new_n1161));
  XOR2_X1   g736(.A(new_n1011), .B(KEYINPUT48), .Z(new_n1162));
  NAND2_X1  g737(.A1(new_n1010), .A2(new_n1162), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n709), .A2(new_n712), .ZN(new_n1164));
  OAI22_X1  g739(.A1(new_n1007), .A2(new_n1164), .B1(G2067), .B2(new_n816), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(new_n1003), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1161), .A2(new_n1163), .A3(new_n1166), .ZN(new_n1167));
  XOR2_X1   g742(.A(new_n1167), .B(KEYINPUT126), .Z(new_n1168));
  NAND2_X1  g743(.A1(new_n1155), .A2(new_n1168), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g744(.A(G227), .ZN(new_n1171));
  INV_X1    g745(.A(new_n457), .ZN(new_n1172));
  AOI21_X1  g746(.A(new_n1172), .B1(new_n698), .B2(new_n700), .ZN(new_n1173));
  NAND3_X1  g747(.A1(new_n661), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g748(.A1(new_n1174), .A2(KEYINPUT127), .ZN(new_n1175));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n1176));
  NAND4_X1  g750(.A1(new_n661), .A2(new_n1176), .A3(new_n1171), .A4(new_n1173), .ZN(new_n1177));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g752(.A1(new_n1178), .A2(new_n912), .A3(new_n992), .ZN(G225));
  INV_X1    g753(.A(G225), .ZN(G308));
endmodule


