//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 0 0 1 1 1 1 1 1 1 1 1 0 1 0 1 0 1 0 0 1 1 1 0 0 1 1 1 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT70), .ZN(new_n189));
  NOR2_X1   g003(.A1(KEYINPUT2), .A2(G113), .ZN(new_n190));
  AOI21_X1  g004(.A(KEYINPUT66), .B1(KEYINPUT2), .B2(G113), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  NAND3_X1  g006(.A1(KEYINPUT66), .A2(KEYINPUT2), .A3(G113), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n190), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G116), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G119), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT67), .B(G119), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n194), .B(new_n196), .C1(new_n195), .C2(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n196), .B1(new_n197), .B2(new_n195), .ZN(new_n199));
  INV_X1    g013(.A(new_n193), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(new_n191), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n199), .B1(new_n190), .B2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT69), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n198), .A2(new_n202), .A3(KEYINPUT69), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G134), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n208), .A2(KEYINPUT65), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(KEYINPUT65), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT11), .ZN(new_n211));
  OAI22_X1  g025(.A1(new_n209), .A2(new_n210), .B1(new_n211), .B2(G137), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  INV_X1    g027(.A(G137), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(KEYINPUT11), .A3(G134), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n211), .A2(G137), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n212), .A2(new_n213), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(G134), .A2(G137), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT65), .B(G134), .ZN(new_n219));
  OAI211_X1 g033(.A(G131), .B(new_n218), .C1(new_n219), .C2(G137), .ZN(new_n220));
  INV_X1    g034(.A(G146), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G143), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G128), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT64), .B(G143), .ZN(new_n227));
  AOI211_X1 g041(.A(new_n223), .B(new_n226), .C1(new_n227), .C2(G146), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n224), .B1(new_n222), .B2(KEYINPUT1), .ZN(new_n229));
  OR2_X1    g043(.A1(KEYINPUT64), .A2(G143), .ZN(new_n230));
  NAND2_X1  g044(.A1(KEYINPUT64), .A2(G143), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n221), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G143), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G146), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n229), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n217), .B(new_n220), .C1(new_n228), .C2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n211), .A2(G137), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n215), .B(new_n216), .C1(new_n219), .C2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G131), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(new_n217), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT0), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n242), .A2(new_n224), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n243), .B1(new_n232), .B2(new_n234), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n224), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n223), .B1(new_n227), .B2(G146), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n244), .A2(new_n245), .B1(new_n246), .B2(new_n243), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n237), .B1(new_n241), .B2(new_n247), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n241), .A2(new_n237), .A3(new_n247), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n207), .B(new_n236), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n241), .A2(new_n247), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT30), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n252), .A2(new_n236), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n236), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n252), .A2(KEYINPUT68), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n241), .A2(new_n237), .A3(new_n247), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n255), .B1(new_n259), .B2(new_n253), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n251), .B1(new_n260), .B2(new_n203), .ZN(new_n261));
  NOR2_X1   g075(.A1(G237), .A2(G953), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G210), .ZN(new_n263));
  XOR2_X1   g077(.A(new_n263), .B(KEYINPUT27), .Z(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(KEYINPUT26), .ZN(new_n265));
  INV_X1    g079(.A(G101), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n265), .B(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n189), .B1(new_n261), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n236), .B1(new_n249), .B2(new_n248), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n254), .B1(new_n269), .B2(KEYINPUT30), .ZN(new_n270));
  INV_X1    g084(.A(new_n203), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n250), .B(new_n267), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n272), .A2(KEYINPUT70), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT31), .B1(new_n268), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n267), .ZN(new_n275));
  XOR2_X1   g089(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n276));
  NAND2_X1  g090(.A1(new_n252), .A2(new_n236), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n203), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n276), .B1(new_n250), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT28), .ZN(new_n280));
  INV_X1    g094(.A(new_n207), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n280), .B1(new_n281), .B2(new_n277), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n275), .B1(new_n279), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n284), .B1(new_n272), .B2(KEYINPUT31), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n188), .B1(new_n274), .B2(new_n286), .ZN(new_n287));
  XOR2_X1   g101(.A(KEYINPUT72), .B(KEYINPUT32), .Z(new_n288));
  OAI21_X1  g102(.A(KEYINPUT73), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT31), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n272), .A2(KEYINPUT70), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n260), .A2(new_n203), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n292), .A2(new_n189), .A3(new_n250), .A4(new_n267), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n290), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  OAI211_X1 g108(.A(KEYINPUT32), .B(new_n187), .C1(new_n294), .C2(new_n285), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n269), .A2(new_n281), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(new_n250), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n283), .B1(new_n297), .B2(KEYINPUT28), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT29), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n275), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(G902), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n299), .B1(new_n261), .B2(new_n267), .ZN(new_n302));
  NOR3_X1   g116(.A1(new_n279), .A2(new_n275), .A3(new_n283), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G472), .ZN(new_n305));
  AND2_X1   g119(.A1(new_n295), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n187), .B1(new_n294), .B2(new_n285), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT73), .ZN(new_n308));
  INV_X1    g122(.A(new_n288), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n289), .A2(new_n306), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G953), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(G221), .A3(G234), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n313), .B(KEYINPUT22), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n314), .B(G137), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT24), .B(G110), .ZN(new_n316));
  INV_X1    g130(.A(G119), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT67), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT67), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G119), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n224), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n317), .A2(G128), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n316), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT23), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n324), .A2(G128), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G119), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(G128), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n326), .B(new_n327), .C1(new_n197), .C2(new_n325), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n323), .B1(new_n328), .B2(G110), .ZN(new_n329));
  INV_X1    g143(.A(G140), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G125), .ZN(new_n331));
  INV_X1    g145(.A(G125), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G140), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n331), .A2(new_n333), .A3(KEYINPUT16), .ZN(new_n334));
  OR3_X1    g148(.A1(new_n332), .A2(KEYINPUT16), .A3(G140), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n334), .A2(G146), .A3(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n331), .A2(new_n333), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n221), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n329), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT74), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n319), .A2(G119), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n317), .A2(KEYINPUT67), .ZN(new_n343));
  OAI22_X1  g157(.A1(new_n342), .A2(new_n343), .B1(new_n324), .B2(G128), .ZN(new_n344));
  INV_X1    g158(.A(G110), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n344), .A2(new_n345), .A3(new_n327), .A4(new_n326), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n336), .B1(new_n346), .B2(new_n323), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT74), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n348), .A3(new_n339), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n341), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(G146), .B1(new_n334), .B2(new_n335), .ZN(new_n351));
  INV_X1    g165(.A(new_n322), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n352), .B1(new_n197), .B2(new_n224), .ZN(new_n353));
  OAI22_X1  g167(.A1(new_n336), .A2(new_n351), .B1(new_n353), .B2(new_n316), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n328), .A2(G110), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n315), .B1(new_n350), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n315), .ZN(new_n359));
  AOI211_X1 g173(.A(new_n356), .B(new_n359), .C1(new_n341), .C2(new_n349), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT75), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT25), .ZN(new_n363));
  INV_X1    g177(.A(G902), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n361), .A2(new_n362), .A3(new_n363), .A4(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G217), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n366), .B1(G234), .B2(new_n364), .ZN(new_n367));
  AND4_X1   g181(.A1(new_n348), .A2(new_n329), .A3(new_n337), .A4(new_n339), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n348), .B1(new_n347), .B2(new_n339), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n357), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n359), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n350), .A2(new_n357), .A3(new_n315), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n364), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n362), .A2(new_n363), .ZN(new_n374));
  NAND2_X1  g188(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n365), .A2(new_n367), .A3(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n367), .A2(G902), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n371), .A2(new_n372), .A3(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(KEYINPUT76), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT77), .B1(new_n311), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(KEYINPUT100), .A2(G952), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(KEYINPUT100), .A2(G952), .ZN(new_n386));
  AOI21_X1  g200(.A(G953), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(G234), .A2(G237), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  XOR2_X1   g203(.A(KEYINPUT21), .B(G898), .Z(new_n390));
  NAND3_X1  g204(.A1(new_n388), .A2(G902), .A3(G953), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G475), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n338), .B(new_n221), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT18), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n262), .A2(G214), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT89), .B1(new_n396), .B2(new_n233), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n227), .A2(new_n396), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT89), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n262), .A2(new_n399), .A3(G143), .A4(G214), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n397), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G131), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n397), .A2(new_n398), .A3(new_n213), .A4(new_n400), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n397), .A2(new_n398), .A3(new_n395), .A4(new_n400), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(new_n404), .A3(KEYINPUT90), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT90), .B1(new_n403), .B2(new_n404), .ZN(new_n407));
  OAI221_X1 g221(.A(new_n394), .B1(new_n395), .B2(new_n402), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT17), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n402), .A2(new_n409), .A3(new_n403), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n336), .A2(new_n351), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n401), .A2(KEYINPUT17), .A3(G131), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(G113), .B(G122), .ZN(new_n415));
  INV_X1    g229(.A(G104), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n415), .B(new_n416), .ZN(new_n417));
  OR2_X1    g231(.A1(new_n417), .A2(KEYINPUT94), .ZN(new_n418));
  OR2_X1    g232(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(G902), .B1(new_n414), .B2(new_n418), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n393), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT91), .ZN(new_n422));
  INV_X1    g236(.A(new_n417), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n423), .B1(new_n408), .B2(new_n413), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n394), .B1(new_n402), .B2(new_n395), .ZN(new_n425));
  INV_X1    g239(.A(new_n407), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n425), .B1(new_n426), .B2(new_n405), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n338), .B(KEYINPUT19), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n336), .B1(new_n428), .B2(new_n221), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n402), .A2(new_n403), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n423), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n427), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n422), .B1(new_n424), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n413), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n417), .B1(new_n435), .B2(new_n427), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n436), .B(KEYINPUT91), .C1(new_n427), .C2(new_n432), .ZN(new_n437));
  NOR2_X1   g251(.A1(G475), .A2(G902), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(KEYINPUT92), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n434), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT20), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n424), .A2(new_n433), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n439), .B1(KEYINPUT93), .B2(KEYINPUT20), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n442), .B(new_n443), .C1(KEYINPUT93), .C2(new_n439), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n421), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G122), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G116), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(KEYINPUT95), .ZN(new_n448));
  XOR2_X1   g262(.A(KEYINPUT80), .B(G107), .Z(new_n449));
  NAND2_X1  g263(.A1(new_n195), .A2(G122), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n448), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n450), .B(KEYINPUT14), .ZN(new_n453));
  OAI21_X1  g267(.A(G107), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n224), .A2(G143), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(KEYINPUT97), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT96), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n457), .B1(new_n227), .B2(G128), .ZN(new_n458));
  AND2_X1   g272(.A1(KEYINPUT64), .A2(G143), .ZN(new_n459));
  NOR2_X1   g273(.A1(KEYINPUT64), .A2(G143), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n457), .B(G128), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n456), .B1(new_n458), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT98), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n459), .A2(new_n460), .ZN(new_n466));
  OAI21_X1  g280(.A(KEYINPUT96), .B1(new_n466), .B2(new_n224), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n461), .ZN(new_n468));
  AOI21_X1  g282(.A(KEYINPUT98), .B1(new_n468), .B2(new_n456), .ZN(new_n469));
  INV_X1    g283(.A(new_n219), .ZN(new_n470));
  NOR3_X1   g284(.A1(new_n465), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n463), .A2(new_n464), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n468), .A2(KEYINPUT98), .A3(new_n456), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n219), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n451), .B(new_n454), .C1(new_n471), .C2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT13), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n468), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n456), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n468), .A2(new_n476), .ZN(new_n479));
  OAI21_X1  g293(.A(G134), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n470), .B1(new_n465), .B2(new_n469), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n448), .A2(new_n450), .ZN(new_n482));
  XOR2_X1   g296(.A(new_n482), .B(new_n449), .Z(new_n483));
  NAND3_X1  g297(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  XOR2_X1   g298(.A(KEYINPUT9), .B(G234), .Z(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NOR3_X1   g300(.A1(new_n486), .A2(new_n366), .A3(G953), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n475), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n487), .B1(new_n475), .B2(new_n484), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n364), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G478), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n491), .A2(KEYINPUT15), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n492), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n364), .B(new_n494), .C1(new_n488), .C2(new_n489), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n493), .A2(KEYINPUT99), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(KEYINPUT99), .B1(new_n493), .B2(new_n495), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n392), .B(new_n445), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT101), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT99), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n475), .A2(new_n484), .ZN(new_n502));
  INV_X1    g316(.A(new_n487), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n475), .A2(new_n484), .A3(new_n487), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n494), .B1(new_n506), .B2(new_n364), .ZN(new_n507));
  INV_X1    g321(.A(new_n495), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n501), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n493), .A2(new_n495), .A3(KEYINPUT99), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n511), .A2(KEYINPUT101), .A3(new_n392), .A4(new_n445), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n500), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(G214), .B1(G237), .B2(G902), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n246), .A2(new_n225), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n232), .A2(new_n234), .ZN(new_n517));
  INV_X1    g331(.A(new_n229), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  OR3_X1    g334(.A1(new_n520), .A2(KEYINPUT85), .A3(G125), .ZN(new_n521));
  OAI21_X1  g335(.A(KEYINPUT85), .B1(new_n520), .B2(G125), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n521), .B(new_n522), .C1(new_n332), .C2(new_n247), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n312), .A2(G224), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(KEYINPUT86), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n523), .B(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n416), .A2(KEYINPUT79), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT79), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(G104), .ZN(new_n529));
  INV_X1    g343(.A(G107), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT3), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT3), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT80), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(G107), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n530), .A2(KEYINPUT80), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n533), .B(G104), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n527), .A2(new_n529), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(G107), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n532), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(G101), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n532), .A2(new_n537), .A3(new_n539), .A4(new_n266), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(KEYINPUT4), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT4), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n540), .A2(new_n544), .A3(G101), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n543), .A2(new_n203), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT5), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n547), .B(G116), .C1(new_n342), .C2(new_n343), .ZN(new_n548));
  OAI211_X1 g362(.A(G113), .B(new_n548), .C1(new_n199), .C2(new_n547), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n198), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n531), .B1(new_n449), .B2(G104), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(G101), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n542), .ZN(new_n553));
  OR2_X1    g367(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n546), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT6), .ZN(new_n556));
  XOR2_X1   g370(.A(G110), .B(G122), .Z(new_n557));
  NAND3_X1  g371(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n555), .A2(new_n557), .ZN(new_n559));
  INV_X1    g373(.A(new_n557), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n546), .A2(new_n554), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n559), .A2(KEYINPUT6), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n526), .A2(new_n558), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT7), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n525), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n523), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n550), .B(new_n553), .ZN(new_n567));
  XOR2_X1   g381(.A(new_n557), .B(KEYINPUT8), .Z(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n561), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n563), .A2(new_n570), .A3(new_n364), .ZN(new_n571));
  OAI21_X1  g385(.A(G210), .B1(G237), .B2(G902), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n572), .B(KEYINPUT88), .Z(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(KEYINPUT87), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n571), .A2(new_n575), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n515), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(G221), .B1(new_n486), .B2(G902), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT84), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n543), .A2(new_n247), .A3(new_n545), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT81), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n224), .B1(new_n232), .B2(KEYINPUT1), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n516), .B1(new_n246), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n586), .A2(new_n542), .A3(new_n552), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT10), .ZN(new_n588));
  INV_X1    g402(.A(new_n553), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n588), .B1(new_n516), .B2(new_n519), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n587), .A2(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n543), .A2(KEYINPUT81), .A3(new_n247), .A4(new_n545), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n584), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n593), .A2(new_n241), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n241), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT83), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n593), .A2(KEYINPUT83), .A3(new_n241), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n594), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n312), .A2(G227), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(KEYINPUT78), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(new_n345), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(new_n330), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n581), .B1(new_n599), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n553), .A2(new_n519), .A3(new_n516), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n587), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n241), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT12), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT82), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT82), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n608), .A2(new_n612), .A3(new_n609), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n611), .B(new_n613), .C1(new_n609), .C2(new_n608), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n594), .A2(new_n603), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n594), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n593), .A2(KEYINPUT83), .A3(new_n241), .ZN(new_n618));
  AOI21_X1  g432(.A(KEYINPUT83), .B1(new_n593), .B2(new_n241), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n620), .A2(KEYINPUT84), .A3(new_n603), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n605), .A2(new_n616), .A3(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(G469), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n622), .A2(new_n623), .A3(new_n364), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n604), .B1(new_n614), .B2(new_n617), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n597), .A2(new_n598), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n625), .B1(new_n615), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(G469), .B1(new_n627), .B2(G902), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n580), .B1(new_n624), .B2(new_n628), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n513), .A2(new_n578), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n311), .A2(KEYINPUT77), .A3(new_n381), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n383), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G101), .ZN(G3));
  OAI21_X1  g447(.A(new_n364), .B1(new_n294), .B2(new_n285), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(G472), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n307), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n629), .A2(new_n381), .A3(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT33), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n639), .B1(new_n488), .B2(new_n489), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n504), .A2(KEYINPUT33), .A3(new_n505), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n640), .A2(new_n641), .A3(G478), .A4(new_n364), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n490), .A2(new_n491), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(new_n445), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n571), .A2(new_n574), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n563), .A2(new_n570), .A3(new_n364), .A4(new_n573), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n648), .A2(new_n514), .A3(new_n392), .A4(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n638), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(new_n416), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT102), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT34), .ZN(G6));
  INV_X1    g469(.A(new_n440), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT20), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n659), .B1(new_n440), .B2(KEYINPUT20), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n656), .A2(new_n659), .A3(new_n657), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR4_X1   g477(.A1(new_n663), .A2(new_n650), .A3(new_n511), .A4(new_n421), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n638), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT35), .B(G107), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G9));
  NAND4_X1  g481(.A1(new_n513), .A2(new_n578), .A3(new_n629), .A4(new_n637), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n359), .A2(KEYINPUT36), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n370), .B(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n378), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n377), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n668), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT37), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G110), .ZN(G12));
  NAND3_X1  g490(.A1(new_n648), .A2(new_n514), .A3(new_n649), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n673), .ZN(new_n678));
  INV_X1    g492(.A(new_n421), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n391), .A2(G900), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n389), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n663), .A2(new_n511), .A3(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n311), .A2(new_n629), .A3(new_n678), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G128), .ZN(G30));
  XOR2_X1   g499(.A(new_n681), .B(KEYINPUT39), .Z(new_n686));
  AOI211_X1 g500(.A(new_n580), .B(new_n686), .C1(new_n624), .C2(new_n628), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT40), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n441), .A2(new_n444), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n679), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n509), .A3(new_n510), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n576), .A2(new_n577), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n694), .B(KEYINPUT38), .Z(new_n695));
  AOI21_X1  g509(.A(new_n695), .B1(new_n687), .B2(new_n688), .ZN(new_n696));
  AOI22_X1  g510(.A1(new_n291), .A2(new_n293), .B1(new_n275), .B2(new_n297), .ZN(new_n697));
  OAI21_X1  g511(.A(G472), .B1(new_n697), .B2(G902), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n289), .A2(new_n295), .A3(new_n310), .A4(new_n698), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n699), .A2(new_n673), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n693), .A2(new_n514), .A3(new_n696), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n466), .ZN(G45));
  NAND3_X1  g516(.A1(new_n691), .A2(new_n644), .A3(new_n681), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n677), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n311), .A2(new_n629), .A3(new_n672), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  AND3_X1   g520(.A1(new_n622), .A2(new_n623), .A3(new_n364), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n623), .B1(new_n622), .B2(new_n364), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n707), .A2(new_n708), .A3(new_n580), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n709), .A2(new_n311), .A3(new_n381), .A4(new_n651), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT104), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT41), .B(G113), .Z(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G15));
  NAND4_X1  g527(.A1(new_n709), .A2(new_n664), .A3(new_n311), .A4(new_n381), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G116), .ZN(G18));
  NAND4_X1  g529(.A1(new_n709), .A2(new_n311), .A3(new_n513), .A4(new_n678), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  NOR4_X1   g531(.A1(new_n707), .A2(new_n708), .A3(new_n692), .A4(new_n580), .ZN(new_n718));
  INV_X1    g532(.A(new_n272), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n290), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n298), .A2(new_n267), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n274), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n187), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT105), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n377), .A2(new_n380), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n724), .B1(new_n377), .B2(new_n380), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n723), .A2(new_n635), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT106), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n723), .A2(new_n635), .A3(new_n727), .A4(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n650), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n718), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G122), .ZN(G24));
  NOR2_X1   g549(.A1(new_n707), .A2(new_n708), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n723), .A2(new_n635), .A3(new_n672), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n736), .A2(new_n579), .A3(new_n737), .A4(new_n704), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  NAND2_X1  g553(.A1(new_n311), .A2(new_n381), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n703), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n576), .A2(new_n577), .A3(new_n514), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n629), .A2(KEYINPUT107), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT107), .B1(new_n629), .B2(new_n744), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n741), .B(new_n742), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT42), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n624), .A2(new_n628), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n579), .A3(new_n744), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT107), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n629), .A2(KEYINPUT107), .A3(new_n744), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n703), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g568(.A(KEYINPUT108), .B1(new_n287), .B2(KEYINPUT32), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT32), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n307), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n755), .A2(new_n306), .A3(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(KEYINPUT42), .A3(new_n727), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  AOI22_X1  g575(.A1(new_n747), .A2(new_n748), .B1(new_n754), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(new_n213), .ZN(G33));
  OAI211_X1 g577(.A(new_n741), .B(new_n683), .C1(new_n745), .C2(new_n746), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G134), .ZN(G36));
  NAND2_X1  g579(.A1(new_n445), .A2(new_n644), .ZN(new_n766));
  NAND2_X1  g580(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g582(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n769));
  OAI21_X1  g583(.A(new_n768), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n636), .A3(new_n672), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT44), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT110), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n627), .A2(KEYINPUT45), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n626), .A2(new_n615), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n776), .B1(new_n777), .B2(new_n625), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n775), .A2(new_n778), .A3(G469), .ZN(new_n779));
  NAND2_X1  g593(.A1(G469), .A2(G902), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT46), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n779), .A2(KEYINPUT46), .A3(new_n780), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(new_n784), .A3(new_n624), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n579), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n686), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n743), .B1(new_n771), .B2(new_n772), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n774), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G137), .ZN(G39));
  NAND2_X1  g604(.A1(new_n786), .A2(KEYINPUT47), .ZN(new_n791));
  INV_X1    g605(.A(new_n311), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n743), .A2(new_n703), .A3(new_n381), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT47), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n785), .A2(new_n794), .A3(new_n579), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n791), .A2(new_n792), .A3(new_n793), .A4(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G140), .ZN(G42));
  NAND2_X1  g611(.A1(new_n791), .A2(new_n795), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n736), .B(KEYINPUT111), .Z(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n580), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n743), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n389), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n770), .A2(new_n802), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n803), .A2(new_n732), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n804), .A2(new_n515), .A3(new_n695), .A4(new_n709), .ZN(new_n806));
  XOR2_X1   g620(.A(new_n806), .B(KEYINPUT50), .Z(new_n807));
  AND3_X1   g621(.A1(new_n803), .A2(new_n709), .A3(new_n744), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n737), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n709), .A2(new_n381), .A3(new_n744), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n810), .A2(new_n389), .A3(new_n699), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n691), .A2(new_n644), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n805), .A2(new_n807), .A3(new_n809), .A4(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n801), .A2(new_n804), .B1(new_n811), .B2(new_n812), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n817), .A2(KEYINPUT51), .A3(new_n809), .A4(new_n807), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n804), .A2(new_n709), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n677), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(KEYINPUT119), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n759), .A2(new_n727), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n808), .A2(new_n822), .ZN(new_n823));
  XOR2_X1   g637(.A(new_n823), .B(KEYINPUT48), .Z(new_n824));
  NAND2_X1  g638(.A1(new_n811), .A2(new_n646), .ZN(new_n825));
  INV_X1    g639(.A(new_n387), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n825), .B1(KEYINPUT118), .B2(new_n826), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n821), .A2(new_n824), .A3(new_n827), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n816), .A2(new_n818), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n826), .A2(KEYINPUT118), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n742), .B(new_n737), .C1(new_n745), .C2(new_n746), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n493), .A2(new_n495), .ZN(new_n832));
  NOR4_X1   g646(.A1(new_n743), .A2(new_n663), .A3(new_n832), .A4(new_n682), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n833), .A2(new_n311), .A3(new_n629), .A4(new_n672), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n764), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n762), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n630), .A2(new_n637), .A3(new_n672), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n646), .A2(KEYINPUT112), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n445), .A2(new_n832), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n646), .A2(KEYINPUT112), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n638), .A2(new_n578), .A3(new_n392), .A4(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n632), .A2(new_n837), .A3(new_n842), .A4(new_n716), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n734), .A2(new_n710), .A3(new_n714), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT114), .B1(new_n389), .B2(new_n680), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n692), .A2(new_n677), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n699), .A2(new_n673), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT114), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n629), .B1(new_n849), .B2(new_n681), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n705), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n738), .A2(new_n684), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT52), .ZN(new_n853));
  OR3_X1    g667(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n853), .B1(new_n851), .B2(new_n852), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n836), .A2(new_n845), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT116), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n855), .A2(KEYINPUT115), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT115), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n861), .B(new_n853), .C1(new_n851), .C2(new_n852), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n705), .B(KEYINPUT52), .C1(new_n848), .C2(new_n850), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT113), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n738), .A2(new_n684), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n852), .A2(KEYINPUT113), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n864), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n860), .A2(new_n862), .A3(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n836), .A2(new_n845), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n858), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n834), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n740), .B1(new_n752), .B2(new_n753), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n873), .B1(new_n874), .B2(new_n683), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT42), .B1(new_n874), .B2(new_n742), .ZN(new_n876));
  AOI211_X1 g690(.A(new_n703), .B(new_n760), .C1(new_n752), .C2(new_n753), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n831), .B(new_n875), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n311), .A2(KEYINPUT77), .A3(new_n381), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(new_n382), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n674), .B1(new_n880), .B2(new_n630), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n734), .A2(new_n710), .A3(new_n714), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n881), .A2(new_n882), .A3(new_n716), .A4(new_n842), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT116), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n884), .A2(new_n885), .A3(KEYINPUT53), .A4(new_n856), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n859), .A2(new_n872), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT54), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n869), .A2(KEYINPUT53), .A3(new_n836), .A4(new_n845), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT117), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n884), .A2(KEYINPUT117), .A3(KEYINPUT53), .A4(new_n869), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n857), .A2(new_n858), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n891), .A2(new_n892), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n829), .A2(new_n830), .A3(new_n888), .A4(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n896), .B1(G952), .B2(G953), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n799), .B(KEYINPUT49), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n695), .A2(new_n727), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n899), .A2(new_n699), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n766), .A2(new_n515), .A3(new_n580), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n898), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n897), .A2(new_n902), .ZN(G75));
  NAND3_X1  g717(.A1(new_n891), .A2(new_n892), .A3(new_n894), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n904), .A2(G902), .A3(new_n573), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT56), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n562), .A2(new_n558), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(new_n526), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT55), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n905), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n909), .B1(new_n905), .B2(new_n906), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n312), .A2(G952), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(G51));
  NAND2_X1  g727(.A1(new_n904), .A2(KEYINPUT54), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n895), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n780), .B(KEYINPUT57), .Z(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n622), .ZN(new_n918));
  INV_X1    g732(.A(new_n779), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n904), .A2(G902), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n912), .B1(new_n918), .B2(new_n920), .ZN(G54));
  AND2_X1   g735(.A1(KEYINPUT58), .A2(G475), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n904), .A2(G902), .A3(new_n922), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n434), .A2(new_n437), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  OR3_X1    g739(.A1(new_n923), .A2(KEYINPUT120), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n912), .B1(new_n923), .B2(new_n925), .ZN(new_n927));
  OAI21_X1  g741(.A(KEYINPUT120), .B1(new_n923), .B2(new_n925), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(G60));
  INV_X1    g743(.A(new_n912), .ZN(new_n930));
  NAND2_X1  g744(.A1(G478), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT59), .Z(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n888), .B2(new_n895), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n640), .A2(new_n641), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n932), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n915), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n935), .A2(new_n937), .ZN(G63));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT60), .Z(new_n940));
  NAND2_X1  g754(.A1(new_n904), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n361), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n904), .A2(new_n670), .A3(new_n940), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n943), .A2(new_n930), .A3(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT61), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n943), .A2(KEYINPUT61), .A3(new_n930), .A4(new_n944), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(G66));
  AOI21_X1  g763(.A(new_n312), .B1(new_n390), .B2(G224), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n883), .B(KEYINPUT121), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n950), .B1(new_n951), .B2(new_n312), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n907), .B1(G898), .B2(new_n312), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT122), .Z(new_n954));
  XNOR2_X1  g768(.A(new_n952), .B(new_n954), .ZN(G69));
  NAND2_X1  g769(.A1(new_n789), .A2(new_n796), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n867), .A2(new_n866), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n957), .A2(new_n701), .A3(new_n705), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n957), .A2(KEYINPUT62), .A3(new_n701), .A4(new_n705), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n956), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n880), .A2(new_n687), .A3(new_n744), .A4(new_n841), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT124), .Z(new_n964));
  AOI21_X1  g778(.A(G953), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT125), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n270), .B(KEYINPUT123), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(new_n428), .Z(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  OR3_X1    g783(.A1(new_n965), .A2(new_n966), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(G900), .A2(G953), .ZN(new_n971));
  INV_X1    g785(.A(new_n956), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n957), .A2(new_n705), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n973), .A2(new_n762), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n692), .A2(new_n677), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n787), .A2(new_n822), .A3(new_n975), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n972), .A2(new_n764), .A3(new_n974), .A4(new_n976), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n969), .B(new_n971), .C1(new_n977), .C2(G953), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n966), .B1(new_n965), .B2(new_n969), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n970), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(G227), .A2(G900), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(G953), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT126), .Z(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n970), .A2(new_n979), .A3(new_n983), .A4(new_n978), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(G72));
  NAND2_X1  g801(.A1(G472), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT63), .Z(new_n989));
  NAND2_X1  g803(.A1(new_n962), .A2(new_n964), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n989), .B1(new_n990), .B2(new_n951), .ZN(new_n991));
  INV_X1    g805(.A(new_n261), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n991), .A2(new_n992), .A3(new_n267), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n989), .B1(new_n977), .B2(new_n951), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n994), .A2(new_n261), .A3(new_n275), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n993), .A2(new_n930), .A3(new_n995), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n268), .A2(new_n273), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n261), .A2(new_n267), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n989), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT127), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n996), .B1(new_n887), .B2(new_n1000), .ZN(G57));
endmodule


