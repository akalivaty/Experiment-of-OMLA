//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 0 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G210), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n190), .B(KEYINPUT27), .Z(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(G101), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G116), .ZN(new_n194));
  OR3_X1    g008(.A1(new_n194), .A2(KEYINPUT69), .A3(G119), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT69), .B1(new_n194), .B2(G119), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(G119), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  XOR2_X1   g012(.A(KEYINPUT2), .B(G113), .Z(new_n199));
  XNOR2_X1  g013(.A(new_n198), .B(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT30), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(KEYINPUT68), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(KEYINPUT68), .ZN(new_n204));
  AND2_X1   g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  AOI21_X1  g025(.A(G146), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n213), .B1(new_n214), .B2(G143), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n208), .A2(KEYINPUT65), .A3(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n207), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n208), .A2(G146), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n209), .A2(new_n211), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n220), .B(new_n205), .C1(new_n221), .C2(new_n214), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n223));
  INV_X1    g037(.A(G137), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AND2_X1   g039(.A1(KEYINPUT11), .A2(G134), .ZN(new_n226));
  NAND2_X1  g040(.A1(KEYINPUT66), .A2(G137), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G131), .ZN(new_n229));
  NAND2_X1  g043(.A1(KEYINPUT11), .A2(G134), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT11), .A2(G134), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(G137), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n228), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n229), .B1(new_n228), .B2(new_n232), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n218), .B(new_n222), .C1(new_n233), .C2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n228), .A2(new_n232), .A3(new_n229), .ZN(new_n237));
  INV_X1    g051(.A(G134), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n225), .A2(new_n238), .A3(new_n227), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n229), .B1(G134), .B2(G137), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G128), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n243), .A2(KEYINPUT1), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n220), .B(new_n244), .C1(new_n221), .C2(new_n214), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT67), .B(G128), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT1), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n247), .B1(G143), .B2(new_n214), .ZN(new_n248));
  OAI22_X1  g062(.A1(new_n212), .A2(new_n217), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n242), .B1(new_n245), .B2(new_n249), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n203), .B(new_n204), .C1(new_n236), .C2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n245), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n237), .A2(new_n241), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n254), .A2(KEYINPUT68), .A3(new_n201), .A4(new_n235), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n200), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n254), .A2(new_n200), .A3(new_n235), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT70), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n254), .A2(KEYINPUT70), .A3(new_n200), .A4(new_n235), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n193), .B1(new_n256), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n200), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n263), .B1(new_n236), .B2(new_n250), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n259), .A2(new_n260), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT28), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT28), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n257), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n193), .B(KEYINPUT71), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT29), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n262), .B1(new_n269), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n268), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n275), .B1(new_n265), .B2(KEYINPUT28), .ZN(new_n276));
  INV_X1    g090(.A(new_n193), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n272), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n187), .B1(new_n274), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G472), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n269), .A2(new_n270), .ZN(new_n281));
  INV_X1    g095(.A(new_n261), .ZN(new_n282));
  INV_X1    g096(.A(new_n204), .ZN(new_n283));
  AOI211_X1 g097(.A(new_n202), .B(new_n283), .C1(new_n254), .C2(new_n235), .ZN(new_n284));
  INV_X1    g098(.A(new_n255), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n263), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n282), .A2(new_n286), .A3(new_n277), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT31), .ZN(new_n288));
  NOR3_X1   g102(.A1(new_n256), .A2(new_n261), .A3(new_n193), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT31), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n281), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G472), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n292), .A2(KEYINPUT32), .A3(new_n293), .A4(new_n187), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n280), .A2(new_n294), .ZN(new_n295));
  OAI22_X1  g109(.A1(new_n289), .A2(new_n290), .B1(new_n276), .B2(new_n271), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n287), .A2(KEYINPUT31), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n293), .B(new_n187), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  XOR2_X1   g112(.A(KEYINPUT72), .B(KEYINPUT32), .Z(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT73), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n298), .A2(KEYINPUT73), .A3(new_n299), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n295), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G119), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G128), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n306), .B(KEYINPUT75), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n246), .A2(G119), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  XOR2_X1   g123(.A(KEYINPUT24), .B(G110), .Z(new_n310));
  NAND3_X1  g124(.A1(new_n246), .A2(KEYINPUT23), .A3(G119), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n305), .A2(G128), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n311), .B(new_n306), .C1(KEYINPUT23), .C2(new_n312), .ZN(new_n313));
  OAI22_X1  g127(.A1(new_n309), .A2(new_n310), .B1(new_n313), .B2(G110), .ZN(new_n314));
  XNOR2_X1  g128(.A(G125), .B(G140), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT16), .ZN(new_n316));
  INV_X1    g130(.A(G140), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G125), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n316), .B(G146), .C1(KEYINPUT16), .C2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n315), .A2(new_n214), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n314), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n316), .B1(KEYINPUT16), .B2(new_n318), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n214), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(new_n319), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n313), .A2(G110), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n309), .A2(new_n310), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n321), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT22), .B(G137), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n329), .B(new_n330), .ZN(new_n331));
  XOR2_X1   g145(.A(new_n331), .B(KEYINPUT76), .Z(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n321), .A2(new_n327), .A3(new_n331), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n187), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT25), .ZN(new_n337));
  NAND2_X1  g151(.A1(G217), .A2(G902), .ZN(new_n338));
  INV_X1    g152(.A(G217), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n338), .B1(new_n339), .B2(G234), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n340), .B(KEYINPUT74), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT25), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n334), .A2(new_n342), .A3(new_n187), .A4(new_n335), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n337), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n334), .A2(new_n335), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n341), .A2(G902), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT77), .B1(new_n304), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT77), .ZN(new_n350));
  INV_X1    g164(.A(new_n348), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n298), .A2(KEYINPUT73), .A3(new_n299), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT73), .B1(new_n298), .B2(new_n299), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n350), .B(new_n351), .C1(new_n354), .C2(new_n295), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n349), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT9), .B(G234), .ZN(new_n357));
  OAI21_X1  g171(.A(G221), .B1(new_n357), .B2(G902), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G107), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G104), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(KEYINPUT78), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT78), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G107), .ZN(new_n364));
  AOI21_X1  g178(.A(G104), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT80), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n361), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(KEYINPUT78), .B(G107), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n368), .A2(KEYINPUT80), .A3(G104), .ZN(new_n369));
  OAI21_X1  g183(.A(G101), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(KEYINPUT81), .ZN(new_n371));
  INV_X1    g185(.A(new_n212), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n243), .B1(new_n372), .B2(KEYINPUT1), .ZN(new_n373));
  INV_X1    g187(.A(new_n221), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n219), .B1(new_n374), .B2(G146), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n245), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G104), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(KEYINPUT3), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n379), .B1(new_n360), .B2(G104), .ZN(new_n380));
  AOI22_X1  g194(.A1(new_n368), .A2(new_n378), .B1(new_n380), .B2(new_n361), .ZN(new_n381));
  INV_X1    g195(.A(G101), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT81), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n384), .B(G101), .C1(new_n367), .C2(new_n369), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n371), .A2(new_n376), .A3(new_n383), .A4(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT10), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n233), .A2(new_n234), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n218), .A2(new_n222), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT4), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n378), .A2(new_n362), .A3(new_n364), .ZN(new_n393));
  AOI21_X1  g207(.A(KEYINPUT3), .B1(new_n377), .B2(G107), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n377), .A2(G107), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT79), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n380), .A2(new_n361), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n378), .A2(new_n362), .A3(new_n364), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT79), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n397), .A2(G101), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n392), .B1(new_n402), .B2(new_n383), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n398), .A2(new_n399), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n382), .B1(new_n404), .B2(KEYINPUT79), .ZN(new_n405));
  AOI21_X1  g219(.A(KEYINPUT4), .B1(new_n405), .B2(new_n401), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n391), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n387), .B1(new_n249), .B2(new_n245), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n371), .A2(new_n383), .A3(new_n385), .A4(new_n408), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n388), .A2(new_n389), .A3(new_n407), .A4(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(G110), .B(G140), .ZN(new_n411));
  INV_X1    g225(.A(G227), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(G953), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n411), .B(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n252), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n385), .A2(new_n383), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n365), .A2(new_n366), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT80), .B1(new_n368), .B2(G104), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(new_n361), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n384), .B1(new_n420), .B2(G101), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n416), .B1(new_n417), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n386), .ZN(new_n423));
  INV_X1    g237(.A(new_n389), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT12), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT12), .ZN(new_n426));
  AOI211_X1 g240(.A(new_n426), .B(new_n389), .C1(new_n422), .C2(new_n386), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n410), .B(new_n415), .C1(new_n425), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(KEYINPUT82), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n423), .A2(new_n424), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n426), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n423), .A2(KEYINPUT12), .A3(new_n424), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n410), .A2(new_n415), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT82), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n407), .A2(new_n409), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n417), .A2(new_n421), .ZN(new_n438));
  AOI21_X1  g252(.A(KEYINPUT10), .B1(new_n438), .B2(new_n376), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n424), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n410), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n414), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n429), .A2(new_n436), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G469), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(new_n444), .A3(new_n187), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n444), .A2(new_n187), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n410), .B1(new_n425), .B2(new_n427), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n447), .A2(new_n414), .B1(new_n434), .B2(new_n440), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n446), .B1(new_n448), .B2(G469), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n359), .B1(new_n445), .B2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(G110), .B(G122), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(G101), .B1(new_n381), .B2(new_n400), .ZN(new_n453));
  INV_X1    g267(.A(new_n401), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n383), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT4), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n392), .B1(new_n453), .B2(new_n454), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n200), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT5), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(new_n305), .A3(G116), .ZN(new_n460));
  OAI211_X1 g274(.A(G113), .B(new_n460), .C1(new_n198), .C2(new_n459), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n199), .A2(new_n196), .A3(new_n195), .A4(new_n197), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR3_X1   g277(.A1(new_n417), .A2(new_n421), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n452), .B1(new_n458), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n464), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n404), .A2(G101), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n467), .B1(new_n405), .B2(new_n401), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n457), .B1(new_n468), .B2(new_n392), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n263), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n466), .A2(new_n470), .A3(new_n451), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n465), .A2(new_n471), .A3(KEYINPUT6), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT6), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n473), .B(new_n452), .C1(new_n458), .C2(new_n464), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n390), .A2(G125), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n252), .A2(G125), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n189), .A2(G224), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n478), .B(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n472), .A2(new_n474), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(KEYINPUT7), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n482), .B1(new_n476), .B2(new_n477), .ZN(new_n483));
  INV_X1    g297(.A(new_n482), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n475), .B(new_n484), .C1(G125), .C2(new_n252), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n463), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n438), .A2(new_n487), .B1(new_n469), .B2(new_n263), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n486), .B1(new_n488), .B2(new_n451), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n451), .B(KEYINPUT8), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n438), .A2(new_n487), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n490), .B1(new_n491), .B2(new_n464), .ZN(new_n492));
  AOI21_X1  g306(.A(G902), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(G210), .B1(G237), .B2(G902), .ZN(new_n494));
  OR2_X1    g308(.A1(new_n494), .A2(KEYINPUT83), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n481), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n495), .B1(new_n481), .B2(new_n493), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(G214), .B1(G237), .B2(G902), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n324), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT87), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n188), .A2(new_n189), .A3(G143), .A4(G214), .ZN(new_n504));
  INV_X1    g318(.A(G214), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n505), .A2(G237), .A3(G953), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n504), .B1(new_n221), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n503), .B1(new_n507), .B2(G131), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n209), .A3(new_n211), .ZN(new_n510));
  AOI211_X1 g324(.A(KEYINPUT87), .B(new_n229), .C1(new_n510), .C2(new_n504), .ZN(new_n511));
  OAI21_X1  g325(.A(KEYINPUT17), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n507), .A2(G131), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT87), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n507), .A2(new_n503), .A3(G131), .ZN(new_n515));
  OAI21_X1  g329(.A(KEYINPUT86), .B1(new_n507), .B2(G131), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT86), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n510), .A2(new_n517), .A3(new_n229), .A4(new_n504), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n514), .A2(new_n515), .A3(new_n516), .A4(new_n518), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n502), .B(new_n512), .C1(new_n519), .C2(KEYINPUT17), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT85), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n320), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(G125), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G140), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n318), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT84), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n315), .A2(KEYINPUT84), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n522), .B1(new_n529), .B2(G146), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n507), .A2(KEYINPUT18), .A3(G131), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n527), .A2(new_n528), .A3(KEYINPUT85), .A4(G146), .ZN(new_n532));
  NAND2_X1  g346(.A1(KEYINPUT18), .A2(G131), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n510), .A2(new_n533), .A3(new_n504), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(G113), .B(G122), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(new_n377), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n520), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n539), .B1(new_n520), .B2(new_n537), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n187), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G475), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT20), .ZN(new_n544));
  NOR2_X1   g358(.A1(G475), .A2(G902), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n519), .A2(KEYINPUT88), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n508), .A2(new_n511), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT88), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n547), .A2(new_n548), .A3(new_n516), .A4(new_n518), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n527), .A2(new_n528), .A3(KEYINPUT19), .ZN(new_n550));
  OR2_X1    g364(.A1(new_n525), .A2(KEYINPUT19), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n550), .A2(new_n214), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n319), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n546), .A2(new_n549), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n539), .B1(new_n555), .B2(new_n537), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n544), .B(new_n545), .C1(new_n556), .C2(new_n540), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n520), .A2(new_n537), .A3(new_n539), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n553), .B1(new_n519), .B2(KEYINPUT88), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n536), .B1(new_n560), .B2(new_n549), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n559), .B1(new_n561), .B2(new_n539), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n544), .B1(new_n562), .B2(new_n545), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n543), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(KEYINPUT91), .A2(G952), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(KEYINPUT91), .A2(G952), .ZN(new_n567));
  AOI21_X1  g381(.A(G953), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(G234), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n568), .B1(new_n569), .B2(new_n188), .ZN(new_n570));
  AOI211_X1 g384(.A(new_n187), .B(new_n189), .C1(G234), .C2(G237), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT21), .B(G898), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n357), .A2(new_n339), .A3(G953), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n209), .A2(new_n211), .A3(G128), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n243), .A2(KEYINPUT67), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT67), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(G128), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n578), .A2(new_n580), .A3(G143), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n577), .A2(new_n581), .A3(new_n238), .ZN(new_n582));
  XNOR2_X1  g396(.A(G116), .B(G122), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n368), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n368), .A2(new_n583), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n582), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n209), .A2(new_n211), .A3(KEYINPUT13), .A4(G128), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n588), .A2(new_n581), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT13), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n577), .A2(KEYINPUT89), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(KEYINPUT89), .B1(new_n577), .B2(new_n590), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n587), .B1(new_n593), .B2(G134), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n194), .A2(G122), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n360), .B1(new_n595), .B2(KEYINPUT14), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT14), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n583), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n584), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n577), .A2(new_n581), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(G134), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n600), .B1(new_n582), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n576), .B1(new_n594), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n582), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n605), .A2(new_n584), .A3(new_n599), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n577), .A2(new_n590), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT89), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n577), .A2(KEYINPUT89), .A3(new_n590), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n238), .B1(new_n611), .B2(new_n589), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n606), .B(new_n575), .C1(new_n612), .C2(new_n587), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n604), .A2(new_n613), .A3(KEYINPUT90), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT90), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n615), .B(new_n576), .C1(new_n594), .C2(new_n603), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n187), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(G478), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(KEYINPUT15), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n617), .B(new_n619), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n564), .A2(new_n574), .A3(new_n620), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n450), .A2(new_n501), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n356), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G101), .ZN(G3));
  OAI21_X1  g438(.A(new_n187), .B1(new_n296), .B2(new_n297), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT92), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n625), .A2(new_n626), .A3(G472), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(G472), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n292), .A2(new_n187), .A3(new_n628), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n627), .A2(new_n351), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n450), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT93), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n481), .A2(new_n493), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n500), .B1(new_n633), .B2(new_n494), .ZN(new_n634));
  INV_X1    g448(.A(new_n574), .ZN(new_n635));
  INV_X1    g449(.A(new_n494), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n481), .A2(new_n493), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n634), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(G475), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n520), .A2(new_n537), .ZN(new_n640));
  INV_X1    g454(.A(new_n539), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n559), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n639), .B1(new_n643), .B2(new_n187), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n562), .A2(new_n545), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(KEYINPUT20), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n644), .B1(new_n646), .B2(new_n557), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT33), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n614), .A2(new_n648), .A3(new_n616), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n604), .A2(new_n613), .A3(KEYINPUT33), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n618), .A2(G902), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  AND3_X1   g466(.A1(new_n617), .A2(KEYINPUT94), .A3(new_n618), .ZN(new_n653));
  AOI21_X1  g467(.A(KEYINPUT94), .B1(new_n617), .B2(new_n618), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n638), .A2(new_n647), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n632), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT95), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT34), .B(G104), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G6));
  INV_X1    g475(.A(KEYINPUT97), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n557), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n562), .A2(KEYINPUT97), .A3(new_n544), .A4(new_n545), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n646), .A2(KEYINPUT96), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n663), .A2(new_n646), .A3(KEYINPUT96), .A4(new_n664), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n669), .A2(new_n543), .A3(new_n620), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n638), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n632), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT35), .B(G107), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G9));
  NAND2_X1  g488(.A1(new_n627), .A2(new_n629), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT98), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n676), .B1(new_n321), .B2(new_n327), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n333), .A2(KEYINPUT36), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n321), .A2(new_n676), .A3(new_n327), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n679), .B1(new_n678), .B2(new_n680), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n346), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n344), .ZN(new_n684));
  INV_X1    g498(.A(new_n620), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n647), .A2(new_n635), .A3(new_n684), .A4(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n675), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n687), .A2(new_n450), .A3(new_n501), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT99), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT37), .B(G110), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G12));
  NAND2_X1  g505(.A1(new_n445), .A2(new_n449), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n358), .ZN(new_n693));
  OR2_X1    g507(.A1(KEYINPUT100), .A2(G900), .ZN(new_n694));
  NAND2_X1  g508(.A1(KEYINPUT100), .A2(G900), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n571), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n570), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT101), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n669), .A2(new_n543), .A3(new_n620), .A4(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n693), .A2(new_n700), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n481), .A2(new_n493), .A3(new_n636), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n636), .B1(new_n481), .B2(new_n493), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n702), .A2(new_n703), .A3(new_n500), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n684), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n302), .A2(new_n303), .ZN(new_n706));
  INV_X1    g520(.A(new_n295), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n701), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G128), .ZN(G30));
  XNOR2_X1  g524(.A(new_n698), .B(KEYINPUT39), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n693), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT104), .ZN(new_n713));
  OR2_X1    g527(.A1(new_n713), .A2(KEYINPUT40), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(KEYINPUT40), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n265), .A2(new_n270), .ZN(new_n716));
  OAI21_X1  g530(.A(KEYINPUT102), .B1(new_n289), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n187), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n289), .A2(new_n716), .A3(KEYINPUT102), .ZN(new_n719));
  OAI21_X1  g533(.A(G472), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n720), .A2(new_n294), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n706), .A2(KEYINPUT103), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(KEYINPUT103), .B1(new_n706), .B2(new_n721), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OR2_X1    g538(.A1(new_n498), .A2(KEYINPUT38), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n498), .A2(KEYINPUT38), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n564), .A2(new_n620), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n683), .A2(new_n344), .A3(new_n499), .ZN(new_n729));
  NOR4_X1   g543(.A1(new_n724), .A2(new_n727), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n714), .A2(new_n715), .A3(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(new_n221), .ZN(G45));
  INV_X1    g546(.A(KEYINPUT105), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n634), .A2(new_n637), .A3(new_n684), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n734), .B1(new_n354), .B2(new_n295), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n564), .A2(new_n655), .A3(new_n699), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n450), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n733), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n450), .A2(new_n736), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n708), .A2(new_n739), .A3(KEYINPUT105), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G146), .ZN(G48));
  AOI21_X1  g556(.A(new_n348), .B1(new_n706), .B2(new_n707), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n443), .A2(new_n187), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(G469), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n358), .A3(new_n445), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT106), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n745), .A2(KEYINPUT106), .A3(new_n358), .A4(new_n445), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n743), .A2(new_n748), .A3(new_n749), .A4(new_n657), .ZN(new_n750));
  XNOR2_X1  g564(.A(KEYINPUT41), .B(G113), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n750), .B(new_n751), .ZN(G15));
  NAND4_X1  g566(.A1(new_n743), .A2(new_n748), .A3(new_n671), .A4(new_n749), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G116), .ZN(G18));
  NAND4_X1  g568(.A1(new_n745), .A2(new_n704), .A3(new_n358), .A4(new_n445), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n304), .A2(new_n755), .A3(new_n686), .ZN(new_n756));
  XOR2_X1   g570(.A(KEYINPUT107), .B(G119), .Z(new_n757));
  XNOR2_X1  g571(.A(new_n756), .B(new_n757), .ZN(G21));
  INV_X1    g572(.A(new_n704), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n625), .A2(G472), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n760), .A2(new_n298), .A3(new_n351), .A4(new_n635), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n759), .A2(new_n761), .A3(new_n728), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n748), .A2(new_n762), .A3(new_n749), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G122), .ZN(G24));
  NAND4_X1  g578(.A1(new_n736), .A2(new_n298), .A3(new_n684), .A4(new_n760), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n755), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(new_n523), .ZN(G27));
  NOR3_X1   g581(.A1(new_n496), .A2(new_n497), .A3(new_n500), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n692), .A2(new_n358), .A3(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT32), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n298), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n348), .B1(new_n707), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n564), .A2(new_n655), .A3(new_n699), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT42), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n769), .A2(new_n772), .A3(new_n775), .ZN(new_n776));
  AOI22_X1  g590(.A1(new_n428), .A2(KEYINPUT82), .B1(new_n441), .B2(new_n414), .ZN(new_n777));
  AOI211_X1 g591(.A(G469), .B(G902), .C1(new_n777), .C2(new_n436), .ZN(new_n778));
  INV_X1    g592(.A(new_n449), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n768), .B(new_n358), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n304), .A2(new_n780), .A3(new_n348), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT108), .B1(new_n781), .B2(new_n736), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n743), .A2(KEYINPUT108), .A3(new_n736), .A4(new_n769), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n774), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n776), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G131), .ZN(G33));
  INV_X1    g600(.A(new_n700), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n743), .A2(new_n787), .A3(new_n769), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G134), .ZN(G36));
  NAND2_X1  g603(.A1(new_n647), .A2(new_n655), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT43), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n675), .A3(new_n684), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT44), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n768), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n796), .A2(KEYINPUT109), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(KEYINPUT109), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n795), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT46), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n448), .A2(KEYINPUT45), .ZN(new_n801));
  OAI21_X1  g615(.A(G469), .B1(new_n448), .B2(KEYINPUT45), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n800), .B1(new_n803), .B2(new_n446), .ZN(new_n804));
  OAI221_X1 g618(.A(KEYINPUT46), .B1(new_n444), .B2(new_n187), .C1(new_n802), .C2(new_n801), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n445), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n358), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(new_n711), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n799), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G137), .ZN(G39));
  AND3_X1   g624(.A1(new_n806), .A2(KEYINPUT47), .A3(new_n358), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT47), .B1(new_n806), .B2(new_n358), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n768), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n815), .A2(new_n351), .A3(new_n773), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n814), .A2(new_n304), .A3(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G140), .ZN(G42));
  INV_X1    g632(.A(new_n790), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n819), .A2(new_n351), .A3(new_n358), .A4(new_n499), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n745), .A2(new_n445), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n820), .B1(KEYINPUT49), .B2(new_n821), .ZN(new_n822));
  XOR2_X1   g636(.A(new_n822), .B(KEYINPUT110), .Z(new_n823));
  OR2_X1    g637(.A1(new_n821), .A2(KEYINPUT49), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n823), .A2(new_n724), .A3(new_n727), .A4(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n570), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n760), .A2(new_n298), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n792), .A2(new_n351), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n815), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n821), .A2(KEYINPUT114), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n358), .B1(new_n821), .B2(KEYINPUT114), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n829), .B1(new_n814), .B2(new_n833), .ZN(new_n834));
  NOR4_X1   g648(.A1(new_n746), .A2(new_n815), .A3(new_n348), .A4(new_n570), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n724), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT117), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n724), .A2(new_n838), .A3(new_n835), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n564), .A2(new_n655), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n837), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n819), .A2(new_n791), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n790), .A2(KEYINPUT43), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n842), .A2(new_n826), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n760), .A2(new_n298), .A3(new_n684), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n746), .A2(new_n815), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n845), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT116), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT116), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n845), .A2(new_n851), .A3(new_n848), .A4(new_n847), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT50), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n499), .B1(new_n725), .B2(new_n726), .ZN(new_n854));
  INV_X1    g668(.A(new_n746), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n853), .B1(new_n856), .B2(new_n828), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n827), .A2(new_n351), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n844), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(KEYINPUT50), .A3(new_n855), .A4(new_n854), .ZN(new_n860));
  AOI22_X1  g674(.A1(new_n850), .A2(new_n852), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n834), .A2(KEYINPUT51), .A3(new_n841), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n841), .A2(new_n861), .ZN(new_n863));
  INV_X1    g677(.A(new_n829), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT115), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n832), .B(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n864), .B1(new_n866), .B2(new_n813), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n862), .B1(new_n868), .B2(KEYINPUT51), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n845), .A2(new_n772), .A3(new_n848), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT48), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n837), .A2(new_n564), .A3(new_n655), .A4(new_n839), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n873));
  INV_X1    g687(.A(new_n568), .ZN(new_n874));
  INV_X1    g688(.A(new_n755), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n874), .B1(new_n859), .B2(new_n875), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n872), .A2(new_n873), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n873), .B1(new_n872), .B2(new_n876), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n871), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n869), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n846), .A2(new_n773), .ZN(new_n882));
  AOI22_X1  g696(.A1(new_n701), .A2(new_n708), .B1(new_n875), .B2(new_n882), .ZN(new_n883));
  NOR4_X1   g697(.A1(new_n728), .A2(new_n500), .A3(new_n702), .A4(new_n703), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n684), .A2(new_n698), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n884), .A2(new_n450), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n886), .B1(new_n722), .B2(new_n723), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n735), .A2(new_n733), .A3(new_n737), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT105), .B1(new_n708), .B2(new_n739), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n883), .B(new_n887), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT52), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n741), .A2(KEYINPUT52), .A3(new_n883), .A4(new_n887), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n706), .A2(new_n707), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n875), .A2(new_n895), .A3(new_n621), .A4(new_n684), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n750), .A2(new_n753), .A3(new_n896), .A4(new_n763), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT111), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n898), .B1(new_n780), .B2(new_n765), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n882), .A2(KEYINPUT111), .A3(new_n450), .A4(new_n768), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n644), .B1(new_n667), .B2(new_n668), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n684), .A2(new_n685), .A3(new_n699), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n769), .A2(new_n895), .A3(new_n902), .A4(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n901), .A2(new_n904), .A3(new_n788), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n897), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n564), .A2(new_n620), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n564), .B2(new_n656), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n499), .B(new_n635), .C1(new_n496), .C2(new_n497), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n688), .B1(new_n631), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n912), .B1(new_n356), .B2(new_n622), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n906), .A2(new_n785), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n881), .B1(new_n894), .B2(new_n914), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n901), .A2(new_n788), .A3(new_n904), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n748), .A2(new_n749), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n895), .A2(new_n351), .A3(new_n657), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n756), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NOR4_X1   g733(.A1(new_n304), .A2(new_n670), .A3(new_n348), .A4(new_n638), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n917), .B1(new_n920), .B2(new_n762), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n916), .A2(new_n913), .A3(new_n919), .A4(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n776), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n783), .A2(new_n774), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT108), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n743), .A2(new_n769), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n925), .B1(new_n926), .B2(new_n773), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n923), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n922), .A2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT113), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n892), .A2(new_n930), .A3(new_n893), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n741), .A2(new_n883), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n932), .A2(KEYINPUT113), .A3(KEYINPUT52), .A4(new_n887), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n929), .A2(new_n931), .A3(KEYINPUT53), .A4(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT54), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n915), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n894), .A2(new_n914), .A3(new_n881), .ZN(new_n937));
  OAI21_X1  g751(.A(KEYINPUT112), .B1(new_n922), .B2(new_n928), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT112), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n906), .A2(new_n785), .A3(new_n939), .A4(new_n913), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n938), .A2(new_n940), .A3(new_n933), .A4(new_n931), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n937), .B1(new_n881), .B2(new_n941), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n880), .B(new_n936), .C1(new_n942), .C2(new_n935), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT119), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OR2_X1    g759(.A1(G952), .A2(G953), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n946), .B1(new_n943), .B2(new_n944), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n825), .B1(new_n945), .B2(new_n947), .ZN(G75));
  NOR2_X1   g762(.A1(new_n189), .A2(G952), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n187), .B1(new_n915), .B2(new_n934), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT56), .B1(new_n951), .B2(G210), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n472), .A2(new_n474), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(new_n480), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT55), .Z(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n950), .B1(new_n952), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n952), .B2(new_n956), .ZN(G51));
  XNOR2_X1  g772(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(new_n446), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n915), .A2(new_n934), .A3(new_n935), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n935), .B1(new_n915), .B2(new_n934), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT121), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g779(.A(KEYINPUT121), .B(new_n960), .C1(new_n961), .C2(new_n962), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n965), .A2(new_n443), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n951), .A2(new_n803), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n949), .B1(new_n967), .B2(new_n968), .ZN(G54));
  NAND2_X1  g783(.A1(KEYINPUT58), .A2(G475), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT122), .Z(new_n971));
  NAND2_X1  g785(.A1(new_n951), .A2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n562), .ZN(new_n973));
  OR3_X1    g787(.A1(new_n972), .A2(KEYINPUT123), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(KEYINPUT123), .B1(new_n972), .B2(new_n973), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n949), .B1(new_n972), .B2(new_n973), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(G60));
  AND2_X1   g791(.A1(new_n649), .A2(new_n650), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n936), .B1(new_n942), .B2(new_n935), .ZN(new_n979));
  XOR2_X1   g793(.A(KEYINPUT124), .B(KEYINPUT59), .Z(new_n980));
  NOR2_X1   g794(.A1(new_n618), .A2(new_n187), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n978), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n978), .B(new_n982), .C1(new_n961), .C2(new_n962), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n950), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n983), .A2(new_n985), .ZN(G63));
  XNOR2_X1  g800(.A(new_n338), .B(KEYINPUT60), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n987), .B1(new_n915), .B2(new_n934), .ZN(new_n988));
  OR2_X1    g802(.A1(new_n988), .A2(new_n345), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n681), .A2(new_n682), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT125), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n989), .A2(new_n950), .A3(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT61), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n989), .A2(KEYINPUT61), .A3(new_n950), .A4(new_n992), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(G66));
  INV_X1    g811(.A(G224), .ZN(new_n998));
  OAI21_X1  g812(.A(G953), .B1(new_n572), .B2(new_n998), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT126), .Z(new_n1000));
  AND3_X1   g814(.A1(new_n913), .A2(new_n919), .A3(new_n921), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n1000), .B1(new_n1001), .B2(G953), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n953), .B1(G898), .B2(new_n189), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1002), .B(new_n1003), .ZN(G69));
  NAND3_X1  g818(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n284), .A2(new_n285), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n550), .A2(new_n551), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1006), .B(new_n1007), .Z(new_n1008));
  NAND2_X1  g822(.A1(new_n731), .A2(new_n932), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(KEYINPUT62), .ZN(new_n1010));
  INV_X1    g824(.A(new_n713), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n1011), .A2(new_n356), .A3(new_n768), .A4(new_n908), .ZN(new_n1012));
  AND3_X1   g826(.A1(new_n809), .A2(new_n817), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT62), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n731), .A2(new_n1014), .A3(new_n932), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1010), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n1005), .B(new_n1008), .C1(new_n1016), .C2(G953), .ZN(new_n1017));
  AND3_X1   g831(.A1(new_n817), .A2(new_n788), .A3(new_n932), .ZN(new_n1018));
  AND2_X1   g832(.A1(new_n772), .A2(new_n884), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n808), .B1(new_n799), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1018), .A2(new_n785), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1021), .A2(KEYINPUT127), .ZN(new_n1022));
  INV_X1    g836(.A(KEYINPUT127), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n1018), .A2(new_n1023), .A3(new_n785), .A4(new_n1020), .ZN(new_n1024));
  AOI21_X1  g838(.A(G953), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  AND3_X1   g839(.A1(new_n412), .A2(G900), .A3(G953), .ZN(new_n1026));
  OR2_X1    g840(.A1(new_n1008), .A2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1017), .B1(new_n1025), .B2(new_n1027), .ZN(G72));
  NAND4_X1  g842(.A1(new_n1010), .A2(new_n1013), .A3(new_n1001), .A4(new_n1015), .ZN(new_n1029));
  NAND2_X1  g843(.A1(G472), .A2(G902), .ZN(new_n1030));
  XOR2_X1   g844(.A(new_n1030), .B(KEYINPUT63), .Z(new_n1031));
  AND2_X1   g845(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n277), .B1(new_n256), .B2(new_n261), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n950), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n282), .A2(new_n286), .A3(new_n193), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n1022), .A2(new_n1001), .A3(new_n1024), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1035), .B1(new_n1036), .B2(new_n1031), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n287), .A2(new_n262), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1038), .A2(new_n1031), .ZN(new_n1039));
  NOR2_X1   g853(.A1(new_n942), .A2(new_n1039), .ZN(new_n1040));
  NOR3_X1   g854(.A1(new_n1034), .A2(new_n1037), .A3(new_n1040), .ZN(G57));
endmodule


