//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 0 0 1 1 1 1 1 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n626, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  NAND3_X1  g035(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g037(.A(KEYINPUT3), .B1(KEYINPUT66), .B2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(G137), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G101), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n469), .A2(new_n471), .A3(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n467), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n466), .A2(new_n474), .ZN(G160));
  OAI21_X1  g050(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(G112), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(new_n470), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(new_n461), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT67), .Z(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(new_n467), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n478), .B1(new_n483), .B2(G124), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n482), .A2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND4_X1  g063(.A1(new_n469), .A2(new_n471), .A3(G138), .A4(new_n467), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(G126), .A2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(KEYINPUT4), .A2(G138), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n481), .A2(new_n494), .ZN(new_n495));
  OR2_X1    g070(.A1(new_n467), .A2(G114), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n491), .A2(new_n495), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(KEYINPUT68), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT68), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT6), .A3(G651), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n502), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G50), .ZN(new_n509));
  XNOR2_X1  g084(.A(new_n509), .B(KEYINPUT69), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(new_n502), .ZN(new_n512));
  NAND3_X1  g087(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n505), .A2(new_n507), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(new_n514), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n515), .A2(new_n504), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n510), .A2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  XNOR2_X1  g096(.A(KEYINPUT73), .B(KEYINPUT7), .ZN(new_n522));
  AND3_X1   g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n522), .B(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n505), .A2(new_n507), .B1(new_n512), .B2(new_n513), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G89), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n514), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n527), .B1(new_n514), .B2(new_n528), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n524), .B(new_n526), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G51), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n516), .A2(G543), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT72), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT72), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n508), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n532), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n531), .A2(new_n537), .ZN(G168));
  NAND2_X1  g113(.A1(new_n534), .A2(new_n536), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G52), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(new_n504), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  OAI211_X1 g118(.A(new_n540), .B(new_n542), .C1(new_n543), .C2(new_n517), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  NAND2_X1  g120(.A1(new_n539), .A2(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(new_n514), .ZN(new_n548));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n550), .A2(G651), .B1(G81), .B2(new_n525), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  INV_X1    g133(.A(KEYINPUT77), .ZN(new_n559));
  INV_X1    g134(.A(G53), .ZN(new_n560));
  AOI211_X1 g135(.A(new_n560), .B(new_n502), .C1(new_n505), .C2(new_n507), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT74), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n561), .A2(KEYINPUT75), .A3(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n516), .A2(G53), .A3(G543), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n563), .B1(new_n566), .B2(new_n562), .ZN(new_n567));
  AND3_X1   g142(.A1(new_n508), .A2(KEYINPUT75), .A3(G53), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n565), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n570), .B1(new_n512), .B2(new_n513), .ZN(new_n571));
  AND2_X1   g146(.A1(G78), .A2(G543), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g148(.A(KEYINPUT76), .B1(new_n525), .B2(G91), .ZN(new_n574));
  AND4_X1   g149(.A1(KEYINPUT76), .A2(new_n516), .A3(new_n514), .A4(G91), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n559), .B1(new_n569), .B2(new_n576), .ZN(new_n577));
  AND4_X1   g152(.A1(KEYINPUT75), .A2(new_n508), .A3(G53), .A4(new_n564), .ZN(new_n578));
  OAI21_X1  g153(.A(KEYINPUT9), .B1(new_n561), .B2(KEYINPUT74), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n561), .A2(KEYINPUT75), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT76), .ZN(new_n582));
  INV_X1    g157(.A(G91), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n517), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n525), .A2(KEYINPUT76), .A3(G91), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n571), .A2(new_n572), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n584), .A2(new_n585), .B1(new_n586), .B2(G651), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n581), .A2(KEYINPUT77), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n577), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G299));
  INV_X1    g165(.A(G168), .ZN(G286));
  NAND2_X1  g166(.A1(new_n508), .A2(G49), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n593));
  INV_X1    g168(.A(G87), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n592), .B(new_n593), .C1(new_n594), .C2(new_n517), .ZN(G288));
  NAND2_X1  g170(.A1(new_n508), .A2(G48), .ZN(new_n596));
  INV_X1    g171(.A(G86), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n517), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(G73), .A2(G543), .ZN(new_n599));
  XOR2_X1   g174(.A(new_n599), .B(KEYINPUT78), .Z(new_n600));
  NAND2_X1  g175(.A1(new_n514), .A2(G61), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n504), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G305));
  AOI22_X1  g179(.A1(new_n539), .A2(G47), .B1(G85), .B2(new_n525), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT79), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n607), .A2(new_n504), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n606), .A2(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n525), .A2(G92), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n539), .A2(G54), .ZN(new_n614));
  NAND2_X1  g189(.A1(G79), .A2(G543), .ZN(new_n615));
  XNOR2_X1  g190(.A(KEYINPUT80), .B(G66), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n548), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G651), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n613), .A2(new_n614), .A3(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n610), .B1(new_n620), .B2(G868), .ZN(G284));
  OAI21_X1  g196(.A(new_n610), .B1(new_n620), .B2(G868), .ZN(G321));
  NAND2_X1  g197(.A1(G286), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(new_n589), .B2(G868), .ZN(G297));
  OAI21_X1  g199(.A(new_n623), .B1(new_n589), .B2(G868), .ZN(G280));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n620), .B1(new_n626), .B2(G860), .ZN(G148));
  NAND2_X1  g202(.A1(new_n620), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n485), .A2(G135), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n483), .A2(G123), .ZN(new_n633));
  OR2_X1    g208(.A1(G99), .A2(G2105), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n634), .B(G2104), .C1(G111), .C2(new_n467), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n632), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n636), .A2(G2096), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(G2096), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT12), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT13), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(G2100), .Z(new_n642));
  NAND3_X1  g217(.A1(new_n637), .A2(new_n638), .A3(new_n642), .ZN(G156));
  INV_X1    g218(.A(KEYINPUT14), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n644), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n647), .B2(new_n646), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n649), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(G14), .A3(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G401));
  XNOR2_X1  g234(.A(G2072), .B(G2078), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT17), .Z(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n666), .B1(new_n662), .B2(new_n660), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT81), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n665), .A2(new_n662), .A3(new_n660), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT18), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n666), .A2(new_n662), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n671), .B1(new_n661), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT82), .ZN(new_n675));
  XOR2_X1   g250(.A(G2096), .B(G2100), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G227));
  XOR2_X1   g252(.A(KEYINPUT83), .B(KEYINPUT19), .Z(new_n678));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1956), .B(G2474), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1961), .B(G1966), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT20), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n681), .A2(new_n682), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n686), .A2(new_n683), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n685), .B(new_n687), .C1(new_n680), .C2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT84), .ZN(new_n690));
  XOR2_X1   g265(.A(G1981), .B(G1986), .Z(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n690), .B(new_n695), .ZN(G229));
  INV_X1    g271(.A(G29), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G32), .ZN(new_n698));
  NAND3_X1  g273(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT92), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT26), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  AND3_X1   g277(.A1(new_n467), .A2(G105), .A3(G2104), .ZN(new_n703));
  AOI211_X1 g278(.A(new_n702), .B(new_n703), .C1(new_n483), .C2(G129), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n485), .A2(G141), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n698), .B1(new_n707), .B2(new_n697), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT27), .B(G1996), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G4), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(new_n620), .B2(new_n712), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(G1348), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n708), .A2(new_n710), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(G1348), .ZN(new_n717));
  NAND4_X1  g292(.A1(new_n711), .A2(new_n715), .A3(new_n716), .A4(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G2090), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n697), .A2(G35), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G162), .B2(new_n697), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT29), .Z(new_n722));
  AOI21_X1  g297(.A(new_n718), .B1(new_n719), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n697), .A2(G33), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT25), .Z(new_n726));
  AND2_X1   g301(.A1(new_n469), .A2(new_n471), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n727), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n726), .B1(new_n728), .B2(new_n467), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n485), .B2(G139), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n724), .B1(new_n730), .B2(new_n697), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G2072), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT24), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n697), .B1(new_n733), .B2(G34), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n733), .B2(G34), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G160), .B2(G29), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n736), .A2(G2084), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n732), .B1(KEYINPUT95), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(G168), .A2(new_n712), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n712), .B2(G21), .ZN(new_n740));
  INV_X1    g315(.A(G1966), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT93), .ZN(new_n743));
  AOI211_X1 g318(.A(new_n738), .B(new_n743), .C1(KEYINPUT95), .C2(new_n737), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n697), .A2(G26), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT28), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n485), .A2(G140), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n483), .A2(G128), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n467), .A2(G116), .ZN(new_n749));
  OAI21_X1  g324(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n747), .B(new_n748), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G29), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n752), .A2(KEYINPUT91), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n752), .A2(KEYINPUT91), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n746), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G2067), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n636), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n758), .A2(G29), .B1(G2084), .B2(new_n736), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n740), .A2(new_n741), .ZN(new_n760));
  INV_X1    g335(.A(G28), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n761), .A2(KEYINPUT30), .ZN(new_n762));
  AOI21_X1  g337(.A(G29), .B1(new_n761), .B2(KEYINPUT30), .ZN(new_n763));
  OR2_X1    g338(.A1(KEYINPUT31), .A2(G11), .ZN(new_n764));
  NAND2_X1  g339(.A1(KEYINPUT31), .A2(G11), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n762), .A2(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(G164), .A2(G29), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G27), .B2(G29), .ZN(new_n768));
  INV_X1    g343(.A(G2078), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n766), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n769), .B2(new_n768), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n712), .A2(G19), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n553), .B2(new_n712), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G1341), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n759), .A2(new_n760), .A3(new_n771), .A4(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G5), .A2(G16), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT94), .Z(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G301), .B2(new_n712), .ZN(new_n778));
  INV_X1    g353(.A(G1961), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G1341), .B2(new_n773), .ZN(new_n781));
  OAI22_X1  g356(.A1(new_n731), .A2(G2072), .B1(new_n778), .B2(new_n779), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n775), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n723), .A2(new_n744), .A3(new_n757), .A4(new_n783), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n722), .A2(new_n719), .ZN(new_n785));
  NAND2_X1  g360(.A1(G299), .A2(G16), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT96), .B(KEYINPUT23), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n712), .A2(G20), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G1956), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n785), .A2(KEYINPUT97), .A3(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(KEYINPUT97), .B1(new_n785), .B2(new_n792), .ZN(new_n795));
  NOR3_X1   g370(.A1(new_n784), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  MUX2_X1   g371(.A(G23), .B(G288), .S(G16), .Z(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT88), .Z(new_n798));
  XOR2_X1   g373(.A(KEYINPUT33), .B(G1976), .Z(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n798), .A2(new_n800), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n712), .A2(G22), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G166), .B2(new_n712), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n804), .A2(G1971), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(G1971), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n801), .A2(new_n802), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n712), .A2(G6), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n603), .B2(new_n712), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT87), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT32), .B(G1981), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT86), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n810), .B(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT89), .ZN(new_n814));
  OR3_X1    g389(.A1(new_n807), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n807), .B2(new_n813), .ZN(new_n816));
  AOI21_X1  g391(.A(KEYINPUT34), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n697), .A2(G25), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n467), .A2(G107), .ZN(new_n819));
  OAI21_X1  g394(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n483), .A2(G119), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n485), .A2(G131), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n818), .B1(new_n824), .B2(new_n697), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT35), .B(G1991), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT85), .Z(new_n827));
  INV_X1    g402(.A(KEYINPUT90), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT36), .ZN(new_n829));
  OAI22_X1  g404(.A1(new_n825), .A2(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(new_n827), .B2(new_n825), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n712), .A2(G24), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n606), .A2(new_n608), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(new_n712), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n834), .A2(G1986), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(G1986), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n831), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n817), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n828), .A2(new_n829), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n815), .A2(KEYINPUT34), .A3(new_n816), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n796), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n839), .B1(new_n838), .B2(new_n840), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n842), .A2(new_n843), .ZN(G311));
  INV_X1    g419(.A(new_n843), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n845), .A2(new_n841), .A3(new_n796), .ZN(G150));
  NAND2_X1  g421(.A1(new_n620), .A2(G559), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT38), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n539), .A2(G55), .ZN(new_n849));
  NAND2_X1  g424(.A1(G80), .A2(G543), .ZN(new_n850));
  INV_X1    g425(.A(G67), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n850), .B1(new_n548), .B2(new_n851), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n852), .A2(G651), .B1(G93), .B2(new_n525), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n552), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n546), .A2(new_n849), .A3(new_n551), .A4(new_n853), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n848), .B(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n859));
  AOI21_X1  g434(.A(G860), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(new_n859), .B2(new_n858), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n854), .A2(G860), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT98), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT37), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(KEYINPUT99), .Z(G145));
  XNOR2_X1  g441(.A(KEYINPUT102), .B(G37), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n487), .B(new_n636), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT100), .ZN(new_n869));
  INV_X1    g444(.A(G160), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n751), .B(new_n500), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n485), .A2(G142), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n483), .A2(G130), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n467), .A2(G118), .ZN(new_n875));
  OAI21_X1  g450(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n873), .B(new_n874), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n872), .B(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n706), .B(new_n730), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n824), .A2(KEYINPUT101), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n822), .A2(new_n823), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n640), .ZN(new_n887));
  INV_X1    g462(.A(new_n640), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n882), .A2(new_n888), .A3(new_n885), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n881), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(new_n889), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n891), .A2(new_n880), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n879), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n869), .A2(new_n870), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n891), .A2(new_n880), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n881), .A2(new_n887), .A3(new_n889), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n895), .A2(new_n896), .A3(new_n878), .ZN(new_n897));
  AND4_X1   g472(.A1(new_n871), .A2(new_n893), .A3(new_n894), .A4(new_n897), .ZN(new_n898));
  AOI22_X1  g473(.A1(new_n893), .A2(new_n897), .B1(new_n871), .B2(new_n894), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n867), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n900), .B(new_n901), .ZN(G395));
  XOR2_X1   g477(.A(new_n603), .B(G288), .Z(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(G290), .A2(G166), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(G290), .A2(G166), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n907), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n909), .A2(new_n903), .A3(new_n905), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT42), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n589), .A2(new_n619), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n620), .A2(new_n577), .A3(new_n588), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n913), .A2(new_n914), .A3(KEYINPUT41), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n628), .B(new_n857), .ZN(new_n920));
  MUX2_X1   g495(.A(new_n919), .B(new_n915), .S(new_n920), .Z(new_n921));
  XNOR2_X1  g496(.A(new_n912), .B(new_n921), .ZN(new_n922));
  MUX2_X1   g497(.A(new_n854), .B(new_n922), .S(G868), .Z(G295));
  MUX2_X1   g498(.A(new_n854), .B(new_n922), .S(G868), .Z(G331));
  AND3_X1   g499(.A1(new_n855), .A2(G301), .A3(new_n856), .ZN(new_n925));
  AOI21_X1  g500(.A(G301), .B1(new_n855), .B2(new_n856), .ZN(new_n926));
  OAI21_X1  g501(.A(G286), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n857), .A2(G171), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n855), .A2(G301), .A3(new_n856), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(G168), .A3(new_n929), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n919), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT104), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n908), .A2(new_n910), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n927), .A2(new_n930), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n915), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n931), .A2(new_n919), .A3(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n933), .A2(new_n934), .A3(new_n936), .A4(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(G37), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n938), .A2(new_n936), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n934), .B1(new_n942), .B2(new_n933), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT43), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n931), .B1(new_n946), .B2(new_n918), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n919), .A2(KEYINPUT105), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n936), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n911), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n950), .A2(new_n951), .A3(new_n939), .A4(new_n867), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n944), .A2(new_n945), .A3(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n941), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n938), .A2(new_n936), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n937), .B1(new_n931), .B2(new_n919), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n911), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n954), .A2(new_n955), .A3(new_n951), .A4(new_n958), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n958), .A2(new_n951), .A3(new_n939), .A4(new_n940), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(KEYINPUT106), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n950), .A2(new_n867), .A3(new_n939), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n959), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n953), .B1(KEYINPUT44), .B2(new_n964), .ZN(G397));
  INV_X1    g540(.A(KEYINPUT112), .ZN(new_n966));
  INV_X1    g541(.A(G1971), .ZN(new_n967));
  INV_X1    g542(.A(new_n474), .ZN(new_n968));
  INV_X1    g543(.A(G137), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n969), .B1(new_n480), .B2(new_n461), .ZN(new_n970));
  INV_X1    g545(.A(new_n465), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n467), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n968), .A2(new_n972), .A3(G40), .ZN(new_n973));
  INV_X1    g548(.A(G1384), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT45), .B1(new_n500), .B2(new_n974), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n973), .B(new_n975), .C1(new_n976), .C2(new_n977), .ZN(new_n978));
  AOI22_X1  g553(.A1(new_n481), .A2(new_n494), .B1(new_n496), .B2(new_n498), .ZN(new_n979));
  AOI21_X1  g554(.A(G1384), .B1(new_n979), .B2(new_n491), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n980), .A2(KEYINPUT110), .A3(KEYINPUT45), .ZN(new_n981));
  OAI211_X1 g556(.A(KEYINPUT111), .B(new_n967), .C1(new_n978), .C2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n983));
  OAI211_X1 g558(.A(G160), .B(G40), .C1(new_n980), .C2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n980), .A2(new_n983), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n719), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n982), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n500), .A2(new_n974), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n990), .A2(new_n977), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT110), .B1(new_n980), .B2(KEYINPUT45), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n992), .A2(new_n993), .A3(new_n973), .A4(new_n975), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT111), .B1(new_n994), .B2(new_n967), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n966), .B1(new_n989), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n967), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n999), .A2(KEYINPUT112), .A3(new_n988), .A4(new_n982), .ZN(new_n1000));
  NAND2_X1  g575(.A1(G303), .A2(G8), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n996), .A2(new_n1000), .A3(G8), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n973), .A2(new_n980), .ZN(new_n1005));
  INV_X1    g580(.A(G1976), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1005), .B(G8), .C1(new_n1006), .C2(G288), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n1007), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT113), .B1(new_n1007), .B2(KEYINPUT52), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G1981), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n603), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n598), .A2(new_n602), .A3(G1981), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1013), .A2(KEYINPUT49), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT49), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1017), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n968), .A2(new_n972), .A3(G40), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n990), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G8), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1016), .A2(new_n1018), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT52), .B1(G288), .B2(new_n1006), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n1024), .B(KEYINPUT114), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1023), .B1(new_n1007), .B2(new_n1025), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n1004), .A2(new_n1010), .A3(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(G288), .A2(G1976), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1014), .B1(new_n1023), .B2(new_n1028), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1029), .A2(KEYINPUT115), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1022), .B1(new_n1029), .B2(KEYINPUT115), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1027), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1001), .B(KEYINPUT55), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n997), .A2(new_n988), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1034), .B1(new_n1021), .B2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1026), .A2(new_n1010), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1004), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n1039));
  AOI211_X1 g614(.A(new_n991), .B(G1384), .C1(new_n979), .C2(new_n491), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n976), .A2(new_n1040), .A3(new_n1019), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(G2078), .ZN(new_n1043));
  MUX2_X1   g618(.A(G2078), .B(new_n1043), .S(KEYINPUT121), .Z(new_n1044));
  NAND2_X1  g619(.A1(new_n990), .A2(KEYINPUT50), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1045), .A2(new_n973), .A3(new_n985), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1041), .A2(new_n1044), .B1(new_n1046), .B2(new_n779), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1040), .A2(new_n1019), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1048), .A2(new_n769), .A3(new_n992), .A4(new_n993), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n1042), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1047), .A2(new_n1050), .A3(G301), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1041), .A2(new_n1043), .B1(new_n1046), .B2(new_n779), .ZN(new_n1052));
  AOI21_X1  g627(.A(G301), .B1(new_n1052), .B2(new_n1050), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1039), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT122), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT122), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1056), .B(new_n1039), .C1(new_n1051), .C2(new_n1053), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT120), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1059), .B1(G168), .B2(new_n1021), .ZN(new_n1060));
  OAI211_X1 g635(.A(KEYINPUT120), .B(G8), .C1(new_n531), .C2(new_n537), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT51), .ZN(new_n1063));
  XOR2_X1   g638(.A(KEYINPUT116), .B(G2084), .Z(new_n1064));
  INV_X1    g639(.A(new_n976), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1065), .A2(new_n973), .A3(new_n975), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n987), .A2(new_n1064), .B1(new_n1066), .B2(new_n741), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1062), .B(new_n1063), .C1(new_n1067), .C2(new_n1021), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT51), .B1(new_n1062), .B2(new_n1067), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1019), .B1(new_n990), .B2(KEYINPUT50), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1071), .A2(new_n985), .A3(new_n1064), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(G1966), .B2(new_n1041), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1070), .B1(new_n1073), .B2(G8), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1068), .B1(new_n1069), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1052), .A2(new_n1050), .A3(G301), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT54), .ZN(new_n1077));
  AOI21_X1  g652(.A(G301), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT123), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1047), .A2(new_n1050), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(G171), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT123), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1081), .A2(new_n1082), .A3(KEYINPUT54), .A4(new_n1076), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1075), .B1(new_n1079), .B2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1038), .A2(new_n1058), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G1348), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1046), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1020), .A2(new_n756), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n619), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1090), .B(new_n565), .C1(new_n567), .C2(new_n568), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1091), .B(new_n1092), .C1(new_n569), .C2(new_n576), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n581), .B(new_n587), .C1(new_n1090), .C2(KEYINPUT57), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  XNOR2_X1  g670(.A(KEYINPUT56), .B(G2072), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1048), .A2(new_n992), .A3(new_n993), .A4(new_n1096), .ZN(new_n1097));
  XOR2_X1   g672(.A(KEYINPUT117), .B(G1956), .Z(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(new_n984), .B2(new_n986), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1089), .B1(new_n1095), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT60), .ZN(new_n1102));
  AOI21_X1  g677(.A(G1348), .B1(new_n1071), .B2(new_n985), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1005), .A2(G2067), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1102), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1087), .A2(KEYINPUT60), .A3(new_n1088), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(new_n1106), .A3(new_n620), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT119), .B(KEYINPUT61), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(new_n1095), .B2(new_n1100), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1087), .A2(KEYINPUT60), .A3(new_n619), .A4(new_n1088), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1107), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n1112));
  INV_X1    g687(.A(G1996), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1048), .A2(new_n1113), .A3(new_n992), .A4(new_n993), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT58), .B(G1341), .Z(new_n1115));
  NAND2_X1  g690(.A1(new_n1005), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1112), .B1(new_n1117), .B2(new_n553), .ZN(new_n1118));
  AOI211_X1 g693(.A(KEYINPUT59), .B(new_n552), .C1(new_n1114), .C2(new_n1116), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1101), .B1(new_n1111), .B2(new_n1120), .ZN(new_n1121));
  OR2_X1    g696(.A1(new_n1095), .A2(new_n1100), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1111), .A2(new_n1120), .ZN(new_n1123));
  AND2_X1   g698(.A1(KEYINPUT119), .A2(KEYINPUT61), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1121), .A2(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1033), .B1(new_n1085), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n996), .A2(G8), .A3(new_n1000), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n1034), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1067), .A2(new_n1021), .A3(G286), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n1129), .A2(KEYINPUT63), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1004), .A2(new_n1037), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT63), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1004), .A2(new_n1037), .A3(new_n1036), .A4(new_n1129), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1131), .A2(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT124), .B1(new_n1126), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1139), .A2(new_n1038), .A3(new_n1058), .A4(new_n1084), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1132), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1134), .A2(new_n1133), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1140), .A2(new_n1141), .A3(new_n1144), .A4(new_n1033), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1075), .ZN(new_n1146));
  OR2_X1    g721(.A1(new_n1146), .A2(KEYINPUT62), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(KEYINPUT62), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1147), .A2(new_n1038), .A3(new_n1053), .A4(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1136), .A2(new_n1145), .A3(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1065), .A2(new_n1019), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n1113), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n706), .A2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1153), .B(KEYINPUT107), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n707), .A2(new_n1113), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n751), .B(G2067), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1151), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT108), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1154), .A2(new_n1157), .A3(KEYINPUT108), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n883), .A2(new_n827), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n883), .A2(new_n827), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1151), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  AND2_X1   g739(.A1(G290), .A2(G1986), .ZN(new_n1165));
  NOR2_X1   g740(.A1(G290), .A2(G1986), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1151), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1160), .A2(new_n1161), .A3(new_n1164), .A4(new_n1167), .ZN(new_n1168));
  XOR2_X1   g743(.A(new_n1168), .B(KEYINPUT109), .Z(new_n1169));
  NAND2_X1  g744(.A1(new_n1150), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n1171));
  XOR2_X1   g746(.A(new_n1163), .B(KEYINPUT125), .Z(new_n1172));
  NAND3_X1  g747(.A1(new_n1160), .A2(new_n1161), .A3(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n751), .A2(G2067), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1174), .ZN(new_n1175));
  AOI211_X1 g750(.A(new_n1065), .B(new_n1019), .C1(new_n1173), .C2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1166), .A2(new_n1151), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT48), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1160), .A2(new_n1178), .A3(new_n1161), .A4(new_n1164), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1151), .B1(new_n1156), .B2(new_n706), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1152), .B(KEYINPUT46), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1182), .B(KEYINPUT47), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1179), .A2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1171), .B1(new_n1176), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(new_n1151), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1187), .A2(KEYINPUT126), .A3(new_n1183), .A4(new_n1179), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1170), .A2(new_n1189), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g765(.A1(G229), .A2(new_n459), .A3(G401), .ZN(new_n1192));
  INV_X1    g766(.A(KEYINPUT127), .ZN(new_n1193));
  OR3_X1    g767(.A1(new_n1192), .A2(new_n1193), .A3(G227), .ZN(new_n1194));
  OAI21_X1  g768(.A(new_n1193), .B1(new_n1192), .B2(G227), .ZN(new_n1195));
  NAND2_X1  g769(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g770(.A1(new_n944), .A2(new_n952), .ZN(new_n1197));
  NAND3_X1  g771(.A1(new_n1196), .A2(new_n900), .A3(new_n1197), .ZN(G225));
  INV_X1    g772(.A(G225), .ZN(G308));
endmodule


