//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 1 1 1 0 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1334, new_n1335, new_n1336, new_n1337, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1397, new_n1398, new_n1399, new_n1400, new_n1401;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n210), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G68), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  INV_X1    g0024(.A(G87), .ZN(new_n225));
  INV_X1    g0025(.A(G250), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n228));
  INV_X1    g0028(.A(G58), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  INV_X1    g0030(.A(G257), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n228), .B1(new_n229), .B2(new_n230), .C1(new_n205), .C2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n212), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n215), .B(new_n221), .C1(KEYINPUT1), .C2(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n230), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n202), .A2(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n223), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n246), .B(new_n251), .Z(G351));
  NAND2_X1  g0052(.A1(new_n203), .A2(G20), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  OAI21_X1  g0054(.A(KEYINPUT65), .B1(new_n254), .B2(G20), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT65), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(new_n210), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT8), .B(G58), .ZN(new_n259));
  OAI21_X1  g0059(.A(KEYINPUT66), .B1(G20), .B2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NOR3_X1   g0061(.A1(KEYINPUT66), .A2(G20), .A3(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G150), .ZN(new_n264));
  OAI221_X1 g0064(.A(new_n253), .B1(new_n258), .B2(new_n259), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n219), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n209), .A2(G20), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G50), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n270), .B(KEYINPUT67), .ZN(new_n271));
  INV_X1    g0071(.A(G13), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G1), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G20), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n275), .A2(new_n267), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n271), .A2(new_n276), .B1(new_n202), .B2(new_n275), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n268), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G169), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(G1), .A3(G13), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT3), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n254), .ZN(new_n284));
  NAND2_X1  g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G1698), .ZN(new_n287));
  INV_X1    g0087(.A(G223), .ZN(new_n288));
  INV_X1    g0088(.A(G77), .ZN(new_n289));
  OAI22_X1  g0089(.A1(new_n287), .A2(new_n288), .B1(new_n289), .B2(new_n286), .ZN(new_n290));
  INV_X1    g0090(.A(G1698), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n286), .A2(G222), .A3(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n282), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT64), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G41), .A2(G45), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n295), .B1(new_n296), .B2(G1), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n209), .B(KEYINPUT64), .C1(G41), .C2(G45), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G274), .ZN(new_n300));
  AND2_X1   g0100(.A1(G1), .A2(G13), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n300), .B1(new_n301), .B2(new_n280), .ZN(new_n302));
  INV_X1    g0102(.A(G41), .ZN(new_n303));
  INV_X1    g0103(.A(G45), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n209), .A2(new_n305), .B1(new_n301), .B2(new_n280), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n299), .A2(new_n302), .B1(new_n306), .B2(G226), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n294), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n278), .B1(new_n279), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G179), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n294), .A2(new_n310), .A3(new_n307), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT10), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n268), .A2(new_n277), .A3(KEYINPUT9), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n315), .B(KEYINPUT69), .ZN(new_n316));
  INV_X1    g0116(.A(G190), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n308), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G200), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(new_n294), .B2(new_n307), .ZN(new_n320));
  AOI21_X1  g0120(.A(KEYINPUT9), .B1(new_n268), .B2(new_n277), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n318), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n314), .B1(new_n316), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n316), .A2(new_n322), .A3(new_n314), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n313), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n276), .A2(G77), .A3(new_n269), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT15), .B(G87), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n258), .A2(new_n328), .B1(new_n210), .B2(new_n289), .ZN(new_n329));
  INV_X1    g0129(.A(new_n262), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n260), .ZN(new_n331));
  INV_X1    g0131(.A(new_n259), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n329), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n267), .ZN(new_n334));
  OAI221_X1 g0134(.A(new_n327), .B1(G77), .B2(new_n274), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n286), .A2(G232), .A3(new_n291), .ZN(new_n336));
  OAI221_X1 g0136(.A(new_n336), .B1(new_n206), .B2(new_n286), .C1(new_n287), .C2(new_n224), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n282), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT68), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n299), .A2(new_n302), .B1(new_n306), .B2(G244), .ZN(new_n340));
  AND3_X1   g0140(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n339), .B1(new_n338), .B2(new_n340), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n335), .B1(new_n343), .B2(G200), .ZN(new_n344));
  OAI21_X1  g0144(.A(G190), .B1(new_n341), .B2(new_n342), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n343), .A2(new_n279), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n310), .B1(new_n341), .B2(new_n342), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n347), .A2(new_n335), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT70), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n326), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  AND3_X1   g0153(.A1(new_n316), .A2(new_n322), .A3(new_n314), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n312), .B1(new_n354), .B2(new_n323), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT70), .B1(new_n355), .B2(new_n350), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n259), .B1(new_n209), .B2(G20), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n276), .A2(new_n358), .B1(new_n275), .B2(new_n259), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  AND2_X1   g0160(.A1(KEYINPUT3), .A2(G33), .ZN(new_n361));
  NOR2_X1   g0161(.A1(KEYINPUT3), .A2(G33), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT7), .B1(new_n363), .B2(new_n210), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT7), .ZN(new_n365));
  NOR4_X1   g0165(.A1(new_n361), .A2(new_n362), .A3(new_n365), .A4(G20), .ZN(new_n366));
  OAI21_X1  g0166(.A(G68), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g0167(.A(G58), .B(G68), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n331), .A2(G159), .B1(new_n368), .B2(G20), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT16), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n334), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n367), .A2(KEYINPUT16), .A3(new_n369), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n360), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI211_X1 g0174(.A(G223), .B(new_n291), .C1(new_n361), .C2(new_n362), .ZN(new_n375));
  OAI211_X1 g0175(.A(G226), .B(G1698), .C1(new_n361), .C2(new_n362), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G33), .A2(G87), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n282), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n299), .A2(new_n302), .B1(new_n306), .B2(G232), .ZN(new_n380));
  AOI21_X1  g0180(.A(G169), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n379), .A2(new_n380), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n382), .B1(G179), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT18), .B1(new_n374), .B2(new_n384), .ZN(new_n385));
  AND3_X1   g0185(.A1(new_n379), .A2(new_n380), .A3(G190), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n319), .B1(new_n379), .B2(new_n380), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n284), .A2(new_n210), .A3(new_n285), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n365), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n363), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n223), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n368), .A2(G20), .ZN(new_n393));
  INV_X1    g0193(.A(G159), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n393), .B1(new_n263), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n371), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(new_n373), .A3(new_n267), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n388), .A2(new_n397), .A3(new_n359), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT17), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n374), .A2(KEYINPUT17), .A3(new_n388), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n397), .A2(new_n359), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT18), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n383), .A2(G179), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n404), .A2(new_n381), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n402), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n385), .A2(new_n400), .A3(new_n401), .A4(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  OAI211_X1 g0208(.A(G232), .B(G1698), .C1(new_n361), .C2(new_n362), .ZN(new_n409));
  OAI211_X1 g0209(.A(G226), .B(new_n291), .C1(new_n361), .C2(new_n362), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G97), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n282), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n299), .A2(new_n302), .B1(new_n306), .B2(G238), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT13), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n415), .B1(new_n413), .B2(new_n414), .ZN(new_n417));
  OAI21_X1  g0217(.A(G169), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT14), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT14), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n420), .B(G169), .C1(new_n416), .C2(new_n417), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n413), .A2(new_n414), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT71), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n413), .A2(new_n414), .A3(KEYINPUT71), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(KEYINPUT13), .A3(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n416), .A2(new_n310), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT72), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n427), .A2(new_n428), .A3(KEYINPUT72), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n422), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(KEYINPUT12), .B1(new_n274), .B2(G68), .ZN(new_n433));
  OR3_X1    g0233(.A1(new_n274), .A2(KEYINPUT12), .A3(G68), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n223), .B1(new_n209), .B2(G20), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n433), .A2(new_n434), .B1(new_n276), .B2(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n263), .A2(new_n202), .ZN(new_n437));
  OAI22_X1  g0237(.A1(new_n258), .A2(new_n289), .B1(new_n210), .B2(G68), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n267), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT11), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n436), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n439), .A2(new_n440), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n432), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n416), .A2(new_n317), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n427), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(G200), .B1(new_n416), .B2(new_n417), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n444), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n357), .A2(new_n408), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT85), .ZN(new_n453));
  INV_X1    g0253(.A(G116), .ZN(new_n454));
  AOI221_X4 g0254(.A(KEYINPUT83), .B1(new_n454), .B2(G20), .C1(new_n266), .C2(new_n219), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT83), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(G20), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n456), .B1(new_n267), .B2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G283), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n460), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT84), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n254), .A2(G97), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n464), .A2(KEYINPUT84), .A3(new_n210), .A4(new_n460), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(KEYINPUT20), .B1(new_n459), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n459), .A2(KEYINPUT20), .A3(new_n466), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n209), .A2(G33), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n334), .A2(new_n274), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G116), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n274), .A2(new_n454), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n468), .A2(new_n469), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(G257), .B(new_n291), .C1(new_n361), .C2(new_n362), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT82), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n286), .A2(KEYINPUT82), .A3(G257), .A4(new_n291), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n363), .A2(G303), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n286), .A2(G264), .A3(G1698), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n477), .A2(new_n478), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n282), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n304), .A2(G1), .ZN(new_n483));
  NAND2_X1  g0283(.A1(KEYINPUT5), .A2(G41), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(G270), .A3(new_n281), .ZN(new_n488));
  INV_X1    g0288(.A(new_n486), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n484), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(new_n302), .A3(new_n483), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT81), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n488), .A2(new_n491), .A3(KEYINPUT81), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n482), .B(G179), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n453), .B1(new_n474), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n472), .A2(new_n473), .ZN(new_n496));
  INV_X1    g0296(.A(new_n458), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n267), .A2(new_n456), .A3(new_n457), .ZN(new_n498));
  AND4_X1   g0298(.A1(KEYINPUT20), .A2(new_n466), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n496), .B1(new_n499), .B2(new_n467), .ZN(new_n500));
  INV_X1    g0300(.A(new_n492), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n488), .A2(new_n491), .A3(KEYINPUT81), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n501), .A2(new_n502), .B1(new_n481), .B2(new_n282), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n500), .A2(new_n503), .A3(KEYINPUT85), .A4(G179), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n495), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n482), .B1(new_n492), .B2(new_n493), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n500), .B1(G200), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(new_n317), .B2(new_n506), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n500), .A2(G169), .A3(new_n506), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n509), .A2(KEYINPUT86), .A3(KEYINPUT21), .ZN(new_n510));
  AOI21_X1  g0310(.A(KEYINPUT21), .B1(new_n509), .B2(KEYINPUT86), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n505), .B(new_n508), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(G244), .B(new_n291), .C1(new_n361), .C2(new_n362), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT4), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n460), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI211_X1 g0315(.A(G250), .B(G1698), .C1(new_n361), .C2(new_n362), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT75), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n286), .A2(KEYINPUT75), .A3(G250), .A4(G1698), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n513), .A2(KEYINPUT74), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT74), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n286), .A2(new_n522), .A3(G244), .A4(new_n291), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(new_n523), .A3(new_n514), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n281), .B1(new_n520), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n487), .A2(G257), .A3(new_n281), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n491), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT76), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT76), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n526), .A2(new_n491), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(KEYINPUT77), .B1(new_n525), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n515), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n518), .A2(new_n519), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n524), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n282), .ZN(new_n536));
  INV_X1    g0336(.A(new_n530), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n529), .B1(new_n526), .B2(new_n491), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT77), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n536), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n532), .A2(G190), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n536), .A2(new_n539), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G200), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT6), .ZN(new_n545));
  NOR3_X1   g0345(.A1(new_n545), .A2(new_n205), .A3(G107), .ZN(new_n546));
  XNOR2_X1  g0346(.A(G97), .B(G107), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n546), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  OAI22_X1  g0348(.A1(new_n548), .A2(new_n210), .B1(new_n289), .B2(new_n263), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n206), .B1(new_n390), .B2(new_n391), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n267), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n471), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G97), .ZN(new_n553));
  OR3_X1    g0353(.A1(new_n274), .A2(KEYINPUT73), .A3(G97), .ZN(new_n554));
  OAI21_X1  g0354(.A(KEYINPUT73), .B1(new_n274), .B2(G97), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n551), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n544), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(G169), .B1(new_n532), .B2(new_n541), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n536), .A2(new_n539), .A3(new_n310), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n557), .ZN(new_n562));
  OAI22_X1  g0362(.A1(new_n542), .A2(new_n559), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n275), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT25), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n274), .B2(G107), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n552), .A2(G107), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n210), .A2(G33), .A3(G116), .ZN(new_n569));
  NOR2_X1   g0369(.A1(KEYINPUT88), .A2(KEYINPUT23), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n570), .A2(G20), .A3(new_n206), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT89), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n572), .A2(KEYINPUT24), .B1(KEYINPUT88), .B2(KEYINPUT23), .ZN(new_n573));
  OAI22_X1  g0373(.A1(new_n210), .A2(G107), .B1(KEYINPUT88), .B2(KEYINPUT23), .ZN(new_n574));
  AND4_X1   g0374(.A1(new_n569), .A2(new_n571), .A3(new_n573), .A4(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n210), .A2(KEYINPUT87), .A3(G87), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n363), .A2(KEYINPUT22), .A3(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT22), .ZN(new_n578));
  INV_X1    g0378(.A(new_n576), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n578), .B1(new_n286), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n575), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT24), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(KEYINPUT89), .ZN(new_n583));
  XNOR2_X1  g0383(.A(new_n581), .B(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n568), .B1(new_n584), .B2(new_n267), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n487), .A2(G264), .A3(new_n281), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G33), .A2(G294), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n226), .A2(new_n291), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n231), .A2(G1698), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n588), .B1(new_n591), .B2(new_n286), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n491), .B(new_n586), .C1(new_n592), .C2(new_n281), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n319), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(G190), .B2(new_n593), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n585), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n581), .A2(new_n583), .ZN(new_n597));
  OAI21_X1  g0397(.A(KEYINPUT22), .B1(new_n363), .B2(new_n576), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n286), .A2(new_n579), .A3(new_n578), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n600), .A2(new_n575), .B1(KEYINPUT89), .B2(new_n582), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n267), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n567), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n593), .A2(G169), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n589), .B(new_n590), .C1(new_n361), .C2(new_n362), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n281), .B1(new_n605), .B2(new_n587), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n607), .A2(G179), .A3(new_n491), .A4(new_n586), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT90), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n604), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n604), .A2(new_n608), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT90), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n603), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n328), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n614), .A2(new_n274), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n471), .A2(new_n225), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT19), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n258), .B2(new_n205), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n286), .A2(KEYINPUT80), .A3(new_n210), .A4(G68), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n210), .B1(new_n411), .B2(new_n617), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(G87), .B2(new_n207), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT80), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n210), .A2(G68), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n622), .B1(new_n363), .B2(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n618), .A2(new_n619), .A3(new_n621), .A4(new_n624), .ZN(new_n625));
  AOI211_X1 g0425(.A(new_n615), .B(new_n616), .C1(new_n625), .C2(new_n267), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n226), .B1(new_n209), .B2(G45), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT78), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n627), .A2(new_n281), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n281), .A2(G274), .A3(new_n483), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n628), .B1(new_n627), .B2(new_n281), .ZN(new_n632));
  OAI21_X1  g0432(.A(KEYINPUT79), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n627), .A2(new_n281), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT78), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT79), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n635), .A2(new_n636), .A3(new_n630), .A4(new_n629), .ZN(new_n637));
  INV_X1    g0437(.A(G244), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(G1698), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(G238), .B2(G1698), .ZN(new_n640));
  OAI22_X1  g0440(.A1(new_n640), .A2(new_n363), .B1(new_n254), .B2(new_n454), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n282), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n633), .A2(new_n637), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(G200), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n633), .A2(G190), .A3(new_n637), .A4(new_n642), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n626), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n615), .B1(new_n625), .B2(new_n267), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n647), .B1(new_n471), .B2(new_n328), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n643), .A2(new_n279), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n633), .A2(new_n310), .A3(new_n637), .A4(new_n642), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n596), .A2(new_n613), .A3(new_n646), .A4(new_n651), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n512), .A2(new_n563), .A3(new_n652), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n452), .A2(new_n653), .ZN(G372));
  AND2_X1   g0454(.A1(new_n400), .A2(new_n401), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n349), .A2(new_n449), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n655), .B1(new_n444), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT94), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n402), .A2(new_n403), .A3(new_n405), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n403), .B1(new_n402), .B2(new_n405), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n385), .A2(KEYINPUT94), .A3(new_n406), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n657), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n354), .A2(new_n323), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n313), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT91), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n254), .A2(new_n454), .ZN(new_n668));
  NOR2_X1   g0468(.A1(G238), .A2(G1698), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n669), .B1(new_n638), .B2(G1698), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n668), .B1(new_n670), .B2(new_n286), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n667), .B1(new_n671), .B2(new_n281), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n641), .A2(KEYINPUT91), .A3(new_n282), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n633), .A2(new_n672), .A3(new_n637), .A4(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n279), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n675), .A2(KEYINPUT92), .A3(new_n650), .ZN(new_n676));
  AOI21_X1  g0476(.A(KEYINPUT92), .B1(new_n675), .B2(new_n650), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n648), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n626), .A2(new_n645), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n674), .A2(G200), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n678), .A2(new_n596), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(KEYINPUT93), .B1(new_n683), .B2(new_n563), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n675), .A2(new_n650), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT92), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n675), .A2(KEYINPUT92), .A3(new_n650), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n681), .B1(new_n689), .B2(new_n648), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n525), .A2(KEYINPUT77), .A3(new_n531), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n540), .B1(new_n536), .B2(new_n539), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n279), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n562), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n532), .A2(G190), .A3(new_n541), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n557), .B1(new_n543), .B2(G200), .ZN(new_n696));
  AOI22_X1  g0496(.A1(new_n693), .A2(new_n694), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT93), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n690), .A2(new_n697), .A3(new_n698), .A4(new_n596), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n510), .A2(new_n511), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n603), .A2(new_n611), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(new_n505), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n684), .A2(new_n699), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n532), .A2(new_n541), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n562), .B1(new_n704), .B2(new_n279), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n651), .A2(new_n646), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(KEYINPUT26), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT26), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n705), .A2(new_n678), .A3(new_n709), .A4(new_n682), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n708), .A2(new_n678), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n703), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n666), .B1(new_n451), .B2(new_n713), .ZN(G369));
  NAND2_X1  g0514(.A1(new_n596), .A2(new_n613), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n273), .A2(new_n210), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n716), .A2(KEYINPUT27), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(KEYINPUT27), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(G213), .A3(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(G343), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n585), .A2(new_n722), .ZN(new_n723));
  OAI22_X1  g0523(.A1(new_n715), .A2(new_n723), .B1(new_n613), .B2(new_n722), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n474), .A2(new_n722), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n512), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT95), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n505), .B1(new_n510), .B2(new_n511), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n725), .ZN(new_n729));
  AND3_X1   g0529(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n727), .B1(new_n726), .B2(new_n729), .ZN(new_n731));
  OAI211_X1 g0531(.A(G330), .B(new_n724), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n728), .A2(new_n613), .A3(new_n596), .A4(new_n722), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n603), .A2(new_n611), .A3(new_n722), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n732), .A2(new_n735), .ZN(G399));
  INV_X1    g0536(.A(new_n213), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G41), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n225), .A2(new_n205), .A3(new_n206), .A4(new_n454), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT96), .ZN(new_n740));
  OR3_X1    g0540(.A1(new_n738), .A2(new_n209), .A3(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT97), .ZN(new_n742));
  INV_X1    g0542(.A(new_n738), .ZN(new_n743));
  OAI22_X1  g0543(.A1(new_n741), .A2(new_n742), .B1(new_n217), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n744), .B1(new_n742), .B2(new_n741), .ZN(new_n745));
  XOR2_X1   g0545(.A(new_n745), .B(KEYINPUT28), .Z(new_n746));
  INV_X1    g0546(.A(new_n683), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n563), .A2(KEYINPUT100), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT100), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n697), .A2(new_n749), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n505), .B(new_n613), .C1(new_n510), .C2(new_n511), .ZN(new_n751));
  AND4_X1   g0551(.A1(new_n747), .A2(new_n748), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n705), .A2(new_n678), .A3(new_n682), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(KEYINPUT26), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n705), .A2(new_n709), .A3(new_n706), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT99), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n678), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n689), .A2(KEYINPUT99), .A3(new_n648), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n754), .A2(new_n755), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n722), .B1(new_n752), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(KEYINPUT29), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n721), .B1(new_n703), .B2(new_n711), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT29), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n563), .A2(new_n652), .ZN(new_n766));
  INV_X1    g0566(.A(new_n512), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n766), .A2(new_n767), .A3(new_n722), .ZN(new_n768));
  INV_X1    g0568(.A(new_n586), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n769), .A2(new_n606), .A3(new_n310), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n770), .A2(new_n637), .A3(new_n633), .A4(new_n642), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n506), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n772), .A2(new_n532), .A3(new_n541), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT30), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n772), .A2(new_n532), .A3(KEYINPUT30), .A4(new_n541), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n593), .A2(new_n310), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n543), .A2(new_n506), .A3(new_n674), .A4(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n779), .A2(KEYINPUT31), .A3(new_n721), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT98), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n779), .A2(KEYINPUT98), .A3(KEYINPUT31), .A4(new_n721), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n779), .A2(new_n721), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT31), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n768), .A2(new_n782), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G330), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n762), .A2(new_n765), .A3(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n746), .B1(new_n790), .B2(G1), .ZN(G364));
  OAI21_X1  g0591(.A(G330), .B1(new_n730), .B2(new_n731), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n272), .A2(G20), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n209), .B1(new_n793), .B2(G45), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n738), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n792), .A2(new_n797), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n730), .A2(new_n731), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(G330), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n210), .A2(new_n310), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n801), .A2(G190), .A3(new_n319), .ZN(new_n802));
  INV_X1    g0602(.A(G322), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(G190), .A2(G200), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G311), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n363), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n210), .A2(G179), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n805), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n804), .B(new_n808), .C1(G329), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n801), .A2(G200), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n317), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G326), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n813), .A2(G190), .ZN(new_n816));
  XNOR2_X1  g0616(.A(KEYINPUT33), .B(G317), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n809), .A2(G190), .A3(G200), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n816), .A2(new_n817), .B1(new_n819), .B2(G303), .ZN(new_n820));
  NOR3_X1   g0620(.A1(new_n317), .A2(G179), .A3(G200), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n210), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n809), .A2(new_n317), .A3(G200), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n823), .A2(G294), .B1(new_n825), .B2(G283), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n812), .A2(new_n815), .A3(new_n820), .A4(new_n826), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n802), .A2(new_n229), .B1(new_n806), .B2(new_n289), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT102), .Z(new_n829));
  AOI21_X1  g0629(.A(new_n363), .B1(new_n823), .B2(G97), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n825), .A2(G107), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n819), .A2(G87), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n829), .A2(new_n830), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n811), .A2(G159), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n834), .A2(KEYINPUT32), .B1(new_n816), .B2(G68), .ZN(new_n835));
  INV_X1    g0635(.A(new_n814), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n835), .B1(KEYINPUT32), .B2(new_n834), .C1(new_n202), .C2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n827), .B1(new_n833), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n219), .B1(G20), .B2(new_n279), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n251), .A2(new_n304), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n737), .A2(new_n286), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n841), .B(new_n843), .C1(new_n304), .C2(new_n218), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n737), .A2(new_n363), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(G355), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(G116), .B2(new_n213), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n844), .B1(KEYINPUT101), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(KEYINPUT101), .B2(new_n847), .ZN(new_n849));
  NOR2_X1   g0649(.A1(G13), .A2(G33), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n851), .A2(G20), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n852), .A2(new_n839), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n797), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n852), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n840), .B(new_n854), .C1(new_n799), .C2(new_n855), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n800), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(G396));
  NAND4_X1  g0658(.A1(new_n347), .A2(new_n335), .A3(new_n348), .A4(new_n722), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n335), .A2(new_n721), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n346), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n860), .B1(new_n862), .B2(new_n349), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n763), .B(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n796), .B1(new_n864), .B2(new_n788), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n788), .B2(new_n864), .ZN(new_n866));
  INV_X1    g0666(.A(new_n802), .ZN(new_n867));
  INV_X1    g0667(.A(new_n806), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n867), .A2(G143), .B1(new_n868), .B2(G159), .ZN(new_n869));
  INV_X1    g0669(.A(new_n816), .ZN(new_n870));
  INV_X1    g0670(.A(G137), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n869), .B1(new_n870), .B2(new_n264), .C1(new_n871), .C2(new_n836), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT34), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n872), .A2(new_n873), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n825), .A2(G68), .ZN(new_n876));
  INV_X1    g0676(.A(G132), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n876), .B(new_n286), .C1(new_n877), .C2(new_n810), .ZN(new_n878));
  OAI22_X1  g0678(.A1(new_n822), .A2(new_n229), .B1(new_n818), .B2(new_n202), .ZN(new_n879));
  NOR4_X1   g0679(.A1(new_n874), .A2(new_n875), .A3(new_n878), .A4(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(G303), .ZN(new_n881));
  OAI22_X1  g0681(.A1(new_n836), .A2(new_n881), .B1(new_n818), .B2(new_n206), .ZN(new_n882));
  XOR2_X1   g0682(.A(KEYINPUT103), .B(G283), .Z(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  AOI22_X1  g0684(.A1(G97), .A2(new_n823), .B1(new_n816), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n286), .B1(new_n867), .B2(G294), .ZN(new_n886));
  AOI22_X1  g0686(.A1(G116), .A2(new_n868), .B1(new_n811), .B2(G311), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n882), .B(new_n888), .C1(G87), .C2(new_n825), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n839), .B1(new_n880), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n839), .A2(new_n850), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n797), .B1(new_n289), .B2(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n890), .B(new_n892), .C1(new_n863), .C2(new_n851), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n866), .A2(new_n893), .ZN(G384));
  INV_X1    g0694(.A(new_n548), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n895), .A2(KEYINPUT35), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(KEYINPUT35), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n896), .A2(G116), .A3(new_n220), .A4(new_n897), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n898), .B(KEYINPUT36), .Z(new_n899));
  OAI211_X1 g0699(.A(new_n218), .B(G77), .C1(new_n229), .C2(new_n223), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n209), .B(G13), .C1(new_n900), .C2(new_n247), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n666), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n747), .A2(new_n748), .A3(new_n750), .A4(new_n751), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n904), .A2(new_n754), .A3(new_n755), .A4(new_n759), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n764), .B1(new_n905), .B2(new_n722), .ZN(new_n906));
  AOI211_X1 g0706(.A(KEYINPUT29), .B(new_n721), .C1(new_n703), .C2(new_n711), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n452), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT104), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n762), .A2(new_n765), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(KEYINPUT104), .A3(new_n452), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n903), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n444), .A2(new_n722), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n402), .A2(new_n405), .ZN(new_n916));
  INV_X1    g0716(.A(new_n719), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n402), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n916), .A2(new_n918), .A3(new_n398), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(KEYINPUT37), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT37), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n916), .A2(new_n918), .A3(new_n921), .A4(new_n398), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n918), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n407), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT38), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n923), .A2(new_n925), .A3(KEYINPUT38), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n928), .A2(KEYINPUT39), .A3(new_n929), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n923), .A2(new_n925), .A3(KEYINPUT38), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n661), .A2(new_n655), .A3(new_n662), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n924), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n923), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n931), .B1(new_n934), .B2(new_n927), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n915), .B(new_n930), .C1(new_n935), .C2(KEYINPUT39), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n661), .A2(new_n662), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n719), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n928), .A2(new_n929), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n860), .B1(new_n763), .B2(new_n863), .ZN(new_n941));
  INV_X1    g0741(.A(new_n449), .ZN(new_n942));
  INV_X1    g0742(.A(new_n443), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n721), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n942), .B(new_n944), .C1(new_n432), .C2(new_n443), .ZN(new_n945));
  AND3_X1   g0745(.A1(new_n427), .A2(KEYINPUT72), .A3(new_n428), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n419), .B(new_n421), .C1(new_n946), .C2(new_n429), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n943), .B(new_n721), .C1(new_n947), .C2(new_n449), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n941), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n939), .B1(new_n940), .B2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n913), .B(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(G330), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n768), .A2(new_n780), .A3(new_n786), .ZN(new_n955));
  INV_X1    g0755(.A(new_n861), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(new_n344), .B2(new_n345), .ZN(new_n957));
  AND3_X1   g0757(.A1(new_n347), .A2(new_n335), .A3(new_n348), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n859), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(new_n945), .B2(new_n948), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n955), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(KEYINPUT40), .B1(new_n961), .B2(new_n935), .ZN(new_n962));
  AOI21_X1  g0762(.A(KEYINPUT40), .B1(new_n928), .B2(new_n929), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n963), .A2(new_n955), .A3(new_n960), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(KEYINPUT31), .B1(new_n779), .B2(new_n721), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(new_n653), .B2(new_n722), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n451), .B1(new_n780), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n954), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n968), .B2(new_n965), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n953), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n209), .B2(new_n793), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n953), .A2(new_n970), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n902), .B1(new_n972), .B2(new_n973), .ZN(G367));
  OAI21_X1  g0774(.A(new_n690), .B1(new_n626), .B2(new_n722), .ZN(new_n975));
  OR3_X1    g0775(.A1(new_n678), .A2(new_n626), .A3(new_n722), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n852), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n853), .B1(new_n213), .B2(new_n328), .C1(new_n843), .C2(new_n242), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n796), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n870), .A2(new_n394), .B1(new_n824), .B2(new_n289), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(G58), .B2(new_n819), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n802), .A2(new_n264), .B1(new_n806), .B2(new_n202), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n363), .B(new_n984), .C1(G137), .C2(new_n811), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n822), .A2(new_n223), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(G143), .B2(new_n814), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n983), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n823), .A2(G107), .B1(new_n884), .B2(new_n868), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n990), .A2(KEYINPUT109), .ZN(new_n991));
  INV_X1    g0791(.A(G294), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n870), .A2(new_n992), .B1(new_n824), .B2(new_n205), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(G311), .B2(new_n814), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n990), .A2(KEYINPUT109), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n991), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n819), .A2(KEYINPUT46), .A3(G116), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n286), .B1(new_n811), .B2(G317), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n867), .A2(G303), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT46), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n818), .B2(new_n454), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n997), .A2(new_n998), .A3(new_n999), .A4(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n988), .B1(new_n996), .B2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT47), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n981), .B1(new_n1004), .B2(new_n839), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n979), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n557), .A2(new_n721), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n748), .A2(new_n750), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n705), .A2(new_n721), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(KEYINPUT105), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT105), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n705), .A2(new_n1011), .A3(new_n721), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1008), .A2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g0814(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n1015));
  AND3_X1   g0815(.A1(new_n1014), .A2(new_n735), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1015), .B1(new_n1014), .B2(new_n735), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT44), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n1014), .B2(new_n735), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n733), .A2(new_n734), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1021), .A2(new_n1008), .A3(KEYINPUT44), .A4(new_n1013), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1018), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n732), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1018), .A2(new_n732), .A3(new_n1023), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n728), .A2(new_n722), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1029), .A2(new_n724), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n733), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n792), .B(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n790), .B1(new_n1028), .B2(new_n1032), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n738), .B(KEYINPUT41), .Z(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n795), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n977), .A2(KEYINPUT43), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT43), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n978), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n705), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1008), .A2(new_n1013), .ZN(new_n1041));
  OAI211_X1 g0841(.A(KEYINPUT106), .B(new_n1040), .C1(new_n1041), .C2(new_n613), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT106), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n613), .B1(new_n1008), .B2(new_n1013), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1043), .B1(new_n1044), .B2(new_n705), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1042), .A2(new_n722), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n733), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1014), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT42), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1048), .B(new_n1049), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1037), .B(new_n1039), .C1(new_n1046), .C2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1046), .A2(new_n1050), .A3(new_n1038), .A4(new_n978), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n1051), .A2(new_n1053), .B1(new_n732), .B2(new_n1041), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1046), .A2(new_n1050), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1037), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1039), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n732), .A2(new_n1041), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1058), .A2(new_n1059), .A3(new_n1052), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1054), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT108), .ZN(new_n1062));
  NOR3_X1   g0862(.A1(new_n1036), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  AND3_X1   g0863(.A1(new_n1018), .A2(new_n732), .A3(new_n1023), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n732), .B1(new_n1018), .B2(new_n1023), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1032), .A2(new_n789), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n789), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n794), .B1(new_n1068), .B2(new_n1034), .ZN(new_n1069));
  AND3_X1   g0869(.A1(new_n1058), .A2(new_n1059), .A3(new_n1052), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1059), .B1(new_n1058), .B2(new_n1052), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(KEYINPUT108), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1006), .B1(new_n1063), .B2(new_n1073), .ZN(G387));
  OR2_X1    g0874(.A1(new_n239), .A2(new_n304), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1075), .A2(new_n842), .B1(new_n740), .B2(new_n845), .ZN(new_n1076));
  OAI21_X1  g0876(.A(KEYINPUT50), .B1(new_n259), .B2(G50), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1077), .B(new_n304), .C1(new_n223), .C2(new_n289), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n259), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n1078), .A2(new_n740), .A3(new_n1079), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n1076), .A2(new_n1080), .B1(G107), .B2(new_n213), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n797), .B1(new_n1081), .B2(new_n853), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n724), .B2(new_n855), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n806), .A2(new_n223), .B1(new_n810), .B2(new_n264), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n363), .B(new_n1084), .C1(G50), .C2(new_n867), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n819), .A2(G77), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n614), .A2(new_n823), .B1(new_n816), .B2(new_n332), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n814), .A2(G159), .B1(new_n825), .B2(G97), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n286), .B1(new_n811), .B2(G326), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n822), .A2(new_n883), .B1(new_n818), .B2(new_n992), .ZN(new_n1091));
  INV_X1    g0891(.A(G317), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n802), .A2(new_n1092), .B1(new_n806), .B2(new_n881), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT110), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(G311), .A2(new_n816), .B1(new_n814), .B2(G322), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1091), .B1(new_n1098), .B2(KEYINPUT48), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT111), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(KEYINPUT48), .B2(new_n1098), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT112), .Z(new_n1102));
  INV_X1    g0902(.A(KEYINPUT49), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1090), .B1(new_n454), .B2(new_n824), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1089), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1083), .B1(new_n1106), .B2(new_n839), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1030), .A2(new_n733), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n792), .B(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1107), .B1(new_n795), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1032), .A2(new_n789), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n790), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1111), .A2(new_n1112), .A3(new_n738), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1110), .A2(new_n1113), .ZN(G393));
  NAND2_X1  g0914(.A1(new_n1041), .A2(new_n852), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT113), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n842), .A2(new_n246), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n852), .B(new_n839), .C1(new_n737), .C2(G97), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n797), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n839), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n836), .A2(new_n264), .B1(new_n394), .B2(new_n802), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT51), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n870), .A2(new_n202), .B1(new_n824), .B2(new_n225), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n363), .B1(new_n811), .B2(G143), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n259), .B2(new_n806), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n822), .A2(new_n289), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n818), .A2(new_n223), .ZN(new_n1127));
  NOR4_X1   g0927(.A1(new_n1123), .A2(new_n1125), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n836), .A2(new_n1092), .B1(new_n807), .B2(new_n802), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT52), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n870), .A2(new_n881), .B1(new_n454), .B2(new_n822), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n831), .B1(new_n818), .B2(new_n883), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n363), .B1(new_n810), .B2(new_n803), .C1(new_n992), .C2(new_n806), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1122), .A2(new_n1128), .B1(new_n1130), .B2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1116), .B(new_n1119), .C1(new_n1120), .C2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n1028), .B2(new_n794), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT114), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1028), .A2(KEYINPUT114), .A3(new_n1112), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n743), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1137), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(G390));
  OAI21_X1  g0944(.A(new_n914), .B1(new_n941), .B2(new_n950), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n930), .B1(new_n935), .B2(KEYINPUT39), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n787), .A2(G330), .A3(new_n863), .A4(new_n949), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT116), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1148), .B(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n862), .A2(new_n349), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n722), .B(new_n1151), .C1(new_n752), .C2(new_n760), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n859), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n949), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n932), .A2(new_n924), .B1(new_n920), .B2(new_n922), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n929), .B1(new_n1155), .B2(KEYINPUT38), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n914), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(KEYINPUT115), .B1(new_n1154), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n950), .B1(new_n1152), .B2(new_n859), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT115), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n1160), .A2(new_n1161), .A3(new_n1157), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1147), .B(new_n1150), .C1(new_n1159), .C2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1154), .A2(KEYINPUT115), .A3(new_n1158), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1161), .B1(new_n1160), .B2(new_n1157), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n1164), .A2(new_n1165), .B1(new_n1146), .B2(new_n1145), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n955), .A2(G330), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n960), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1163), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1170), .A2(new_n794), .ZN(new_n1171));
  INV_X1    g0971(.A(G283), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n836), .A2(new_n1172), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1126), .B(new_n1173), .C1(G107), .C2(new_n816), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n802), .A2(new_n454), .B1(new_n810), .B2(new_n992), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n286), .B(new_n1175), .C1(G97), .C2(new_n868), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1174), .A2(new_n832), .A3(new_n876), .A4(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n286), .B1(new_n824), .B2(new_n202), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT117), .Z(new_n1179));
  OAI22_X1  g0979(.A1(new_n870), .A2(new_n871), .B1(new_n394), .B2(new_n822), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(G128), .B2(new_n814), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n818), .A2(new_n264), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT53), .ZN(new_n1183));
  INV_X1    g0983(.A(G125), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n802), .A2(new_n877), .B1(new_n810), .B2(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(KEYINPUT54), .B(G143), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1185), .B1(new_n868), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1181), .A2(new_n1183), .A3(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1177), .B1(new_n1179), .B2(new_n1189), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1190), .A2(new_n839), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n891), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n796), .B1(new_n332), .B2(new_n1192), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1191), .B(new_n1193), .C1(new_n1146), .C2(new_n850), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1171), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n452), .A2(new_n1168), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT104), .B1(new_n911), .B2(new_n452), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n909), .B(new_n451), .C1(new_n762), .C2(new_n765), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n666), .B(new_n1196), .C1(new_n1197), .C2(new_n1198), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1152), .A2(new_n859), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n950), .B1(new_n1167), .B2(new_n959), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n712), .A2(new_n722), .A3(new_n863), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n859), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n950), .B1(new_n788), .B2(new_n959), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n1169), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1150), .A2(new_n1202), .B1(new_n1204), .B2(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1199), .A2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1147), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1209), .A2(new_n960), .A3(new_n1168), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1208), .A2(new_n1210), .A3(new_n1163), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1206), .A2(new_n1204), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1148), .B(KEYINPUT116), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1212), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1215), .A2(new_n913), .A3(new_n1196), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1170), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1211), .A2(new_n1217), .A3(new_n738), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1195), .A2(new_n1218), .ZN(G378));
  NOR2_X1   g1019(.A1(new_n278), .A2(new_n719), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n355), .A2(new_n1220), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n312), .B1(new_n278), .B2(new_n719), .C1(new_n354), .C2(new_n323), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1223), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n850), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n363), .A2(new_n303), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G283), .B2(new_n811), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1229), .B(new_n1086), .C1(new_n229), .C2(new_n824), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT118), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n802), .A2(new_n206), .B1(new_n806), .B2(new_n328), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n205), .A2(new_n870), .B1(new_n836), .B2(new_n454), .ZN(new_n1233));
  NOR4_X1   g1033(.A1(new_n1231), .A2(new_n986), .A3(new_n1232), .A4(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(G50), .B1(new_n254), .B2(new_n303), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1234), .A2(KEYINPUT58), .B1(new_n1228), .B2(new_n1235), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n1184), .A2(new_n836), .B1(new_n870), .B2(new_n877), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n867), .A2(G128), .B1(new_n868), .B2(G137), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n818), .B2(new_n1186), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1237), .B(new_n1239), .C1(G150), .C2(new_n823), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(KEYINPUT59), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n825), .A2(G159), .ZN(new_n1243));
  AOI211_X1 g1043(.A(G33), .B(G41), .C1(new_n811), .C2(G124), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1241), .A2(KEYINPUT59), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n1236), .B1(KEYINPUT58), .B2(new_n1234), .C1(new_n1245), .C2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n839), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n797), .B1(new_n202), .B2(new_n891), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1227), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1204), .A2(new_n940), .A3(new_n949), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1252), .A2(new_n938), .A3(new_n936), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1226), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n965), .B2(G330), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n954), .B(new_n1226), .C1(new_n962), .C2(new_n964), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1253), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1156), .A2(new_n955), .A3(new_n960), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n949), .A2(new_n863), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n780), .B2(new_n967), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(KEYINPUT40), .A2(new_n1258), .B1(new_n1260), .B2(new_n963), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1226), .B1(new_n1261), .B2(new_n954), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n965), .A2(G330), .A3(new_n1254), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n952), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT119), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1257), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(KEYINPUT119), .A3(new_n1253), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1251), .B1(new_n1269), .B2(new_n795), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT121), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1257), .A2(new_n1271), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1253), .B(KEYINPUT121), .C1(new_n1255), .C2(new_n1256), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT120), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1274), .B1(new_n1275), .B2(new_n952), .ZN(new_n1276));
  AND4_X1   g1076(.A1(new_n1274), .A2(new_n952), .A3(new_n1262), .A4(new_n1263), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1272), .B(new_n1273), .C1(new_n1276), .C2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1199), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n1170), .B2(new_n1216), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1278), .A2(new_n1280), .A3(KEYINPUT57), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n738), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT57), .B1(new_n1269), .B2(new_n1280), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1270), .B1(new_n1282), .B2(new_n1283), .ZN(G375));
  NOR2_X1   g1084(.A1(new_n1207), .A2(new_n794), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n949), .A2(new_n851), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(new_n1286), .B(KEYINPUT122), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(G107), .A2(new_n868), .B1(new_n811), .B2(G303), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1288), .B1(new_n1172), .B2(new_n802), .ZN(new_n1289));
  OAI22_X1  g1089(.A1(new_n870), .A2(new_n454), .B1(new_n328), .B2(new_n822), .ZN(new_n1290));
  OAI22_X1  g1090(.A1(new_n836), .A2(new_n992), .B1(new_n818), .B2(new_n205), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1289), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n363), .B1(new_n824), .B2(new_n289), .ZN(new_n1293));
  XOR2_X1   g1093(.A(new_n1293), .B(KEYINPUT123), .Z(new_n1294));
  AOI21_X1  g1094(.A(new_n363), .B1(new_n811), .B2(G128), .ZN(new_n1295));
  OAI221_X1 g1095(.A(new_n1295), .B1(new_n871), .B2(new_n802), .C1(new_n264), .C2(new_n806), .ZN(new_n1296));
  OAI22_X1  g1096(.A1(new_n870), .A2(new_n1186), .B1(new_n824), .B2(new_n229), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  OAI22_X1  g1098(.A1(new_n822), .A2(new_n202), .B1(new_n818), .B2(new_n394), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1299), .B1(G132), .B2(new_n814), .ZN(new_n1300));
  AOI22_X1  g1100(.A1(new_n1292), .A2(new_n1294), .B1(new_n1298), .B2(new_n1300), .ZN(new_n1301));
  OAI221_X1 g1101(.A(new_n796), .B1(G68), .B2(new_n1192), .C1(new_n1301), .C2(new_n1120), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1287), .A2(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(KEYINPUT124), .B1(new_n1285), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1215), .A2(new_n795), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT124), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1303), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1305), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1304), .A2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1199), .A2(new_n1207), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1216), .A2(new_n1310), .A3(new_n1035), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1309), .A2(new_n1311), .ZN(G381));
  NAND2_X1  g1112(.A1(new_n1269), .A2(new_n795), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1250), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT57), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1273), .ZN(new_n1316));
  AOI21_X1  g1116(.A(KEYINPUT121), .B1(new_n1267), .B2(new_n1253), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1275), .A2(new_n1274), .A3(new_n952), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1264), .A2(KEYINPUT120), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1315), .B1(new_n1318), .B2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n743), .B1(new_n1322), .B2(new_n1280), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1283), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1314), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1110), .A2(new_n857), .A3(new_n1113), .ZN(new_n1326));
  NOR4_X1   g1126(.A1(G381), .A2(G390), .A3(G384), .A4(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1006), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1062), .B1(new_n1036), .B2(new_n1061), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1069), .A2(new_n1072), .A3(KEYINPUT108), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1328), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(G378), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1325), .A2(new_n1327), .A3(new_n1331), .A4(new_n1332), .ZN(G407));
  INV_X1    g1133(.A(G213), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1334), .A2(G343), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1325), .A2(new_n1332), .A3(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(G407), .A2(G213), .A3(new_n1336), .ZN(new_n1337));
  XNOR2_X1  g1137(.A(new_n1337), .B(KEYINPUT125), .ZN(G409));
  XOR2_X1   g1138(.A(KEYINPUT126), .B(KEYINPUT60), .Z(new_n1339));
  NAND2_X1  g1139(.A1(new_n1310), .A2(new_n1339), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1199), .A2(new_n1207), .A3(KEYINPUT60), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1340), .A2(new_n738), .A3(new_n1216), .A4(new_n1341), .ZN(new_n1342));
  AND3_X1   g1142(.A1(new_n1342), .A2(new_n1309), .A3(G384), .ZN(new_n1343));
  AOI21_X1  g1143(.A(G384), .B1(new_n1342), .B2(new_n1309), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1335), .A2(G2897), .ZN(new_n1345));
  NOR3_X1   g1145(.A1(new_n1343), .A2(new_n1344), .A3(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1345), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1340), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1341), .A2(new_n1216), .A3(new_n738), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1306), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1350));
  AOI211_X1 g1150(.A(KEYINPUT124), .B(new_n1303), .C1(new_n1215), .C2(new_n795), .ZN(new_n1351));
  OAI22_X1  g1151(.A1(new_n1348), .A2(new_n1349), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(G384), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1352), .A2(new_n1353), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1342), .A2(new_n1309), .A3(G384), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1347), .B1(new_n1354), .B2(new_n1355), .ZN(new_n1356));
  NOR2_X1   g1156(.A1(new_n1346), .A2(new_n1356), .ZN(new_n1357));
  OAI211_X1 g1157(.A(G378), .B(new_n1270), .C1(new_n1282), .C2(new_n1283), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1251), .B1(new_n1278), .B2(new_n795), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1269), .A2(new_n1280), .A3(new_n1035), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1359), .A2(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1332), .A2(new_n1361), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n1335), .B1(new_n1358), .B2(new_n1362), .ZN(new_n1363));
  AOI21_X1  g1163(.A(new_n1357), .B1(new_n1363), .B2(KEYINPUT127), .ZN(new_n1364));
  INV_X1    g1164(.A(KEYINPUT127), .ZN(new_n1365));
  AOI21_X1  g1165(.A(G378), .B1(new_n1360), .B2(new_n1359), .ZN(new_n1366));
  AOI21_X1  g1166(.A(new_n1366), .B1(new_n1325), .B2(G378), .ZN(new_n1367));
  OAI21_X1  g1167(.A(new_n1365), .B1(new_n1367), .B2(new_n1335), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1364), .A2(new_n1368), .ZN(new_n1369));
  NOR2_X1   g1169(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1363), .A2(KEYINPUT63), .A3(new_n1370), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(G393), .A2(G396), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1372), .A2(new_n1326), .ZN(new_n1373));
  NOR2_X1   g1173(.A1(new_n1331), .A2(G390), .ZN(new_n1374));
  AOI211_X1 g1174(.A(new_n1328), .B(new_n1143), .C1(new_n1329), .C2(new_n1330), .ZN(new_n1375));
  OAI21_X1  g1175(.A(new_n1373), .B1(new_n1374), .B2(new_n1375), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(G387), .A2(new_n1143), .ZN(new_n1377));
  INV_X1    g1177(.A(new_n1373), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1331), .A2(G390), .ZN(new_n1379));
  NAND3_X1  g1179(.A1(new_n1377), .A2(new_n1378), .A3(new_n1379), .ZN(new_n1380));
  INV_X1    g1180(.A(KEYINPUT61), .ZN(new_n1381));
  NAND3_X1  g1181(.A1(new_n1376), .A2(new_n1380), .A3(new_n1381), .ZN(new_n1382));
  NAND2_X1  g1182(.A1(new_n1358), .A2(new_n1362), .ZN(new_n1383));
  INV_X1    g1183(.A(new_n1335), .ZN(new_n1384));
  NAND3_X1  g1184(.A1(new_n1383), .A2(new_n1384), .A3(new_n1370), .ZN(new_n1385));
  INV_X1    g1185(.A(KEYINPUT63), .ZN(new_n1386));
  AOI21_X1  g1186(.A(new_n1382), .B1(new_n1385), .B2(new_n1386), .ZN(new_n1387));
  NAND3_X1  g1187(.A1(new_n1369), .A2(new_n1371), .A3(new_n1387), .ZN(new_n1388));
  INV_X1    g1188(.A(KEYINPUT62), .ZN(new_n1389));
  AND3_X1   g1189(.A1(new_n1363), .A2(new_n1389), .A3(new_n1370), .ZN(new_n1390));
  OAI21_X1  g1190(.A(new_n1381), .B1(new_n1363), .B2(new_n1357), .ZN(new_n1391));
  AOI21_X1  g1191(.A(new_n1389), .B1(new_n1363), .B2(new_n1370), .ZN(new_n1392));
  NOR3_X1   g1192(.A1(new_n1390), .A2(new_n1391), .A3(new_n1392), .ZN(new_n1393));
  NAND2_X1  g1193(.A1(new_n1376), .A2(new_n1380), .ZN(new_n1394));
  INV_X1    g1194(.A(new_n1394), .ZN(new_n1395));
  OAI21_X1  g1195(.A(new_n1388), .B1(new_n1393), .B2(new_n1395), .ZN(G405));
  NAND2_X1  g1196(.A1(G375), .A2(new_n1332), .ZN(new_n1397));
  NAND2_X1  g1197(.A1(new_n1397), .A2(new_n1358), .ZN(new_n1398));
  NAND2_X1  g1198(.A1(new_n1398), .A2(new_n1370), .ZN(new_n1399));
  OAI211_X1 g1199(.A(new_n1397), .B(new_n1358), .C1(new_n1344), .C2(new_n1343), .ZN(new_n1400));
  NAND2_X1  g1200(.A1(new_n1399), .A2(new_n1400), .ZN(new_n1401));
  XNOR2_X1  g1201(.A(new_n1401), .B(new_n1394), .ZN(G402));
endmodule


