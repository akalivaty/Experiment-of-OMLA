//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 0 0 1 1 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 1 1 1 0 1 0 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1274, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT0), .Z(new_n208));
  AOI22_X1  g0008(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n209));
  INV_X1    g0009(.A(G58), .ZN(new_n210));
  INV_X1    g0010(.A(G232), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n205), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT1), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g0022(.A1(G58), .A2(G68), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT64), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n225), .A2(G50), .A3(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  AOI211_X1 g0028(.A(new_n208), .B(new_n219), .C1(new_n222), .C2(new_n228), .ZN(G361));
  XOR2_X1   g0029(.A(G226), .B(G232), .Z(new_n230));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XNOR2_X1  g0038(.A(G68), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT66), .ZN(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(G97), .B(G107), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  INV_X1    g0046(.A(G1), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n247), .B1(G41), .B2(G45), .ZN(new_n248));
  INV_X1    g0048(.A(G274), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  OAI211_X1 g0052(.A(G1), .B(G13), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n248), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  AND2_X1   g0055(.A1(new_n255), .A2(G244), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n220), .B1(G33), .B2(G41), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT3), .B(G33), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(G232), .A3(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n258), .A2(G238), .A3(G1698), .ZN(new_n261));
  INV_X1    g0061(.A(G107), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n260), .B(new_n261), .C1(new_n262), .C2(new_n258), .ZN(new_n263));
  AOI211_X1 g0063(.A(new_n250), .B(new_n256), .C1(new_n257), .C2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G179), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XOR2_X1   g0066(.A(KEYINPUT8), .B(G58), .Z(new_n267));
  NOR2_X1   g0067(.A1(G20), .A2(G33), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n267), .A2(new_n268), .B1(G20), .B2(G77), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n221), .A2(G33), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT15), .B(G87), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n220), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n274), .B1(new_n247), .B2(G20), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G77), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n247), .A2(G13), .A3(G20), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n275), .B(new_n277), .C1(G77), .C2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n279), .B1(new_n264), .B2(G169), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n266), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G200), .ZN(new_n282));
  OR2_X1    g0082(.A1(new_n264), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n279), .B1(G190), .B2(new_n264), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n281), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n258), .A2(G232), .A3(G1698), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n258), .A2(G226), .A3(new_n259), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G97), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n257), .ZN(new_n290));
  INV_X1    g0090(.A(new_n250), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n291), .B1(new_n254), .B2(new_n213), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT68), .B(KEYINPUT13), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  AND3_X1   g0095(.A1(new_n290), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n295), .B1(new_n290), .B2(new_n293), .ZN(new_n297));
  OAI21_X1  g0097(.A(G169), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT14), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n290), .A2(new_n293), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT69), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n300), .A2(new_n301), .A3(KEYINPUT13), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n292), .B1(new_n289), .B2(new_n257), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT13), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT69), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n295), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n302), .A2(new_n305), .A3(G179), .A4(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT14), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n308), .B(G169), .C1(new_n296), .C2(new_n297), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n299), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n278), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n212), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n312), .B(KEYINPUT12), .ZN(new_n313));
  INV_X1    g0113(.A(new_n276), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT11), .ZN(new_n315));
  INV_X1    g0115(.A(new_n268), .ZN(new_n316));
  INV_X1    g0116(.A(G50), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n270), .A2(new_n202), .B1(new_n221), .B2(G68), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n274), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI221_X1 g0120(.A(new_n313), .B1(new_n212), .B2(new_n314), .C1(new_n315), .C2(new_n320), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n320), .A2(new_n315), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n310), .A2(new_n324), .ZN(new_n325));
  AND4_X1   g0125(.A1(G190), .A2(new_n302), .A3(new_n305), .A4(new_n306), .ZN(new_n326));
  OAI21_X1  g0126(.A(G200), .B1(new_n296), .B2(new_n297), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n323), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n267), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(new_n270), .ZN(new_n331));
  INV_X1    g0131(.A(G150), .ZN(new_n332));
  OAI22_X1  g0132(.A1(new_n332), .A2(new_n316), .B1(new_n201), .B2(new_n221), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n274), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n278), .A2(G50), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n335), .B1(new_n276), .B2(G50), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n250), .B1(new_n255), .B2(G226), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT3), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G33), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n202), .ZN(new_n343));
  MUX2_X1   g0143(.A(G222), .B(G223), .S(G1698), .Z(new_n344));
  OAI211_X1 g0144(.A(new_n343), .B(new_n257), .C1(new_n342), .C2(new_n344), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n338), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n337), .B1(new_n346), .B2(G169), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n347), .B1(new_n265), .B2(new_n346), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n346), .A2(new_n282), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(G190), .B2(new_n346), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n337), .B(KEYINPUT9), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT10), .B1(new_n349), .B2(KEYINPUT67), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n350), .A2(new_n351), .A3(new_n353), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n348), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n285), .A2(new_n325), .A3(new_n329), .A4(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n267), .A2(new_n311), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n359), .B1(new_n314), .B2(new_n267), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT16), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT7), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(new_n258), .B2(G20), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n342), .A2(KEYINPUT7), .A3(new_n221), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n212), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n210), .A2(new_n212), .ZN(new_n366));
  OAI21_X1  g0166(.A(G20), .B1(new_n366), .B2(new_n223), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n268), .A2(G159), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI211_X1 g0169(.A(KEYINPUT70), .B(new_n361), .C1(new_n365), .C2(new_n369), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n370), .A2(new_n274), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n361), .B1(new_n365), .B2(new_n369), .ZN(new_n372));
  NOR3_X1   g0172(.A1(new_n365), .A2(new_n361), .A3(new_n369), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT70), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n360), .B1(new_n371), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n291), .B1(new_n254), .B2(new_n211), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n339), .A2(new_n341), .A3(G226), .A4(G1698), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n378), .A2(KEYINPUT71), .B1(G33), .B2(G87), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT72), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n258), .A2(new_n380), .A3(G223), .A4(new_n259), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT71), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n258), .A2(new_n382), .A3(G226), .A4(G1698), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n339), .A2(new_n341), .A3(G223), .A4(new_n259), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT72), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n379), .A2(new_n381), .A3(new_n383), .A4(new_n385), .ZN(new_n386));
  AOI211_X1 g0186(.A(new_n265), .B(new_n377), .C1(new_n386), .C2(new_n257), .ZN(new_n387));
  INV_X1    g0187(.A(G169), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n385), .A2(new_n381), .A3(new_n383), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n378), .A2(KEYINPUT71), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G33), .A2(G87), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n257), .B1(new_n389), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n377), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n388), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n387), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT18), .B1(new_n376), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n371), .A2(new_n375), .ZN(new_n398));
  INV_X1    g0198(.A(new_n360), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT18), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n393), .A2(G179), .A3(new_n394), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n377), .B1(new_n386), .B2(new_n257), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n402), .B1(new_n388), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n400), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n282), .B1(new_n393), .B2(new_n394), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n406), .B1(G190), .B2(new_n403), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT17), .ZN(new_n408));
  AND3_X1   g0208(.A1(new_n376), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n408), .B1(new_n376), .B2(new_n407), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n397), .B(new_n405), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n358), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT78), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n340), .A2(G33), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n415));
  OAI21_X1  g0215(.A(G303), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n339), .A2(new_n341), .A3(G257), .A4(new_n259), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n339), .A2(new_n341), .A3(G264), .A4(G1698), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n257), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n252), .A2(KEYINPUT5), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n247), .B(G45), .C1(new_n252), .C2(KEYINPUT5), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n421), .B1(new_n422), .B2(KEYINPUT74), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT74), .ZN(new_n424));
  INV_X1    g0224(.A(G45), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n425), .A2(G1), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT5), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(G41), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n424), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(G270), .B(new_n253), .C1(new_n423), .C2(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n257), .A2(new_n249), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n426), .A2(new_n424), .A3(new_n428), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n422), .A2(KEYINPUT74), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n431), .A2(new_n432), .A3(new_n433), .A4(new_n421), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n420), .A2(new_n430), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(G169), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n278), .A2(G116), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n273), .A2(new_n220), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n247), .A2(G33), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n439), .A2(new_n278), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G116), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n438), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(G33), .A2(G283), .ZN(new_n444));
  INV_X1    g0244(.A(G97), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n444), .B(new_n221), .C1(G33), .C2(new_n445), .ZN(new_n446));
  AOI221_X4 g0246(.A(KEYINPUT76), .B1(new_n442), .B2(G20), .C1(new_n273), .C2(new_n220), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT76), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n442), .A2(G20), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n448), .B1(new_n274), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n446), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT20), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(KEYINPUT20), .B(new_n446), .C1(new_n447), .C2(new_n450), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n443), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n413), .B1(new_n436), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n423), .A2(new_n429), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n457), .A2(new_n431), .B1(new_n419), .B2(new_n257), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n388), .B1(new_n458), .B2(new_n430), .ZN(new_n459));
  INV_X1    g0259(.A(new_n443), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n274), .A2(new_n449), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT76), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n274), .A2(new_n448), .A3(new_n449), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT20), .B1(new_n464), .B2(new_n446), .ZN(new_n465));
  INV_X1    g0265(.A(new_n454), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n459), .A2(new_n467), .A3(KEYINPUT78), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT21), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n456), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT79), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n456), .A2(new_n468), .A3(KEYINPUT79), .A4(new_n469), .ZN(new_n473));
  OAI22_X1  g0273(.A1(new_n436), .A2(new_n469), .B1(new_n265), .B2(new_n435), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n467), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT77), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n474), .A2(KEYINPUT77), .A3(new_n467), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n472), .A2(new_n473), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n435), .A2(G200), .ZN(new_n480));
  INV_X1    g0280(.A(G190), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n480), .B(new_n455), .C1(new_n481), .C2(new_n435), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g0283(.A(G257), .B(new_n253), .C1(new_n423), .C2(new_n429), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n484), .A2(new_n434), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n339), .A2(new_n341), .A3(G244), .A4(new_n259), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT4), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n258), .A2(G250), .A3(G1698), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(new_n444), .A3(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n486), .A2(new_n487), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n257), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n485), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G200), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n485), .A2(new_n492), .A3(G190), .ZN(new_n495));
  NOR3_X1   g0295(.A1(new_n258), .A2(new_n362), .A3(G20), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT7), .B1(new_n342), .B2(new_n221), .ZN(new_n497));
  OAI21_X1  g0297(.A(G107), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n316), .A2(new_n202), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n262), .A2(G97), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n445), .A2(G107), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT6), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n503), .B1(new_n502), .B2(new_n500), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n499), .B1(new_n504), .B2(G20), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n439), .B1(new_n498), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT73), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n278), .A2(G97), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n439), .A2(new_n278), .A3(new_n440), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n508), .B1(new_n509), .B2(G97), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n506), .A2(new_n507), .A3(new_n511), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n502), .A2(new_n445), .A3(G107), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n513), .B1(new_n502), .B2(new_n244), .ZN(new_n514));
  OAI22_X1  g0314(.A1(new_n514), .A2(new_n221), .B1(new_n202), .B2(new_n316), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n262), .B1(new_n363), .B2(new_n364), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n274), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT73), .B1(new_n517), .B2(new_n510), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n494), .B(new_n495), .C1(new_n512), .C2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT75), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n339), .A2(new_n341), .A3(G238), .A4(new_n259), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n339), .A2(new_n341), .A3(G244), .A4(G1698), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n521), .B(new_n522), .C1(new_n251), .C2(new_n442), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n257), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n426), .A2(G274), .ZN(new_n525));
  OAI21_X1  g0325(.A(G250), .B1(new_n425), .B2(G1), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n525), .B1(new_n257), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n520), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  AOI211_X1 g0329(.A(KEYINPUT75), .B(new_n527), .C1(new_n523), .C2(new_n257), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n265), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT19), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n221), .B1(new_n288), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(G87), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n534), .A2(new_n445), .A3(new_n262), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n339), .A2(new_n341), .A3(new_n221), .A4(G68), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n532), .B1(new_n270), .B2(new_n445), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n274), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n271), .A2(new_n311), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n540), .B(new_n541), .C1(new_n271), .C2(new_n441), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n524), .A2(new_n528), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT75), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n524), .A2(new_n520), .A3(new_n528), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n531), .B(new_n542), .C1(new_n546), .C2(G169), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n544), .A2(G200), .A3(new_n545), .ZN(new_n548));
  OAI21_X1  g0348(.A(G190), .B1(new_n529), .B2(new_n530), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n509), .A2(G87), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n540), .A2(new_n550), .A3(new_n541), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n517), .A2(new_n510), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n485), .A2(new_n492), .A3(G179), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n388), .B1(new_n485), .B2(new_n492), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n519), .A2(new_n547), .A3(new_n552), .A4(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n339), .A2(new_n341), .A3(G257), .A4(G1698), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n339), .A2(new_n341), .A3(G250), .A4(new_n259), .ZN(new_n559));
  NAND2_X1  g0359(.A1(G33), .A2(G294), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT81), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n558), .A2(new_n559), .A3(KEYINPUT81), .A4(new_n560), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n563), .A2(new_n257), .A3(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(G264), .B(new_n253), .C1(new_n423), .C2(new_n429), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT82), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n433), .A2(new_n421), .A3(new_n432), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n569), .A2(KEYINPUT82), .A3(G264), .A4(new_n253), .ZN(new_n570));
  AND3_X1   g0370(.A1(new_n565), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n571), .A2(new_n265), .A3(new_n434), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n339), .A2(new_n341), .A3(new_n221), .A4(G87), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT22), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT22), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n258), .A2(new_n575), .A3(new_n221), .A4(G87), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT23), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n221), .B2(G107), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n262), .A2(KEYINPUT23), .A3(G20), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n221), .A2(G33), .A3(G116), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n577), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT24), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n439), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n583), .B1(new_n574), .B2(new_n576), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT24), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n247), .A2(new_n262), .A3(G13), .A4(G20), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT80), .ZN(new_n592));
  XNOR2_X1  g0392(.A(new_n591), .B(new_n592), .ZN(new_n593));
  AOI22_X1  g0393(.A1(KEYINPUT25), .A2(new_n593), .B1(new_n509), .B2(G107), .ZN(new_n594));
  XNOR2_X1  g0394(.A(new_n591), .B(KEYINPUT80), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT25), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n590), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n565), .A2(new_n568), .A3(new_n570), .A4(new_n434), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n388), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n572), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(G200), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n593), .A2(KEYINPUT25), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n597), .B(new_n604), .C1(new_n262), .C2(new_n441), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n605), .B1(new_n587), .B2(new_n589), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n603), .B(new_n606), .C1(new_n481), .C2(new_n600), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n557), .A2(new_n608), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n412), .A2(new_n483), .A3(new_n609), .ZN(G372));
  AOI21_X1  g0410(.A(new_n282), .B1(new_n485), .B2(new_n492), .ZN(new_n611));
  INV_X1    g0411(.A(new_n493), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n611), .B1(new_n612), .B2(G190), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n507), .B1(new_n506), .B2(new_n511), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n517), .A2(KEYINPUT73), .A3(new_n510), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n493), .A2(G169), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n485), .A2(new_n492), .A3(G179), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n613), .A2(new_n616), .B1(new_n619), .B2(new_n553), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n543), .A2(G200), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n621), .A2(KEYINPUT83), .A3(new_n551), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT83), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n282), .B1(new_n524), .B2(new_n528), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n540), .A2(new_n550), .A3(new_n541), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n622), .A2(new_n549), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n543), .A2(new_n388), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n531), .A2(new_n542), .A3(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n620), .A2(new_n630), .A3(new_n607), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n472), .A2(new_n473), .B1(new_n467), .B2(new_n474), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n631), .B1(new_n632), .B2(new_n602), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT26), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n630), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n547), .A2(new_n552), .A3(new_n553), .A4(new_n619), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(KEYINPUT26), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n636), .A2(new_n638), .A3(new_n629), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n412), .B1(new_n633), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT84), .B1(new_n376), .B2(new_n396), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT84), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n370), .A2(new_n274), .ZN(new_n643));
  OAI21_X1  g0443(.A(G68), .B1(new_n496), .B2(new_n497), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n644), .A2(KEYINPUT16), .A3(new_n368), .A4(new_n367), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT70), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n643), .B1(new_n646), .B2(new_n372), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n642), .B(new_n404), .C1(new_n647), .C2(new_n360), .ZN(new_n648));
  XNOR2_X1  g0448(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n641), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n649), .B1(new_n641), .B2(new_n648), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n329), .A2(new_n281), .B1(new_n324), .B2(new_n310), .ZN(new_n653));
  INV_X1    g0453(.A(new_n410), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n376), .A2(new_n407), .A3(new_n408), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n652), .B1(new_n653), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n355), .A2(new_n356), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n348), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n640), .A2(new_n660), .ZN(G369));
  INV_X1    g0461(.A(G213), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n221), .A2(G13), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n247), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n662), .B1(new_n664), .B2(KEYINPUT27), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(KEYINPUT27), .B2(new_n664), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n666), .B(KEYINPUT86), .ZN(new_n667));
  INV_X1    g0467(.A(G343), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(new_n455), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n483), .A2(new_n672), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n632), .A2(new_n672), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G330), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT87), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n669), .A2(new_n599), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n602), .A2(new_n607), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(KEYINPUT88), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n602), .A2(new_n670), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT88), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n602), .A2(new_n607), .A3(new_n682), .A4(new_n678), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n680), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n677), .A2(new_n684), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n680), .A2(new_n681), .A3(new_n683), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n477), .A2(new_n478), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n459), .A2(new_n467), .ZN(new_n688));
  AOI21_X1  g0488(.A(KEYINPUT21), .B1(new_n688), .B2(new_n413), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT79), .B1(new_n689), .B2(new_n468), .ZN(new_n690));
  INV_X1    g0490(.A(new_n473), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n687), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT89), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(new_n693), .A3(new_n670), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT89), .B1(new_n479), .B2(new_n669), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n686), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n602), .A2(new_n669), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT90), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n693), .B1(new_n692), .B2(new_n670), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n479), .A2(KEYINPUT89), .A3(new_n669), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n684), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT90), .ZN(new_n702));
  INV_X1    g0502(.A(new_n697), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n685), .A2(new_n698), .A3(new_n704), .ZN(G399));
  INV_X1    g0505(.A(new_n206), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G41), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n535), .A2(G116), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G1), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n227), .B2(new_n708), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n479), .A2(new_n609), .A3(new_n482), .A4(new_n670), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n435), .A2(new_n265), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n546), .A2(new_n612), .A3(new_n571), .A4(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT30), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n493), .A2(new_n265), .A3(new_n435), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(KEYINPUT30), .A3(new_n571), .A4(new_n546), .ZN(new_n719));
  AOI21_X1  g0519(.A(G179), .B1(new_n524), .B2(new_n528), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n600), .A2(new_n493), .A3(new_n435), .A4(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n717), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT91), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n670), .B1(new_n722), .B2(new_n723), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n713), .A2(KEYINPUT31), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n722), .A2(KEYINPUT31), .A3(new_n669), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G330), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n631), .B1(new_n479), .B2(new_n602), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n627), .A2(new_n629), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n619), .A2(new_n614), .A3(new_n615), .ZN(new_n732));
  OAI21_X1  g0532(.A(KEYINPUT26), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT92), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n629), .B(new_n734), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n733), .B(new_n735), .C1(KEYINPUT26), .C2(new_n637), .ZN(new_n736));
  OAI211_X1 g0536(.A(KEYINPUT29), .B(new_n670), .C1(new_n730), .C2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n631), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n475), .B(new_n602), .C1(new_n690), .C2(new_n691), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AND3_X1   g0540(.A1(new_n636), .A2(new_n638), .A3(new_n629), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n669), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n737), .B1(new_n742), .B2(KEYINPUT29), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n729), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n712), .B1(new_n745), .B2(G1), .ZN(G364));
  INV_X1    g0546(.A(KEYINPUT87), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n676), .B(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n247), .B1(new_n663), .B2(G45), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n707), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n748), .B(new_n752), .C1(G330), .C2(new_n675), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n706), .A2(new_n342), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G355), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(G116), .B2(new_n206), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n242), .A2(G45), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n706), .A2(new_n258), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n759), .B1(new_n228), .B2(new_n425), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n756), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n220), .B1(G20), .B2(new_n388), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n751), .B1(new_n761), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n221), .A2(G190), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n769), .A2(new_n265), .A3(new_n282), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT95), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n221), .A2(new_n481), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n265), .A2(new_n282), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT94), .ZN(new_n778));
  AND3_X1   g0578(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n778), .B1(new_n776), .B2(new_n777), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n775), .A2(G329), .B1(G326), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n265), .A2(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n776), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n282), .A2(G179), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n769), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G322), .A2(new_n786), .B1(new_n789), .B2(G283), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n777), .A2(new_n769), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(KEYINPUT33), .B(G317), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n776), .A2(new_n787), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n792), .A2(new_n793), .B1(new_n795), .B2(G303), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n784), .A2(new_n769), .ZN(new_n797));
  INV_X1    g0597(.A(G311), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n342), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n481), .A2(G179), .A3(G200), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n221), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n799), .B1(G294), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n783), .A2(new_n790), .A3(new_n796), .A4(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(G159), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n774), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT97), .ZN(new_n807));
  XNOR2_X1  g0607(.A(KEYINPUT96), .B(KEYINPUT32), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n807), .B(new_n808), .Z(new_n809));
  NOR2_X1   g0609(.A1(new_n781), .A2(new_n317), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n801), .A2(new_n445), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n258), .B1(new_n791), .B2(new_n212), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n794), .A2(new_n534), .B1(new_n788), .B2(new_n262), .ZN(new_n813));
  NOR4_X1   g0613(.A1(new_n810), .A2(new_n811), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n785), .A2(new_n210), .B1(new_n797), .B2(new_n202), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT93), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n804), .B1(new_n809), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n768), .B1(new_n818), .B2(new_n765), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n764), .B(KEYINPUT98), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n819), .B1(new_n675), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n753), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(G396));
  OR2_X1    g0624(.A1(new_n266), .A2(new_n280), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(new_n669), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n283), .A2(new_n284), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n669), .A2(new_n279), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n826), .B1(new_n829), .B2(new_n825), .ZN(new_n830));
  OR2_X1    g0630(.A1(new_n742), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n670), .B(new_n830), .C1(new_n633), .C2(new_n639), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n834), .A2(new_n729), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n751), .B1(new_n834), .B2(new_n729), .ZN(new_n837));
  INV_X1    g0637(.A(new_n826), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n829), .A2(new_n825), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n762), .ZN(new_n841));
  INV_X1    g0641(.A(new_n765), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n788), .A2(new_n212), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n342), .B(new_n843), .C1(G50), .C2(new_n795), .ZN(new_n844));
  INV_X1    g0644(.A(G132), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n844), .B1(new_n210), .B2(new_n801), .C1(new_n845), .C2(new_n774), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n846), .A2(KEYINPUT99), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(KEYINPUT99), .ZN(new_n848));
  INV_X1    g0648(.A(new_n797), .ZN(new_n849));
  AOI22_X1  g0649(.A1(G143), .A2(new_n786), .B1(new_n849), .B2(G159), .ZN(new_n850));
  INV_X1    g0650(.A(G137), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n850), .B1(new_n332), .B2(new_n791), .C1(new_n781), .C2(new_n851), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT34), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n847), .A2(new_n848), .A3(new_n853), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n775), .A2(G311), .B1(G303), .B2(new_n782), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n788), .A2(new_n534), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n794), .A2(new_n262), .B1(new_n797), .B2(new_n442), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n856), .B(new_n857), .C1(G294), .C2(new_n786), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n258), .B(new_n811), .C1(G283), .C2(new_n792), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n855), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n842), .B1(new_n854), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n765), .A2(new_n762), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n752), .B(new_n861), .C1(new_n202), .C2(new_n862), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT100), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n836), .A2(new_n837), .B1(new_n841), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(G384));
  OAI211_X1 g0666(.A(G116), .B(new_n222), .C1(new_n504), .C2(KEYINPUT35), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(KEYINPUT35), .B2(new_n504), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT36), .ZN(new_n869));
  OR3_X1    g0669(.A1(new_n227), .A2(new_n202), .A3(new_n366), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n317), .A2(G68), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n247), .B(G13), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n713), .A2(KEYINPUT31), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n724), .A2(new_n725), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n724), .A2(KEYINPUT31), .A3(new_n725), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT40), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT102), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n372), .A2(new_n274), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n399), .B1(new_n881), .B2(new_n373), .ZN(new_n882));
  INV_X1    g0682(.A(new_n667), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n411), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n404), .A2(new_n882), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n403), .A2(G190), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n282), .B2(new_n403), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n884), .B(new_n887), .C1(new_n400), .C2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n400), .A2(new_n404), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n883), .B1(new_n647), .B2(new_n360), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT37), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n376), .A2(new_n407), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n892), .A2(new_n893), .A3(new_n894), .A4(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  AND4_X1   g0697(.A1(new_n880), .A2(new_n886), .A3(KEYINPUT38), .A4(new_n897), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n411), .A2(new_n885), .B1(new_n891), .B2(new_n896), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n880), .B1(new_n899), .B2(KEYINPUT38), .ZN(new_n900));
  INV_X1    g0700(.A(new_n649), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n642), .B1(new_n400), .B2(new_n404), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n376), .A2(new_n396), .A3(KEYINPUT84), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n641), .A2(new_n648), .A3(new_n649), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n904), .A2(new_n656), .A3(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n893), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n641), .A2(new_n648), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n893), .A2(new_n895), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT37), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n906), .A2(new_n907), .B1(new_n896), .B2(new_n910), .ZN(new_n911));
  OAI22_X1  g0711(.A1(new_n898), .A2(new_n900), .B1(KEYINPUT38), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n324), .A2(new_n669), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n329), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n325), .A2(KEYINPUT101), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT101), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n310), .A2(new_n916), .A3(new_n324), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n914), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n325), .A2(new_n670), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n830), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(new_n876), .B2(new_n877), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n879), .B1(new_n912), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n886), .A2(new_n897), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT38), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n886), .A2(KEYINPUT38), .A3(new_n897), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT40), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n920), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n927), .A2(new_n878), .A3(new_n928), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n412), .B(new_n878), .C1(new_n922), .C2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(G330), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n926), .A2(KEYINPUT102), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n899), .A2(new_n880), .A3(KEYINPUT38), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n906), .A2(new_n907), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n910), .A2(new_n896), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n932), .A2(new_n933), .B1(new_n936), .B2(new_n924), .ZN(new_n937));
  INV_X1    g0737(.A(new_n877), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n928), .B1(new_n726), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(KEYINPUT40), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n921), .A2(new_n927), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n931), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n878), .A2(new_n412), .A3(G330), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n930), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n737), .B(new_n412), .C1(new_n742), .C2(KEYINPUT29), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n660), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n945), .B(new_n947), .Z(new_n948));
  NAND2_X1  g0748(.A1(new_n925), .A2(new_n926), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n832), .A2(new_n838), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n918), .A2(new_n919), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n949), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n667), .B1(new_n650), .B2(new_n651), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n932), .A2(new_n933), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT39), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n893), .B1(new_n652), .B2(new_n656), .ZN(new_n958));
  INV_X1    g0758(.A(new_n935), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n924), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n956), .A2(new_n957), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n957), .B1(new_n925), .B2(new_n926), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n915), .A2(new_n670), .A3(new_n917), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n955), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n948), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n247), .B2(new_n663), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n948), .A2(new_n967), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n873), .B1(new_n969), .B2(new_n970), .ZN(G367));
  NOR2_X1   g0771(.A1(new_n237), .A2(new_n759), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n766), .B1(new_n206), .B2(new_n271), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n751), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  AOI22_X1  g0774(.A1(G294), .A2(new_n792), .B1(new_n786), .B2(G303), .ZN(new_n975));
  INV_X1    g0775(.A(G283), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n975), .B1(new_n976), .B2(new_n797), .C1(new_n798), .C2(new_n781), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n342), .B1(new_n788), .B2(new_n445), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n794), .A2(new_n442), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n978), .B1(KEYINPUT46), .B2(new_n979), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n980), .B1(KEYINPUT46), .B2(new_n979), .C1(new_n262), .C2(new_n801), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n977), .B(new_n981), .C1(G317), .C2(new_n775), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT104), .ZN(new_n983));
  AOI22_X1  g0783(.A1(G159), .A2(new_n792), .B1(new_n849), .B2(G50), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n984), .A2(KEYINPUT105), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(G137), .B2(new_n775), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n258), .B1(new_n794), .B2(new_n210), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n785), .A2(new_n332), .B1(new_n788), .B2(new_n202), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n987), .B(new_n988), .C1(G68), .C2(new_n802), .ZN(new_n989));
  AOI22_X1  g0789(.A1(G143), .A2(new_n782), .B1(new_n984), .B2(KEYINPUT105), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n986), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(KEYINPUT47), .B1(new_n983), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n992), .A2(new_n842), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n983), .A2(KEYINPUT47), .A3(new_n991), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n974), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n630), .B1(new_n551), .B2(new_n670), .ZN(new_n996));
  OR3_X1    g0796(.A1(new_n629), .A2(new_n670), .A3(new_n551), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n995), .B1(new_n821), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n748), .A2(new_n686), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n620), .B1(new_n616), .B2(new_n670), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n635), .A2(new_n669), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n698), .B2(new_n704), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT44), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n698), .A2(new_n704), .A3(new_n1003), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT45), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1000), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1004), .B(KEYINPUT44), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT45), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1007), .B(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1010), .A2(new_n685), .A3(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n686), .A2(new_n694), .A3(new_n695), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n748), .A2(new_n701), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n701), .A2(new_n1014), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n677), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n744), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1009), .A2(new_n1013), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n745), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n707), .B(KEYINPUT41), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n750), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n703), .A2(KEYINPUT42), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1003), .B(new_n1023), .C1(new_n696), .C2(new_n697), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1003), .ZN(new_n1025));
  OAI21_X1  g0825(.A(KEYINPUT42), .B1(new_n701), .B2(new_n1025), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1024), .B(new_n1026), .C1(new_n556), .C2(new_n669), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n998), .A2(KEYINPUT43), .ZN(new_n1028));
  OR3_X1    g0828(.A1(new_n1027), .A2(KEYINPUT103), .A3(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(KEYINPUT103), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n998), .A2(KEYINPUT43), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1027), .A2(new_n1028), .A3(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1033), .B(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n999), .B1(new_n1022), .B2(new_n1035), .ZN(G387));
  NAND2_X1  g0836(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n745), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1015), .A2(new_n1017), .A3(new_n744), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(new_n1039), .A3(new_n707), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n686), .A2(new_n820), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G311), .A2(new_n792), .B1(new_n849), .B2(G303), .ZN(new_n1042));
  INV_X1    g0842(.A(G317), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1042), .B1(new_n1043), .B2(new_n785), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G322), .B2(new_n782), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT48), .Z(new_n1046));
  INV_X1    g0846(.A(G294), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1046), .B1(new_n976), .B2(new_n801), .C1(new_n1047), .C2(new_n794), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT49), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n775), .A2(G326), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n258), .B1(new_n789), .B2(G116), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n795), .A2(G77), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n797), .B2(new_n212), .C1(new_n330), .C2(new_n791), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n342), .B(new_n1054), .C1(G97), .C2(new_n789), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n775), .A2(G150), .B1(G159), .B2(new_n782), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n801), .A2(new_n271), .B1(new_n785), .B2(new_n317), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT110), .Z(new_n1058));
  NAND3_X1  g0858(.A1(new_n1055), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n842), .B1(new_n1052), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n267), .A2(new_n317), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT108), .Z(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(KEYINPUT50), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n709), .B(new_n425), .C1(new_n212), .C2(new_n202), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT107), .Z(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1062), .A2(KEYINPUT50), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n758), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT109), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n234), .A2(G45), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT106), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1070), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n709), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n754), .A2(new_n1075), .B1(new_n262), .B2(new_n706), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n767), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n1060), .A2(new_n752), .A3(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1037), .A2(new_n750), .B1(new_n1041), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1040), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT111), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1040), .A2(KEYINPUT111), .A3(new_n1079), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(G393));
  INV_X1    g0884(.A(KEYINPUT113), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1019), .A2(new_n707), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1018), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1006), .A2(new_n1008), .A3(new_n1000), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n685), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1038), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1091), .A2(KEYINPUT113), .A3(new_n707), .A4(new_n1019), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1009), .A2(new_n750), .A3(new_n1013), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n245), .A2(new_n759), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n766), .B1(new_n445), .B2(new_n206), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n751), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n342), .B1(new_n788), .B2(new_n262), .C1(new_n801), .C2(new_n442), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n792), .A2(G303), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1098), .B1(new_n976), .B2(new_n794), .C1(new_n1047), .C2(new_n797), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1097), .B(new_n1099), .C1(G322), .C2(new_n775), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n781), .A2(new_n1043), .B1(new_n798), .B2(new_n785), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT52), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n781), .A2(new_n332), .B1(new_n805), .B2(new_n785), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT51), .Z(new_n1105));
  INV_X1    g0905(.A(G143), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n774), .A2(new_n1106), .B1(new_n212), .B2(new_n794), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n1107), .A2(KEYINPUT112), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(KEYINPUT112), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n330), .A2(new_n797), .B1(new_n317), .B2(new_n791), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n801), .A2(new_n202), .ZN(new_n1111));
  NOR4_X1   g0911(.A1(new_n1110), .A2(new_n1111), .A3(new_n342), .A4(new_n856), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1108), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1103), .B1(new_n1105), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1096), .B1(new_n1114), .B2(new_n765), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n764), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1115), .B1(new_n1003), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1093), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1088), .A2(new_n1092), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(KEYINPUT114), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1091), .A2(new_n707), .A3(new_n1019), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1118), .B1(new_n1122), .B2(new_n1085), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT114), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1123), .A2(new_n1124), .A3(new_n1092), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1121), .A2(new_n1125), .ZN(G390));
  OAI211_X1 g0926(.A(new_n670), .B(new_n839), .C1(new_n730), .C2(new_n736), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n838), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT115), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1127), .A2(KEYINPUT115), .A3(new_n838), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1130), .A2(new_n952), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n966), .B1(new_n956), .B2(new_n960), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n826), .B1(new_n742), .B2(new_n830), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n965), .B1(new_n1135), .B2(new_n951), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1136), .A2(new_n963), .A3(new_n961), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n728), .A2(G330), .A3(new_n928), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n1134), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n878), .A2(G330), .A3(new_n928), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n962), .B1(new_n937), .B2(new_n957), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n762), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n775), .A2(G294), .B1(G283), .B2(new_n782), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n785), .A2(new_n442), .B1(new_n797), .B2(new_n445), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n843), .B(new_n1146), .C1(G107), .C2(new_n792), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n258), .B(new_n1111), .C1(G87), .C2(new_n795), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1145), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n845), .A2(new_n785), .B1(new_n791), .B2(new_n851), .ZN(new_n1150));
  XOR2_X1   g0950(.A(KEYINPUT54), .B(G143), .Z(new_n1151));
  AOI21_X1  g0951(.A(new_n1150), .B1(new_n849), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(G125), .ZN(new_n1153));
  INV_X1    g0953(.A(G128), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n1152), .B1(new_n1153), .B2(new_n774), .C1(new_n1154), .C2(new_n781), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n794), .A2(new_n332), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT53), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n342), .B1(new_n789), .B2(G50), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1157), .B(new_n1158), .C1(new_n805), .C2(new_n801), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1149), .B1(new_n1155), .B2(new_n1159), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n1160), .A2(new_n765), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n752), .B(new_n1161), .C1(new_n330), .C2(new_n862), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n1142), .A2(new_n750), .B1(new_n1144), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT116), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1134), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n1143), .A2(new_n1136), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1165), .B1(new_n1166), .B2(new_n1140), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n943), .A2(new_n660), .A3(new_n946), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1170));
  OAI211_X1 g0970(.A(G330), .B(new_n830), .C1(new_n726), .C2(new_n938), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n951), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1138), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(G330), .B(new_n830), .C1(new_n726), .C2(new_n727), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n951), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1135), .B1(new_n1175), .B2(new_n1140), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1169), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1164), .B1(new_n1167), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1141), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1175), .A2(new_n1140), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n950), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1138), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1168), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1179), .A2(new_n1183), .A3(KEYINPUT116), .A4(new_n1165), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1178), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT117), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n708), .B1(new_n1167), .B2(new_n1177), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1186), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1163), .B1(new_n1188), .B2(new_n1189), .ZN(G378));
  AOI21_X1  g0990(.A(KEYINPUT116), .B1(new_n1142), .B2(new_n1183), .ZN(new_n1191));
  NOR3_X1   g0991(.A1(new_n1167), .A2(new_n1177), .A3(new_n1164), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1169), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n357), .B(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n883), .A2(new_n337), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT118), .Z(new_n1197));
  XOR2_X1   g0997(.A(new_n1195), .B(new_n1197), .Z(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n954), .B(new_n953), .C1(new_n1143), .C2(new_n965), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1200), .A2(new_n942), .ZN(new_n1201));
  OAI21_X1  g1001(.A(G330), .B1(new_n922), .B2(new_n929), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n967), .A2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1199), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1200), .A2(new_n942), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n967), .A2(new_n1202), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(new_n1198), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1204), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1193), .A2(KEYINPUT57), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT57), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1168), .B1(new_n1178), .B2(new_n1184), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1211), .B1(new_n1212), .B2(new_n1208), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1210), .A2(new_n1213), .A3(new_n707), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n251), .A2(new_n252), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n317), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n252), .B2(new_n342), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n774), .A2(new_n976), .B1(new_n442), .B2(new_n781), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1053), .B1(new_n785), .B2(new_n262), .C1(new_n801), .C2(new_n212), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n791), .A2(new_n445), .B1(new_n797), .B2(new_n271), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n252), .B(new_n342), .C1(new_n788), .C2(new_n210), .ZN(new_n1221));
  NOR4_X1   g1021(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1217), .B1(new_n1222), .B2(KEYINPUT58), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n1154), .A2(new_n785), .B1(new_n791), .B2(new_n845), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1151), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n1225), .A2(new_n794), .B1(new_n797), .B2(new_n851), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1224), .B(new_n1226), .C1(G150), .C2(new_n802), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n1153), .B2(new_n781), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n775), .A2(G124), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1215), .B1(new_n789), .B2(G159), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1223), .B1(KEYINPUT58), .B2(new_n1222), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n765), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n752), .B1(new_n317), .B2(new_n862), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1235), .B(new_n1236), .C1(new_n1198), .C2(new_n763), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n1208), .B2(new_n749), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1214), .A2(new_n1239), .ZN(G375));
  NAND2_X1  g1040(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1241));
  OR3_X1    g1041(.A1(new_n1241), .A2(KEYINPUT119), .A3(new_n1169), .ZN(new_n1242));
  OAI21_X1  g1042(.A(KEYINPUT119), .B1(new_n1241), .B2(new_n1169), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1244), .A2(new_n1021), .A3(new_n1177), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1241), .A2(new_n750), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n752), .B1(new_n212), .B2(new_n862), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n258), .B1(new_n788), .B2(new_n210), .C1(new_n801), .C2(new_n317), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n1225), .A2(new_n791), .B1(new_n805), .B2(new_n794), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n785), .A2(new_n851), .B1(new_n797), .B2(new_n332), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n775), .A2(G128), .B1(G132), .B2(new_n782), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n775), .A2(G303), .B1(G294), .B2(new_n782), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n342), .B1(new_n788), .B2(new_n202), .C1(new_n801), .C2(new_n271), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n785), .A2(new_n976), .B1(new_n797), .B2(new_n262), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n445), .A2(new_n794), .B1(new_n791), .B2(new_n442), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1251), .A2(new_n1252), .B1(new_n1253), .B2(new_n1257), .ZN(new_n1258));
  OAI221_X1 g1058(.A(new_n1247), .B1(new_n842), .B2(new_n1258), .C1(new_n952), .C2(new_n763), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1246), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1245), .A2(new_n1261), .ZN(G381));
  NOR2_X1   g1062(.A1(G393), .A2(G396), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n865), .ZN(new_n1264));
  NOR3_X1   g1064(.A1(new_n1264), .A2(G387), .A3(G381), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1121), .A2(new_n1125), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1208), .B1(new_n1185), .B2(new_n1169), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n708), .B1(new_n1267), .B2(KEYINPUT57), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1238), .B1(new_n1268), .B2(new_n1213), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1163), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1265), .A2(new_n1266), .A3(new_n1269), .A4(new_n1272), .ZN(G407));
  NAND3_X1  g1073(.A1(new_n1269), .A2(new_n668), .A3(new_n1272), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(G407), .A2(G213), .A3(new_n1274), .ZN(G409));
  XOR2_X1   g1075(.A(KEYINPUT123), .B(KEYINPUT61), .Z(new_n1276));
  NOR2_X1   g1076(.A1(new_n662), .A2(G343), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1021), .ZN(new_n1278));
  NOR3_X1   g1078(.A1(new_n1212), .A2(new_n1278), .A3(new_n1208), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT120), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1239), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NOR4_X1   g1081(.A1(new_n1212), .A2(new_n1208), .A3(KEYINPUT120), .A4(new_n1278), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1272), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1214), .A2(G378), .A3(new_n1239), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1277), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1177), .A2(KEYINPUT60), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1244), .A2(new_n1286), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1181), .A2(KEYINPUT60), .A3(new_n1182), .A4(new_n1168), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n707), .ZN(new_n1289));
  OAI211_X1 g1089(.A(G384), .B(new_n1261), .C1(new_n1287), .C2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1289), .B1(new_n1244), .B2(new_n1286), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n865), .B1(new_n1292), .B2(new_n1260), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  OAI211_X1 g1094(.A(G2897), .B(new_n1277), .C1(new_n1291), .C2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1277), .A2(G2897), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1290), .A2(new_n1293), .A3(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1276), .B1(new_n1285), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT124), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  OAI211_X1 g1101(.A(KEYINPUT124), .B(new_n1276), .C1(new_n1285), .C2(new_n1298), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1291), .A2(new_n1294), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1285), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(KEYINPUT62), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT62), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1285), .A2(new_n1306), .A3(new_n1303), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1301), .A2(new_n1302), .A3(new_n1305), .A4(new_n1307), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1266), .A2(G387), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1121), .A2(new_n1125), .A3(G387), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n823), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1311));
  OR2_X1    g1111(.A1(new_n1263), .A2(new_n1311), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1310), .A2(new_n1312), .A3(KEYINPUT122), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT121), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1312), .B1(new_n1310), .B2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1309), .B1(new_n1313), .B2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1310), .A2(new_n1314), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1312), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  OAI211_X1 g1119(.A(G390), .B(new_n999), .C1(new_n1022), .C2(new_n1035), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1310), .A2(new_n1312), .A3(KEYINPUT122), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1319), .A2(new_n1320), .A3(new_n1321), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1316), .A2(new_n1322), .A3(KEYINPUT125), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT125), .B1(new_n1316), .B2(new_n1322), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1308), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  NOR3_X1   g1125(.A1(new_n1313), .A2(new_n1315), .A3(new_n1309), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1320), .B1(new_n1319), .B2(new_n1321), .ZN(new_n1327));
  NOR3_X1   g1127(.A1(new_n1326), .A2(new_n1327), .A3(KEYINPUT61), .ZN(new_n1328));
  OAI21_X1  g1128(.A(KEYINPUT63), .B1(new_n1285), .B2(new_n1298), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(new_n1304), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1285), .A2(KEYINPUT63), .A3(new_n1303), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1328), .A2(new_n1330), .A3(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1325), .A2(new_n1332), .ZN(G405));
  INV_X1    g1133(.A(KEYINPUT126), .ZN(new_n1334));
  OAI211_X1 g1134(.A(new_n1284), .B(new_n1334), .C1(new_n1269), .C2(new_n1271), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT127), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1335), .A2(new_n1336), .A3(new_n1303), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1336), .B1(new_n1335), .B2(new_n1303), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(G375), .A2(new_n1272), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1334), .B1(new_n1340), .B2(new_n1284), .ZN(new_n1341));
  NOR3_X1   g1141(.A1(new_n1338), .A2(new_n1339), .A3(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1341), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1335), .A2(new_n1303), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1344), .A2(KEYINPUT127), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1343), .B1(new_n1345), .B2(new_n1337), .ZN(new_n1346));
  OAI22_X1  g1146(.A1(new_n1323), .A2(new_n1324), .B1(new_n1342), .B2(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT125), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1348), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1316), .A2(new_n1322), .A3(KEYINPUT125), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1345), .A2(new_n1337), .A3(new_n1343), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1341), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1349), .A2(new_n1350), .A3(new_n1351), .A4(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1347), .A2(new_n1353), .ZN(G402));
endmodule


