//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 0 0 1 0 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G250), .ZN(new_n205));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  OR3_X1    g0006(.A1(new_n206), .A2(KEYINPUT64), .A3(G13), .ZN(new_n207));
  OAI21_X1  g0007(.A(KEYINPUT64), .B1(new_n206), .B2(G13), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  INV_X1    g0011(.A(G264), .ZN(new_n212));
  AOI211_X1 g0012(.A(new_n205), .B(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n213), .A2(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(KEYINPUT0), .ZN(new_n215));
  AND2_X1   g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G20), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT65), .Z(new_n218));
  OAI21_X1  g0018(.A(G50), .B1(G58), .B2(G68), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT66), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n214), .B(new_n215), .C1(new_n218), .C2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT67), .Z(new_n223));
  NAND2_X1  g0023(.A1(G116), .A2(G270), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G87), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n224), .B1(new_n202), .B2(new_n225), .C1(new_n226), .C2(new_n205), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n228));
  INV_X1    g0028(.A(G50), .ZN(new_n229));
  INV_X1    g0029(.A(G226), .ZN(new_n230));
  INV_X1    g0030(.A(G68), .ZN(new_n231));
  INV_X1    g0031(.A(G238), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n228), .B1(new_n229), .B2(new_n230), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n227), .B(new_n233), .C1(G97), .C2(G257), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(G1), .B2(G20), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(KEYINPUT1), .Z(new_n236));
  NOR2_X1   g0036(.A1(new_n223), .A2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  INV_X1    g0038(.A(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G250), .B(G257), .Z(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G358));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G222), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G223), .A2(G1698), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n255), .A2(new_n257), .A3(new_n259), .A4(new_n260), .ZN(new_n261));
  AND2_X1   g0061(.A1(G33), .A2(G41), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G1), .A2(G13), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT3), .B(G33), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n261), .B(new_n264), .C1(G77), .C2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n262), .A2(KEYINPUT68), .A3(new_n263), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT68), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n270), .B1(new_n216), .B2(new_n271), .ZN(new_n272));
  OAI211_X1 g0072(.A(G226), .B(new_n268), .C1(new_n269), .C2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  INV_X1    g0074(.A(G45), .ZN(new_n275));
  AOI21_X1  g0075(.A(G1), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI211_X1 g0076(.A(G274), .B(new_n276), .C1(new_n269), .C2(new_n272), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n266), .A2(new_n273), .A3(new_n277), .A4(G190), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT74), .ZN(new_n279));
  XNOR2_X1  g0079(.A(new_n278), .B(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G13), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(G1), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G20), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n229), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n229), .B1(new_n267), .B2(G20), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n263), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT69), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(KEYINPUT69), .B1(new_n287), .B2(new_n263), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n283), .B(new_n286), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G20), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n256), .ZN(new_n294));
  INV_X1    g0094(.A(G150), .ZN(new_n295));
  OAI22_X1  g0095(.A1(new_n201), .A2(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT72), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(new_n256), .B2(G20), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n293), .A2(KEYINPUT72), .A3(G33), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(KEYINPUT71), .A2(KEYINPUT8), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G58), .ZN(new_n303));
  INV_X1    g0103(.A(G58), .ZN(new_n304));
  NOR3_X1   g0104(.A1(new_n304), .A2(KEYINPUT70), .A3(KEYINPUT71), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT70), .ZN(new_n306));
  OAI21_X1  g0106(.A(KEYINPUT8), .B1(new_n306), .B2(G58), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n303), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n296), .B1(new_n301), .B2(new_n308), .ZN(new_n309));
  OR2_X1    g0109(.A1(new_n290), .A2(new_n291), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n285), .B(new_n292), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT9), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n290), .A2(new_n291), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n304), .A2(KEYINPUT70), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n306), .A2(G58), .ZN(new_n315));
  OAI211_X1 g0115(.A(KEYINPUT8), .B(new_n314), .C1(new_n315), .C2(KEYINPUT71), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n300), .B1(new_n316), .B2(new_n303), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n313), .B1(new_n317), .B2(new_n296), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT9), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n318), .A2(new_n319), .A3(new_n285), .A4(new_n292), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n312), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT10), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n266), .A2(new_n273), .A3(new_n277), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G200), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n280), .A2(new_n321), .A3(new_n322), .A4(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT76), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT75), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n280), .A2(new_n321), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n328), .B1(new_n280), .B2(new_n321), .ZN(new_n330));
  INV_X1    g0130(.A(new_n324), .ZN(new_n331));
  NOR3_X1   g0131(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n327), .B1(new_n332), .B2(new_n322), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n280), .A2(new_n321), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT75), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n280), .A2(new_n321), .A3(new_n328), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(new_n336), .A3(new_n324), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n337), .A2(KEYINPUT76), .A3(KEYINPUT10), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n326), .B1(new_n333), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT15), .B(G87), .ZN(new_n340));
  OR2_X1    g0140(.A1(new_n300), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT73), .ZN(new_n342));
  INV_X1    g0142(.A(new_n294), .ZN(new_n343));
  XOR2_X1   g0143(.A(KEYINPUT8), .B(G58), .Z(new_n344));
  AOI22_X1  g0144(.A1(new_n341), .A2(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI221_X1 g0145(.A(new_n345), .B1(new_n342), .B2(new_n341), .C1(new_n293), .C2(new_n202), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n346), .A2(new_n288), .B1(new_n202), .B2(new_n284), .ZN(new_n347));
  INV_X1    g0147(.A(new_n288), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n267), .A2(G20), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(G77), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G274), .ZN(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT68), .B1(new_n262), .B2(new_n263), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n216), .A2(new_n270), .A3(new_n271), .ZN(new_n354));
  AOI211_X1 g0154(.A(new_n352), .B(new_n268), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n276), .B1(new_n353), .B2(new_n354), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n355), .B1(G244), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n255), .A2(new_n257), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n358), .B1(G232), .B2(new_n258), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n232), .B2(new_n258), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(G107), .B2(new_n265), .ZN(new_n361));
  INV_X1    g0161(.A(new_n264), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n357), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G169), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n363), .A2(G179), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n351), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G190), .ZN(new_n369));
  OR2_X1    g0169(.A1(new_n363), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n363), .A2(G200), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n370), .A2(new_n347), .A3(new_n350), .A4(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  OR2_X1    g0173(.A1(new_n323), .A2(G179), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n323), .A2(new_n364), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n374), .A2(new_n311), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NOR3_X1   g0177(.A1(new_n368), .A2(new_n373), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT77), .B1(new_n339), .B2(new_n379), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n332), .A2(new_n327), .A3(new_n322), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT76), .B1(new_n337), .B2(KEYINPUT10), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n325), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT77), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(new_n384), .A3(new_n378), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n230), .A2(new_n258), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n239), .A2(G1698), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n265), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G97), .ZN(new_n390));
  AOI211_X1 g0190(.A(KEYINPUT78), .B(new_n362), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT78), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n389), .A2(new_n390), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n392), .B1(new_n393), .B2(new_n264), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n356), .A2(G238), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n277), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n395), .A2(KEYINPUT13), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT13), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n393), .A2(new_n264), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT78), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n393), .A2(new_n392), .A3(new_n264), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n397), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n399), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(G169), .B1(new_n398), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT14), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT13), .B1(new_n395), .B2(new_n397), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n403), .A2(new_n399), .A3(new_n404), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT14), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(new_n411), .A3(G169), .ZN(new_n412));
  INV_X1    g0212(.A(G179), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n407), .B(new_n412), .C1(new_n413), .C2(new_n410), .ZN(new_n414));
  OAI22_X1  g0214(.A1(new_n300), .A2(new_n202), .B1(new_n229), .B2(new_n294), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n293), .A2(G68), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n313), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT11), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n348), .A2(G68), .A3(new_n349), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n417), .B2(new_n418), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n282), .A2(new_n416), .ZN(new_n422));
  XOR2_X1   g0222(.A(new_n422), .B(KEYINPUT12), .Z(new_n423));
  NOR3_X1   g0223(.A1(new_n419), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n414), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n410), .A2(G200), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n408), .A2(new_n409), .A3(G190), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT87), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT18), .ZN(new_n432));
  NAND2_X1  g0232(.A1(G33), .A2(G87), .ZN(new_n433));
  XOR2_X1   g0233(.A(new_n433), .B(KEYINPUT84), .Z(new_n434));
  AND2_X1   g0234(.A1(KEYINPUT79), .A2(G33), .ZN(new_n435));
  NOR2_X1   g0235(.A1(KEYINPUT79), .A2(G33), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT3), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT80), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n438), .A2(new_n254), .A3(G33), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n255), .A2(KEYINPUT80), .ZN(new_n440));
  OR2_X1    g0240(.A1(G223), .A2(G1698), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n437), .A2(new_n439), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n258), .A2(G226), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n434), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n264), .ZN(new_n445));
  AOI211_X1 g0245(.A(new_n239), .B(new_n276), .C1(new_n353), .C2(new_n354), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n445), .A2(new_n413), .A3(new_n277), .A4(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT85), .ZN(new_n449));
  AOI211_X1 g0249(.A(new_n355), .B(new_n446), .C1(new_n444), .C2(new_n264), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n448), .B(new_n449), .C1(new_n450), .C2(G169), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n445), .A2(new_n277), .A3(new_n447), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n364), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n449), .B1(new_n454), .B2(new_n448), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n313), .A2(new_n284), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n308), .A2(new_n349), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(new_n283), .B2(new_n308), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT83), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT82), .ZN(new_n463));
  AOI21_X1  g0263(.A(G20), .B1(new_n255), .B2(new_n257), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n463), .B1(new_n464), .B2(KEYINPUT7), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT7), .ZN(new_n466));
  OAI211_X1 g0266(.A(KEYINPUT82), .B(new_n466), .C1(new_n265), .C2(G20), .ZN(new_n467));
  OR2_X1    g0267(.A1(KEYINPUT79), .A2(G33), .ZN(new_n468));
  NAND2_X1  g0268(.A1(KEYINPUT79), .A2(G33), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n468), .A2(new_n254), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(G20), .B1(new_n470), .B2(new_n257), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n465), .A2(new_n467), .B1(new_n471), .B2(KEYINPUT7), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n462), .B1(new_n472), .B2(new_n231), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n470), .A2(new_n257), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(KEYINPUT7), .A3(new_n293), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n358), .A2(new_n293), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT82), .B1(new_n476), .B2(new_n466), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n464), .A2(new_n463), .A3(KEYINPUT7), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n479), .A2(KEYINPUT83), .A3(G68), .ZN(new_n480));
  NOR2_X1   g0280(.A1(G58), .A2(G68), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n314), .A2(new_n315), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n481), .B1(new_n482), .B2(G68), .ZN(new_n483));
  INV_X1    g0283(.A(G159), .ZN(new_n484));
  OAI22_X1  g0284(.A1(new_n483), .A2(new_n293), .B1(new_n484), .B2(new_n294), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n473), .A2(new_n480), .A3(new_n486), .ZN(new_n487));
  XOR2_X1   g0287(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n437), .A2(new_n439), .A3(new_n440), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n293), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n231), .B1(new_n492), .B2(KEYINPUT7), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n491), .A2(new_n466), .A3(new_n293), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n485), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n348), .B1(new_n495), .B2(KEYINPUT16), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n461), .B1(new_n490), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n432), .B1(new_n456), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n448), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n446), .B1(new_n444), .B2(new_n264), .ZN(new_n500));
  AOI21_X1  g0300(.A(G169), .B1(new_n500), .B2(new_n277), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT85), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n451), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n492), .A2(KEYINPUT7), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(G68), .A3(new_n494), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(KEYINPUT16), .A3(new_n486), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n288), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n507), .B1(new_n489), .B2(new_n487), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n503), .B(KEYINPUT18), .C1(new_n508), .C2(new_n461), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n498), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n490), .A2(new_n496), .ZN(new_n511));
  INV_X1    g0311(.A(new_n461), .ZN(new_n512));
  INV_X1    g0312(.A(G200), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n453), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(G190), .B2(new_n453), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n511), .A2(KEYINPUT86), .A3(new_n512), .A4(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT17), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n497), .A2(KEYINPUT86), .A3(KEYINPUT17), .A4(new_n515), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n431), .B1(new_n510), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n498), .A2(new_n509), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n522), .A2(KEYINPUT87), .A3(new_n518), .A4(new_n519), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n430), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n386), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT88), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT88), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n386), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT24), .ZN(new_n530));
  NOR4_X1   g0330(.A1(new_n358), .A2(KEYINPUT22), .A3(G20), .A4(new_n226), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n438), .B1(new_n254), .B2(G33), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n468), .A2(new_n469), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n532), .B1(new_n533), .B2(KEYINPUT3), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n534), .A2(new_n293), .A3(G87), .A4(new_n439), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n531), .B1(new_n535), .B2(KEYINPUT22), .ZN(new_n536));
  INV_X1    g0336(.A(G107), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G20), .ZN(new_n538));
  XOR2_X1   g0338(.A(new_n538), .B(KEYINPUT23), .Z(new_n539));
  INV_X1    g0339(.A(G116), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n533), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT93), .B1(new_n541), .B2(new_n293), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n435), .A2(new_n436), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n543), .A2(new_n293), .A3(G116), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT93), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n539), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n530), .B1(new_n536), .B2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n437), .A2(new_n293), .A3(new_n439), .A4(new_n440), .ZN(new_n549));
  OAI21_X1  g0349(.A(KEYINPUT22), .B1(new_n549), .B2(new_n226), .ZN(new_n550));
  INV_X1    g0350(.A(new_n531), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g0352(.A(new_n544), .B(new_n545), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n552), .A2(KEYINPUT24), .A3(new_n539), .A4(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n548), .A2(new_n554), .A3(new_n288), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n282), .A2(G20), .A3(new_n537), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(KEYINPUT25), .ZN(new_n557));
  OR2_X1    g0357(.A1(new_n556), .A2(KEYINPUT25), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n267), .A2(G33), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n283), .B(new_n559), .C1(new_n290), .C2(new_n291), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n557), .B(new_n558), .C1(new_n560), .C2(new_n537), .ZN(new_n561));
  XNOR2_X1  g0361(.A(new_n561), .B(KEYINPUT94), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(G257), .A2(G1698), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n205), .B2(G1698), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n437), .A2(new_n439), .A3(new_n440), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n543), .A2(G294), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n264), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n353), .A2(new_n354), .ZN(new_n570));
  OR2_X1    g0370(.A1(new_n274), .A2(KEYINPUT5), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n274), .A2(KEYINPUT5), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n275), .A2(G1), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n570), .A2(G264), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n572), .A2(KEYINPUT90), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n267), .B(G45), .C1(new_n274), .C2(KEYINPUT5), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n572), .A2(KEYINPUT90), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n576), .A2(new_n276), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n569), .A2(new_n575), .A3(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n582), .A2(G190), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT95), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n569), .A2(new_n584), .A3(new_n575), .ZN(new_n585));
  INV_X1    g0385(.A(new_n575), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n362), .B1(new_n566), .B2(new_n567), .ZN(new_n587));
  OAI21_X1  g0387(.A(KEYINPUT95), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n585), .A2(new_n588), .A3(new_n581), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n583), .B1(new_n589), .B2(new_n513), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n563), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n585), .A2(new_n588), .A3(G179), .A4(new_n581), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n582), .A2(G169), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n555), .A2(new_n562), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n358), .A2(G303), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n211), .A2(new_n258), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n437), .A2(new_n439), .A3(new_n440), .A4(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n258), .A2(G264), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n595), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n264), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n570), .A2(G270), .A3(new_n574), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n600), .A2(G190), .A3(new_n581), .A4(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n282), .A2(G20), .A3(new_n540), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n348), .A2(new_n283), .A3(G116), .A4(new_n559), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n287), .A2(new_n263), .B1(G20), .B2(new_n540), .ZN(new_n605));
  AOI21_X1  g0405(.A(G20), .B1(G33), .B2(G283), .ZN(new_n606));
  INV_X1    g0406(.A(G97), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n606), .B1(G33), .B2(new_n607), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n605), .A2(new_n608), .A3(KEYINPUT20), .ZN(new_n609));
  AOI21_X1  g0409(.A(KEYINPUT20), .B1(new_n605), .B2(new_n608), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n603), .B(new_n604), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n598), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n534), .A2(new_n439), .A3(new_n613), .A4(new_n596), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n362), .B1(new_n614), .B2(new_n595), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n581), .A2(new_n601), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n602), .B(new_n612), .C1(new_n617), .C2(new_n513), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT21), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n611), .A2(G169), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n619), .B1(new_n617), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n600), .A2(new_n581), .A3(new_n601), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n622), .A2(KEYINPUT21), .A3(G169), .A4(new_n611), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n617), .A2(G179), .A3(new_n611), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n618), .A2(new_n621), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n591), .A2(new_n594), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n343), .A2(G77), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n537), .A2(KEYINPUT6), .A3(G97), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n607), .A2(new_n537), .ZN(new_n629));
  NOR2_X1   g0429(.A1(G97), .A2(G107), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n628), .B1(new_n631), .B2(KEYINPUT6), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(G20), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n627), .B(new_n633), .C1(new_n472), .C2(new_n537), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n288), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n284), .A2(new_n607), .ZN(new_n636));
  INV_X1    g0436(.A(new_n560), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(G97), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n635), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT4), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n225), .A2(G1698), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n640), .B1(new_n491), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n641), .A2(new_n255), .A3(new_n257), .A4(KEYINPUT4), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n645), .A2(KEYINPUT89), .B1(G33), .B2(G283), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n265), .A2(G250), .A3(G1698), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT89), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n265), .A2(new_n648), .A3(KEYINPUT4), .A4(new_n641), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n646), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n264), .B1(new_n644), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n570), .A2(G257), .A3(new_n574), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(new_n581), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n364), .ZN(new_n654));
  INV_X1    g0454(.A(new_n581), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n643), .A2(new_n647), .A3(new_n649), .A4(new_n646), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n655), .B1(new_n656), .B2(new_n264), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n657), .A2(new_n413), .A3(new_n652), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n639), .A2(new_n654), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n653), .A2(G200), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n657), .A2(G190), .A3(new_n652), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n634), .A2(new_n288), .B1(new_n607), .B2(new_n284), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n660), .A2(new_n661), .A3(new_n662), .A4(new_n638), .ZN(new_n663));
  INV_X1    g0463(.A(new_n541), .ZN(new_n664));
  NOR2_X1   g0464(.A1(G238), .A2(G1698), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n665), .B1(new_n225), .B2(G1698), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n666), .A2(new_n437), .A3(new_n439), .A4(new_n440), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n264), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n275), .A2(G1), .A3(G274), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n570), .B(new_n671), .C1(G250), .C2(new_n573), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n364), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n226), .A2(new_n607), .A3(new_n537), .ZN(new_n675));
  AND2_X1   g0475(.A1(KEYINPUT91), .A2(KEYINPUT19), .ZN(new_n676));
  NOR2_X1   g0476(.A1(KEYINPUT91), .A2(KEYINPUT19), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n676), .A2(new_n677), .A3(new_n390), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n675), .B1(new_n678), .B2(G20), .ZN(new_n679));
  OAI22_X1  g0479(.A1(new_n300), .A2(new_n607), .B1(new_n677), .B2(new_n676), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n679), .B(new_n680), .C1(new_n549), .C2(new_n231), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n288), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n340), .B(KEYINPUT92), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n637), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n284), .A2(new_n340), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n682), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n669), .A2(new_n413), .A3(new_n672), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n674), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n681), .A2(new_n288), .B1(new_n284), .B2(new_n340), .ZN(new_n689));
  INV_X1    g0489(.A(new_n672), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n362), .B1(new_n664), .B2(new_n667), .ZN(new_n691));
  OAI21_X1  g0491(.A(G200), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n669), .A2(G190), .A3(new_n672), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n637), .A2(G87), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n689), .A2(new_n692), .A3(new_n693), .A4(new_n694), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n688), .A2(new_n695), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n659), .A2(new_n663), .A3(new_n696), .ZN(new_n697));
  AND3_X1   g0497(.A1(new_n529), .A2(new_n626), .A3(new_n697), .ZN(G372));
  INV_X1    g0498(.A(new_n659), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(KEYINPUT26), .A3(new_n695), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n663), .A2(new_n695), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n621), .A2(new_n623), .A3(new_n624), .ZN(new_n702));
  OAI22_X1  g0502(.A1(new_n594), .A2(new_n702), .B1(new_n563), .B2(new_n590), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n701), .B1(new_n703), .B2(new_n659), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n700), .B1(new_n704), .B2(KEYINPUT26), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n688), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n529), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n429), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n426), .B1(new_n367), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n520), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(KEYINPUT96), .B1(new_n498), .B2(new_n509), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n498), .A2(KEYINPUT96), .A3(new_n509), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT97), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n383), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n339), .A2(KEYINPUT97), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n377), .B1(new_n714), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n707), .A2(new_n719), .ZN(G369));
  NOR2_X1   g0520(.A1(new_n281), .A2(G20), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n267), .ZN(new_n722));
  OR2_X1    g0522(.A1(new_n722), .A2(KEYINPUT27), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(KEYINPUT27), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(G213), .A3(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G343), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n612), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n625), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n702), .B2(new_n728), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G330), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT98), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n591), .A2(new_n594), .ZN(new_n735));
  INV_X1    g0535(.A(new_n727), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n563), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n594), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n738), .B1(new_n739), .B2(new_n727), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n734), .A2(new_n740), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n702), .A2(new_n727), .ZN(new_n742));
  AOI22_X1  g0542(.A1(new_n735), .A2(new_n742), .B1(new_n594), .B2(new_n727), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n741), .A2(new_n743), .ZN(G399));
  NOR2_X1   g0544(.A1(new_n210), .A2(G41), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n675), .A2(G116), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n745), .A2(new_n267), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n747), .B1(new_n220), .B2(new_n745), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT28), .Z(new_n749));
  NOR2_X1   g0549(.A1(KEYINPUT100), .A2(KEYINPUT29), .ZN(new_n750));
  AOI211_X1 g0550(.A(new_n736), .B(new_n750), .C1(new_n705), .C2(new_n688), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n736), .B1(new_n705), .B2(new_n688), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  XNOR2_X1  g0553(.A(KEYINPUT100), .B(KEYINPUT29), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n751), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n626), .A2(new_n697), .A3(new_n727), .ZN(new_n756));
  NOR3_X1   g0556(.A1(new_n622), .A2(new_n673), .A3(new_n413), .ZN(new_n757));
  AND3_X1   g0557(.A1(new_n651), .A2(new_n581), .A3(new_n652), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n585), .A2(new_n588), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT30), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(G179), .B1(new_n657), .B2(new_n652), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n763), .A2(new_n589), .A3(new_n622), .A4(new_n673), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n757), .A2(new_n758), .A3(KEYINPUT30), .A4(new_n759), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n762), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(new_n736), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n756), .A2(KEYINPUT31), .A3(new_n767), .ZN(new_n768));
  XOR2_X1   g0568(.A(KEYINPUT99), .B(KEYINPUT31), .Z(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n766), .A2(new_n736), .A3(new_n770), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n771), .A2(G330), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n755), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n749), .B1(new_n774), .B2(G1), .ZN(G364));
  NOR2_X1   g0575(.A1(new_n210), .A2(new_n358), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G355), .ZN(new_n777));
  INV_X1    g0577(.A(new_n491), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n210), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(new_n221), .B2(G45), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n249), .A2(new_n275), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n777), .B1(G116), .B2(new_n209), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G13), .A2(G33), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(G20), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n263), .B1(G20), .B2(new_n364), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n782), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n267), .B1(new_n721), .B2(G45), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n745), .A2(new_n790), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n791), .B(KEYINPUT101), .Z(new_n792));
  NOR2_X1   g0592(.A1(new_n293), .A2(new_n413), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G190), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(G200), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n793), .A2(new_n369), .A3(G200), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n482), .A2(new_n795), .B1(new_n797), .B2(G68), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n293), .A2(G179), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n799), .A2(new_n369), .A3(G200), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n798), .B1(new_n537), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n793), .A2(new_n369), .A3(new_n513), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n794), .A2(new_n513), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n265), .B1(new_n202), .B2(new_n802), .C1(new_n804), .C2(new_n229), .ZN(new_n805));
  NOR2_X1   g0605(.A1(G179), .A2(G200), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n806), .A2(G20), .A3(new_n369), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n807), .A2(KEYINPUT32), .A3(new_n484), .ZN(new_n808));
  NOR3_X1   g0608(.A1(new_n801), .A2(new_n805), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(KEYINPUT32), .B1(new_n807), .B2(new_n484), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n293), .B1(new_n806), .B2(G190), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n811), .A2(KEYINPUT103), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(KEYINPUT103), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G97), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n799), .A2(G190), .A3(G200), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT102), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(G87), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n809), .A2(new_n810), .A3(new_n816), .A4(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(G311), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n802), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n807), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(G329), .ZN(new_n828));
  INV_X1    g0628(.A(G326), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n358), .B(new_n828), .C1(new_n804), .C2(new_n829), .ZN(new_n830));
  XOR2_X1   g0630(.A(KEYINPUT104), .B(G317), .Z(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT33), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n830), .B1(new_n797), .B2(new_n832), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n822), .A2(G303), .B1(new_n815), .B2(G294), .ZN(new_n834));
  INV_X1    g0634(.A(new_n800), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n795), .A2(G322), .B1(new_n835), .B2(G283), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n824), .B1(new_n826), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n792), .B1(new_n838), .B2(new_n786), .ZN(new_n839));
  INV_X1    g0639(.A(new_n785), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n788), .B(new_n839), .C1(new_n731), .C2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n791), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n731), .B2(G330), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n841), .B1(new_n734), .B2(new_n843), .ZN(G396));
  NAND2_X1  g0644(.A1(new_n368), .A2(new_n727), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n727), .B1(new_n347), .B2(new_n350), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n367), .B1(new_n373), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n752), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(new_n773), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n842), .ZN(new_n852));
  INV_X1    g0652(.A(G283), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n802), .A2(new_n540), .B1(new_n796), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(G303), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n358), .B1(new_n807), .B2(new_n825), .C1(new_n804), .C2(new_n855), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n854), .B(new_n856), .C1(G87), .C2(new_n835), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n795), .A2(G294), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n822), .A2(G107), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n857), .A2(new_n816), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(G143), .A2(new_n795), .B1(new_n797), .B2(G150), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n803), .A2(G137), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n861), .B(new_n862), .C1(new_n484), .C2(new_n802), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n863), .B(KEYINPUT34), .Z(new_n864));
  AOI22_X1  g0664(.A1(new_n815), .A2(new_n482), .B1(G68), .B2(new_n835), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n491), .B1(G132), .B2(new_n827), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n865), .B(new_n866), .C1(new_n229), .C2(new_n821), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n860), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n792), .B1(new_n868), .B2(new_n786), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n786), .A2(new_n783), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n869), .B1(G77), .B2(new_n871), .C1(new_n849), .C2(new_n784), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n852), .A2(new_n872), .ZN(G384));
  INV_X1    g0673(.A(new_n218), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n540), .B1(new_n632), .B2(KEYINPUT35), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n874), .B(new_n875), .C1(KEYINPUT35), .C2(new_n632), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n876), .B(KEYINPUT36), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n482), .A2(G68), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n220), .A2(G77), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(G50), .B2(new_n231), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n880), .A2(G1), .A3(new_n281), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n425), .A2(new_n736), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n408), .A2(new_n409), .A3(G179), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n407), .A2(new_n883), .A3(new_n412), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n429), .B(new_n882), .C1(new_n884), .C2(new_n424), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n425), .B(new_n736), .C1(new_n414), .C2(new_n708), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n848), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT31), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n766), .A2(new_n888), .A3(new_n736), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n756), .A2(new_n769), .A3(new_n767), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT106), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT40), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n887), .A2(new_n889), .A3(new_n890), .A4(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n497), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n503), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n726), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT37), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n511), .A2(new_n512), .A3(new_n515), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n895), .A2(new_n896), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n488), .B1(new_n505), .B2(new_n486), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT105), .B1(new_n900), .B2(new_n310), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT105), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n902), .B(new_n313), .C1(new_n495), .C2(new_n488), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n901), .A2(new_n506), .A3(new_n903), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n904), .A2(new_n512), .B1(new_n502), .B2(new_n451), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n725), .B1(new_n904), .B2(new_n512), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n511), .A2(new_n512), .A3(new_n515), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n899), .B1(new_n908), .B2(new_n897), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n906), .B1(new_n510), .B2(new_n520), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT38), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n909), .A2(new_n910), .A3(KEYINPUT38), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n893), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n885), .A2(new_n886), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n916), .A2(new_n890), .A3(new_n849), .A4(new_n889), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n891), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n710), .B1(new_n713), .B2(new_n712), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n497), .A2(new_n725), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n898), .B1(new_n497), .B2(new_n725), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n898), .B(KEYINPUT96), .C1(new_n497), .C2(new_n725), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n923), .A2(new_n895), .B1(new_n924), .B2(KEYINPUT37), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n456), .A2(new_n497), .ZN(new_n926));
  NOR4_X1   g0726(.A1(new_n922), .A2(new_n926), .A3(KEYINPUT96), .A4(new_n897), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT38), .B1(new_n921), .B2(new_n928), .ZN(new_n929));
  AND3_X1   g0729(.A1(new_n909), .A2(new_n910), .A3(KEYINPUT38), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n893), .B(new_n918), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n915), .B1(new_n931), .B2(KEYINPUT40), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n890), .A2(new_n889), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n529), .A2(new_n933), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n932), .B(new_n934), .Z(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(G330), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n426), .A2(new_n736), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n913), .A2(new_n914), .A3(KEYINPUT39), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n921), .A2(new_n928), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n930), .B1(new_n939), .B2(new_n912), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n937), .B(new_n938), .C1(new_n940), .C2(KEYINPUT39), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n913), .A2(new_n914), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n706), .A2(new_n727), .A3(new_n849), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n845), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n942), .A2(new_n916), .A3(new_n944), .ZN(new_n945));
  OR3_X1    g0745(.A1(new_n713), .A2(new_n712), .A3(new_n726), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n941), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n719), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(new_n529), .B2(new_n755), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n947), .B(new_n949), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n936), .A2(new_n950), .B1(new_n267), .B2(new_n721), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n951), .B(KEYINPUT107), .Z(new_n952));
  AND2_X1   g0752(.A1(new_n936), .A2(new_n950), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n877), .B(new_n881), .C1(new_n952), .C2(new_n953), .ZN(G367));
  INV_X1    g0754(.A(new_n779), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n787), .B1(new_n209), .B2(new_n340), .C1(new_n955), .C2(new_n245), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT110), .ZN(new_n957));
  INV_X1    g0757(.A(new_n792), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT111), .Z(new_n960));
  NAND2_X1  g0760(.A1(new_n689), .A2(new_n694), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n736), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n696), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n688), .B2(new_n962), .ZN(new_n964));
  INV_X1    g0764(.A(new_n802), .ZN(new_n965));
  AOI22_X1  g0765(.A1(G303), .A2(new_n795), .B1(new_n965), .B2(G283), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n825), .B2(new_n804), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n778), .B1(G317), .B2(new_n827), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n607), .B2(new_n800), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n967), .B(new_n969), .C1(G107), .C2(new_n815), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT112), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n971), .A2(KEYINPUT46), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n822), .A2(G116), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(KEYINPUT46), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(new_n973), .B2(new_n972), .ZN(new_n976));
  INV_X1    g0776(.A(G294), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n970), .B(new_n976), .C1(new_n977), .C2(new_n796), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n265), .B1(new_n800), .B2(new_n202), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT113), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n795), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n982), .A2(new_n295), .B1(new_n229), .B2(new_n802), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(G159), .B2(new_n797), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n979), .A2(new_n980), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n815), .A2(G68), .ZN(new_n986));
  AND4_X1   g0786(.A1(new_n981), .A2(new_n984), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n803), .A2(G143), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n822), .A2(new_n482), .B1(G137), .B2(new_n827), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(KEYINPUT114), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n989), .A2(KEYINPUT114), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n987), .A2(new_n988), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n978), .A2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT47), .Z(new_n994));
  INV_X1    g0794(.A(new_n786), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n960), .B1(new_n840), .B2(new_n964), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n741), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n639), .A2(new_n736), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n659), .A2(new_n663), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n659), .B2(new_n727), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n743), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT44), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1003), .A2(KEYINPUT109), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n743), .A2(new_n1000), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT45), .Z(new_n1007));
  OAI211_X1 g0807(.A(new_n1005), .B(new_n1007), .C1(KEYINPUT109), .C2(new_n1004), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n997), .B(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n735), .A2(new_n742), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n740), .B2(new_n742), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n733), .B(new_n1011), .Z(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n774), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1009), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n774), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n745), .B(KEYINPUT41), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n790), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1010), .A2(new_n999), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT42), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n659), .B1(new_n999), .B2(new_n739), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n727), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(KEYINPUT108), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT43), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1024), .A2(new_n1022), .A3(new_n964), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n1024), .B2(new_n964), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n997), .A2(new_n1000), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1026), .B(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n996), .B1(new_n1017), .B2(new_n1028), .ZN(G387));
  OR2_X1    g0829(.A1(new_n1012), .A2(new_n774), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1030), .A2(new_n745), .A3(new_n1013), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1012), .A2(new_n790), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n955), .B1(new_n242), .B2(G45), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(new_n746), .B2(new_n776), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n344), .A2(new_n229), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n746), .B1(new_n1035), .B2(KEYINPUT50), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1036), .B(new_n275), .C1(KEYINPUT50), .C2(new_n1035), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(G68), .B2(G77), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n1034), .A2(new_n1038), .B1(G107), .B2(new_n209), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n792), .B1(new_n1039), .B2(new_n787), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT115), .Z(new_n1041));
  AOI22_X1  g0841(.A1(G317), .A2(new_n795), .B1(new_n797), .B2(G311), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n855), .B2(new_n802), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(G322), .B2(new_n803), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT116), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n1045), .A2(KEYINPUT48), .B1(G283), .B2(new_n815), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(KEYINPUT48), .B2(new_n1045), .C1(new_n977), .C2(new_n821), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT49), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n491), .B1(new_n540), .B2(new_n800), .C1(new_n829), .C2(new_n807), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT117), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1049), .A2(new_n1052), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(G68), .A2(new_n965), .B1(new_n835), .B2(G97), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1056), .B1(new_n229), .B2(new_n982), .C1(new_n484), .C2(new_n804), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n491), .B(new_n1057), .C1(new_n308), .C2(new_n797), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n821), .A2(new_n202), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n683), .B2(new_n815), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1058), .B(new_n1060), .C1(new_n295), .C2(new_n807), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1055), .A2(new_n1061), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1041), .B1(new_n740), .B2(new_n840), .C1(new_n1062), .C2(new_n995), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1031), .A2(new_n1032), .A3(new_n1063), .ZN(G393));
  INV_X1    g0864(.A(new_n745), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1014), .A2(new_n1066), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n821), .A2(new_n231), .B1(new_n226), .B2(new_n800), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n491), .B(new_n1068), .C1(G143), .C2(new_n827), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1069), .A2(KEYINPUT118), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n797), .A2(G50), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n814), .A2(new_n202), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n795), .A2(G159), .B1(new_n803), .B2(G150), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT51), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n1072), .B(new_n1074), .C1(new_n344), .C2(new_n965), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1069), .A2(KEYINPUT118), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1070), .A2(new_n1071), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n795), .A2(G311), .B1(new_n803), .B2(G317), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1078), .A2(KEYINPUT52), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n822), .A2(G283), .B1(new_n815), .B2(G116), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n827), .A2(G322), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1081), .B1(new_n802), .B2(new_n977), .C1(new_n855), .C2(new_n796), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n1078), .B2(KEYINPUT52), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n265), .B1(new_n835), .B2(G107), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1080), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1077), .B1(new_n1079), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n792), .B1(new_n1086), .B2(new_n786), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n787), .B1(new_n607), .B2(new_n209), .C1(new_n955), .C2(new_n252), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1087), .B(new_n1088), .C1(new_n840), .C2(new_n1000), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n1009), .B2(new_n789), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1067), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(G390));
  AND3_X1   g0892(.A1(new_n386), .A2(new_n527), .A3(new_n524), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n527), .B1(new_n386), .B2(new_n524), .ZN(new_n1094));
  OAI211_X1 g0894(.A(G330), .B(new_n933), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n916), .B1(new_n773), .B2(new_n849), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n890), .A2(G330), .A3(new_n849), .A4(new_n889), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n916), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n944), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n752), .A2(new_n847), .B1(new_n368), .B2(new_n727), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n773), .A2(new_n849), .A3(new_n916), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1100), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n755), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1095), .A2(new_n1105), .A3(new_n1106), .A4(new_n719), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(KEYINPUT119), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT119), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n949), .A2(new_n1109), .A3(new_n1095), .A4(new_n1105), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT39), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n929), .B2(new_n930), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n937), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n1101), .B2(new_n1098), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1112), .A2(new_n1114), .A3(new_n938), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n940), .B(new_n1113), .C1(new_n1098), .C2(new_n1101), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1102), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1115), .B(new_n1116), .C1(new_n1098), .C2(new_n1097), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1108), .A2(new_n1110), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1108), .A2(new_n1110), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1122), .A2(new_n745), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(KEYINPUT120), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n789), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n821), .A2(new_n295), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT53), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n358), .B1(new_n835), .B2(G50), .ZN(new_n1129));
  INV_X1    g0929(.A(G128), .ZN(new_n1130));
  INV_X1    g0930(.A(G132), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1129), .B1(new_n804), .B2(new_n1130), .C1(new_n1131), .C2(new_n982), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(G159), .B2(new_n815), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n827), .A2(G125), .ZN(new_n1134));
  XOR2_X1   g0934(.A(KEYINPUT54), .B(G143), .Z(new_n1135));
  AOI22_X1  g0935(.A1(new_n797), .A2(G137), .B1(new_n965), .B2(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT121), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1128), .A2(new_n1133), .A3(new_n1134), .A4(new_n1137), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n358), .B1(new_n807), .B2(new_n977), .C1(new_n800), .C2(new_n231), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n804), .A2(new_n853), .B1(new_n607), .B2(new_n802), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1139), .B(new_n1140), .C1(G116), .C2(new_n795), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1072), .B1(G87), .B2(new_n822), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(new_n537), .C2(new_n796), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n1138), .A2(new_n1143), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n958), .B1(new_n308), .B2(new_n871), .C1(new_n1144), .C2(new_n995), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT122), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1112), .A2(new_n938), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1146), .B1(new_n1147), .B2(new_n783), .ZN(new_n1148));
  OAI21_X1  g0948(.A(KEYINPUT123), .B1(new_n1126), .B2(new_n1148), .ZN(new_n1149));
  OR3_X1    g0949(.A1(new_n1126), .A2(KEYINPUT123), .A3(new_n1148), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT120), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1122), .A2(new_n1151), .A3(new_n745), .A4(new_n1123), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1125), .A2(new_n1149), .A3(new_n1150), .A4(new_n1152), .ZN(G378));
  NAND3_X1  g0953(.A1(new_n1095), .A2(new_n719), .A3(new_n1106), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n311), .A2(new_n726), .ZN(new_n1155));
  XOR2_X1   g0955(.A(new_n1155), .B(KEYINPUT56), .Z(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT55), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n718), .B2(new_n376), .ZN(new_n1159));
  AOI211_X1 g0959(.A(KEYINPUT55), .B(new_n377), .C1(new_n716), .C2(new_n717), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1157), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n383), .A2(new_n715), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n339), .A2(KEYINPUT97), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n376), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(KEYINPUT55), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n718), .A2(new_n1158), .A3(new_n376), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1165), .A2(new_n1166), .A3(new_n1156), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1161), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(G330), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1168), .B1(new_n932), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1161), .A2(new_n1167), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT40), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n918), .A2(new_n893), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n924), .A2(KEYINPUT37), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n895), .A2(new_n896), .A3(new_n898), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT37), .A4(new_n895), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n920), .B2(new_n919), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n914), .B1(new_n1179), .B2(KEYINPUT38), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1172), .B1(new_n1173), .B2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1171), .B(G330), .C1(new_n1181), .C2(new_n915), .ZN(new_n1182));
  AND3_X1   g0982(.A1(new_n1170), .A2(new_n947), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n947), .B1(new_n1170), .B2(new_n1182), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n1121), .A2(new_n1154), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT57), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n745), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(KEYINPUT125), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT125), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1190), .B(new_n745), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1188), .A2(new_n1189), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1168), .A2(new_n783), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n965), .A2(G137), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n803), .A2(G125), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n1131), .B2(new_n796), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1194), .B(new_n1196), .C1(new_n822), .C2(new_n1135), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1197), .B1(new_n1130), .B2(new_n982), .C1(new_n295), .C2(new_n814), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT59), .Z(new_n1199));
  AOI21_X1  g0999(.A(G41), .B1(new_n835), .B2(G159), .ZN(new_n1200));
  AOI21_X1  g1000(.A(G33), .B1(new_n827), .B2(G124), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(G41), .B1(new_n778), .B2(G33), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1202), .B1(G50), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n683), .A2(new_n965), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n827), .A2(G283), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n986), .A2(new_n274), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(G97), .A2(new_n797), .B1(new_n835), .B2(new_n482), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n537), .B2(new_n982), .C1(new_n540), .C2(new_n804), .ZN(new_n1209));
  NOR4_X1   g1009(.A1(new_n1207), .A2(new_n1209), .A3(new_n778), .A4(new_n1059), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT58), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n786), .B1(new_n1204), .B2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n791), .B1(G50), .B2(new_n871), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT124), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1193), .A2(new_n1212), .A3(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1215), .B1(new_n1216), .B2(new_n789), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1192), .A2(new_n1218), .ZN(G375));
  NAND2_X1  g1019(.A1(new_n1105), .A2(new_n790), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n358), .B1(new_n807), .B2(new_n855), .C1(new_n800), .C2(new_n202), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n982), .A2(new_n853), .B1(new_n804), .B2(new_n977), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n1221), .B(new_n1222), .C1(G116), .C2(new_n797), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n815), .A2(new_n683), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n965), .A2(G107), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n822), .A2(G97), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n822), .A2(G159), .B1(new_n815), .B2(G50), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n795), .A2(G137), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n965), .A2(G150), .B1(new_n827), .B2(G128), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n803), .A2(G132), .B1(new_n797), .B2(new_n1135), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .A4(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n491), .B1(new_n482), .B2(new_n835), .ZN(new_n1233));
  XOR2_X1   g1033(.A(new_n1233), .B(KEYINPUT126), .Z(new_n1234));
  OAI21_X1  g1034(.A(new_n1227), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n792), .B1(new_n1235), .B2(new_n786), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(G68), .B2(new_n871), .C1(new_n916), .C2(new_n784), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1220), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1105), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1154), .A2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1108), .A2(new_n1110), .A3(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1016), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1239), .B1(new_n1242), .B2(new_n1243), .ZN(G381));
  INV_X1    g1044(.A(G375), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1126), .A2(new_n1148), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1124), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1248));
  OR4_X1    g1048(.A1(G396), .A2(G381), .A3(G384), .A4(G393), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1091), .B(new_n996), .C1(new_n1017), .C2(new_n1028), .ZN(new_n1250));
  OR3_X1    g1050(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .ZN(G407));
  OAI211_X1 g1051(.A(G407), .B(G213), .C1(G343), .C2(new_n1248), .ZN(G409));
  INV_X1    g1052(.A(G213), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1253), .A2(G343), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1192), .A2(G378), .A3(new_n1218), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1185), .A2(new_n1243), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1247), .B1(new_n1256), .B2(new_n1217), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1254), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  AND2_X1   g1058(.A1(new_n1254), .A2(G2897), .ZN(new_n1259));
  INV_X1    g1059(.A(G384), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT60), .B1(new_n1154), .B2(new_n1240), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n1065), .B(new_n1261), .C1(new_n1242), .C2(KEYINPUT60), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1260), .B1(new_n1262), .B2(new_n1238), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1242), .A2(KEYINPUT60), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1261), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1264), .A2(new_n745), .A3(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1266), .A2(G384), .A3(new_n1239), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1263), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT127), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1259), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1268), .A2(new_n1269), .A3(new_n1259), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(KEYINPUT63), .B1(new_n1258), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1268), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1258), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1278));
  AND2_X1   g1078(.A1(G387), .A2(G390), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1250), .ZN(new_n1280));
  XOR2_X1   g1080(.A(G393), .B(G396), .Z(new_n1281));
  OR3_X1    g1081(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1281), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  AOI211_X1 g1084(.A(new_n1254), .B(new_n1268), .C1(new_n1255), .C2(new_n1257), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1284), .B1(new_n1285), .B2(KEYINPUT63), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT61), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1278), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT62), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1258), .A2(new_n1289), .A3(new_n1276), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1287), .B1(new_n1258), .B2(new_n1274), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1289), .B1(new_n1258), .B2(new_n1276), .ZN(new_n1292));
  NOR3_X1   g1092(.A1(new_n1290), .A2(new_n1291), .A3(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1284), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1288), .B1(new_n1293), .B2(new_n1294), .ZN(G405));
  NAND2_X1  g1095(.A1(G375), .A2(new_n1247), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1255), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1276), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1296), .A2(new_n1255), .A3(new_n1268), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  XNOR2_X1  g1100(.A(new_n1300), .B(new_n1284), .ZN(G402));
endmodule


