//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 1 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n815, new_n817, new_n818, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT12), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G229gat), .A2(G233gat), .ZN(new_n208));
  XOR2_X1   g007(.A(new_n208), .B(KEYINPUT13), .Z(new_n209));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT83), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT14), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n211), .B(new_n212), .C1(G29gat), .C2(G36gat), .ZN(new_n213));
  INV_X1    g012(.A(G29gat), .ZN(new_n214));
  INV_X1    g013(.A(G36gat), .ZN(new_n215));
  OAI221_X1 g014(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n210), .C2(KEYINPUT15), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(KEYINPUT83), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n211), .B1(G29gat), .B2(G36gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT14), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  OAI211_X1 g019(.A(KEYINPUT15), .B(new_n210), .C1(new_n216), .C2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n210), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT15), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n222), .A2(new_n223), .B1(G29gat), .B2(G36gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n210), .A2(KEYINPUT15), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n224), .A2(new_n225), .A3(new_n219), .A4(new_n213), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n221), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G15gat), .B(G22gat), .ZN(new_n228));
  INV_X1    g027(.A(G1gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT16), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT84), .B1(new_n228), .B2(G1gat), .ZN(new_n233));
  OAI21_X1  g032(.A(G8gat), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  XOR2_X1   g033(.A(G15gat), .B(G22gat), .Z(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(new_n229), .ZN(new_n236));
  INV_X1    g035(.A(G8gat), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n236), .A2(new_n231), .A3(KEYINPUT84), .A4(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n227), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n227), .A2(new_n239), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n209), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT87), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n227), .B(new_n239), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT87), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n244), .A2(new_n245), .A3(new_n209), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n227), .A2(new_n239), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n208), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n239), .A2(KEYINPUT85), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT85), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n234), .A2(new_n251), .A3(new_n238), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT17), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n227), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n221), .A2(new_n226), .A3(KEYINPUT17), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT86), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n221), .A2(KEYINPUT17), .A3(new_n226), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT17), .B1(new_n221), .B2(new_n226), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n262), .A2(KEYINPUT86), .A3(new_n253), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n249), .B1(new_n259), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n247), .B1(new_n264), .B2(KEYINPUT18), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT18), .ZN(new_n266));
  AOI211_X1 g065(.A(new_n266), .B(new_n249), .C1(new_n259), .C2(new_n263), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n207), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n249), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n257), .A2(new_n258), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT86), .B1(new_n262), .B2(new_n253), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(new_n266), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n264), .A2(KEYINPUT18), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n273), .A2(new_n274), .A3(new_n206), .A4(new_n247), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n268), .A2(new_n275), .A3(KEYINPUT88), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT88), .B1(new_n268), .B2(new_n275), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G113gat), .B(G120gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT71), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT1), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(KEYINPUT72), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G127gat), .ZN(new_n284));
  INV_X1    g083(.A(G134gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(G127gat), .A2(G134gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n283), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n290));
  OAI21_X1  g089(.A(KEYINPUT71), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n280), .A2(KEYINPUT1), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT69), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT68), .B(KEYINPUT26), .ZN(new_n296));
  NOR2_X1   g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n295), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT68), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n300), .A2(KEYINPUT26), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT26), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(KEYINPUT68), .ZN(new_n303));
  OAI211_X1 g102(.A(KEYINPUT69), .B(new_n297), .C1(new_n301), .C2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G169gat), .ZN(new_n305));
  INV_X1    g104(.A(G176gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n302), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(new_n298), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n299), .A2(new_n304), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT70), .ZN(new_n310));
  NAND2_X1  g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311));
  AND3_X1   g110(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n310), .B1(new_n309), .B2(new_n311), .ZN(new_n313));
  XOR2_X1   g112(.A(KEYINPUT27), .B(G183gat), .Z(new_n314));
  OAI21_X1  g113(.A(KEYINPUT28), .B1(new_n314), .B2(G190gat), .ZN(new_n315));
  INV_X1    g114(.A(G183gat), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT27), .B1(new_n316), .B2(KEYINPUT67), .ZN(new_n317));
  NOR2_X1   g116(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n318));
  OR2_X1    g117(.A1(new_n316), .A2(KEYINPUT27), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n317), .B(new_n318), .C1(KEYINPUT67), .C2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  NOR3_X1   g120(.A1(new_n312), .A2(new_n313), .A3(new_n321), .ZN(new_n322));
  OAI22_X1  g121(.A1(new_n311), .A2(KEYINPUT24), .B1(new_n305), .B2(new_n306), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(G190gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n316), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n326), .A2(KEYINPUT24), .A3(new_n311), .ZN(new_n327));
  OR2_X1    g126(.A1(new_n297), .A2(KEYINPUT23), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT25), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n329), .B1(new_n297), .B2(KEYINPUT23), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n324), .A2(new_n327), .A3(new_n328), .A4(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT66), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n297), .A2(KEYINPUT23), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n323), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT66), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n334), .A2(new_n335), .A3(new_n327), .A4(new_n330), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT23), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT65), .B1(new_n298), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT65), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n297), .A2(new_n339), .A3(KEYINPUT23), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n334), .A2(new_n327), .A3(new_n338), .A4(new_n340), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n332), .A2(new_n336), .B1(new_n341), .B2(new_n329), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n294), .B1(new_n322), .B2(new_n342), .ZN(new_n343));
  AOI22_X1  g142(.A1(new_n283), .A2(new_n288), .B1(new_n291), .B2(new_n292), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n332), .A2(new_n336), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n341), .A2(new_n329), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n321), .ZN(new_n348));
  INV_X1    g147(.A(new_n311), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n297), .B1(new_n301), .B2(new_n303), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n350), .A2(new_n295), .B1(new_n298), .B2(new_n307), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n349), .B1(new_n351), .B2(new_n304), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n348), .B1(new_n352), .B2(new_n310), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n344), .B(new_n347), .C1(new_n353), .C2(new_n312), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n343), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G227gat), .A2(G233gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n356), .B(KEYINPUT64), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT73), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n357), .A3(new_n354), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT32), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n357), .B1(new_n343), .B2(new_n354), .ZN(new_n363));
  OAI211_X1 g162(.A(KEYINPUT32), .B(new_n360), .C1(new_n363), .C2(KEYINPUT73), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT33), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n360), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G15gat), .B(G43gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(G71gat), .B(G99gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n368), .B(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT34), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n370), .B1(new_n360), .B2(new_n366), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT34), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n365), .A2(new_n371), .A3(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n372), .A2(new_n373), .ZN(new_n376));
  AOI211_X1 g175(.A(KEYINPUT34), .B(new_n370), .C1(new_n360), .C2(new_n366), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n364), .B(new_n362), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT36), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n375), .A2(new_n378), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT36), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(G226gat), .A2(G233gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n309), .A2(new_n311), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n321), .B1(new_n386), .B2(KEYINPUT70), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n352), .A2(new_n310), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n342), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n385), .B1(new_n389), .B2(KEYINPUT29), .ZN(new_n390));
  XNOR2_X1  g189(.A(G197gat), .B(G204gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(G211gat), .A2(G218gat), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT22), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(G211gat), .B(G218gat), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n391), .A3(new_n394), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n347), .B1(new_n353), .B2(new_n312), .ZN(new_n401));
  INV_X1    g200(.A(new_n385), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n390), .A2(new_n400), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n400), .B1(new_n390), .B2(new_n403), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT37), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n400), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT29), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n402), .B1(new_n401), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n389), .A2(new_n385), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n407), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT37), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n390), .A2(new_n403), .A3(new_n400), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G8gat), .B(G36gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(G64gat), .B(G92gat), .ZN(new_n416));
  XOR2_X1   g215(.A(new_n415), .B(new_n416), .Z(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n406), .A2(new_n414), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT38), .ZN(new_n420));
  OR2_X1    g219(.A1(G141gat), .A2(G148gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(G141gat), .A2(G148gat), .ZN(new_n422));
  AND2_X1   g221(.A1(G155gat), .A2(G162gat), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT2), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n421), .B(new_n422), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  OR2_X1    g224(.A1(new_n423), .A2(KEYINPUT74), .ZN(new_n426));
  NOR2_X1   g225(.A1(G155gat), .A2(G162gat), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT74), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n425), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  XOR2_X1   g228(.A(KEYINPUT75), .B(G155gat), .Z(new_n430));
  AOI21_X1  g229(.A(new_n424), .B1(new_n430), .B2(G162gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(G155gat), .B(G162gat), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n432), .A2(new_n421), .A3(new_n422), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n429), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT3), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT3), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n429), .B(new_n436), .C1(new_n431), .C2(new_n433), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n435), .A2(new_n344), .A3(new_n437), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n426), .A2(new_n428), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n432), .A2(new_n421), .A3(new_n422), .ZN(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT75), .B(G155gat), .ZN(new_n441));
  INV_X1    g240(.A(G162gat), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT2), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n439), .A2(new_n425), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n294), .A2(KEYINPUT4), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(G225gat), .A2(G233gat), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT4), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n447), .B1(new_n344), .B2(new_n434), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n438), .A2(new_n445), .A3(new_n446), .A4(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT5), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n294), .A2(new_n444), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n344), .A2(new_n434), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n446), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n449), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n445), .A2(new_n448), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n455), .A2(KEYINPUT5), .A3(new_n446), .A4(new_n438), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT81), .ZN(new_n458));
  XOR2_X1   g257(.A(G1gat), .B(G29gat), .Z(new_n459));
  XNOR2_X1  g258(.A(G57gat), .B(G85gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n459), .B(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n461), .B(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT81), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n454), .A2(new_n456), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n458), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n463), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT6), .B1(new_n457), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n457), .A2(new_n467), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n466), .A2(new_n468), .B1(KEYINPUT6), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT38), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n406), .A2(new_n414), .A3(new_n471), .A4(new_n418), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n411), .A2(new_n413), .A3(new_n417), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n420), .A2(new_n470), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(G78gat), .B(G106gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(KEYINPUT31), .B(G50gat), .ZN(new_n476));
  XOR2_X1   g275(.A(new_n475), .B(new_n476), .Z(new_n477));
  INV_X1    g276(.A(G22gat), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n400), .B1(new_n437), .B2(new_n408), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n400), .A2(new_n408), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(new_n436), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n434), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT78), .ZN(new_n484));
  NAND2_X1  g283(.A1(G228gat), .A2(G233gat), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n480), .B(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  OAI211_X1 g286(.A(G228gat), .B(G233gat), .C1(new_n479), .C2(KEYINPUT78), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n444), .B1(new_n481), .B2(new_n436), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n489), .A2(new_n479), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n478), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT80), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n477), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT79), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n495), .B1(new_n487), .B2(new_n491), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n485), .B1(new_n480), .B2(new_n484), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n483), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(KEYINPUT79), .A3(new_n486), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n496), .A2(new_n500), .A3(G22gat), .ZN(new_n501));
  AOI21_X1  g300(.A(G22gat), .B1(new_n499), .B2(new_n486), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT80), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n494), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  NOR3_X1   g303(.A1(new_n487), .A2(new_n491), .A3(new_n478), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n477), .B1(new_n505), .B2(new_n502), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n438), .A2(new_n448), .A3(new_n445), .ZN(new_n508));
  OR3_X1    g307(.A1(new_n508), .A2(KEYINPUT39), .A3(new_n446), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n451), .A2(new_n452), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(new_n446), .ZN(new_n511));
  OAI211_X1 g310(.A(KEYINPUT39), .B(new_n511), .C1(new_n508), .C2(new_n446), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n509), .A2(new_n512), .A3(KEYINPUT40), .A4(new_n467), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT82), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n509), .A2(new_n467), .A3(new_n512), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT40), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n515), .A2(new_n466), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n418), .B1(new_n404), .B2(new_n405), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n520), .A2(KEYINPUT30), .A3(new_n473), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT30), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n411), .A2(new_n522), .A3(new_n413), .A4(new_n417), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n474), .B(new_n507), .C1(new_n519), .C2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT77), .B1(new_n457), .B2(new_n467), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT77), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n454), .A2(new_n456), .A3(new_n527), .A4(new_n463), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n526), .A2(new_n468), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n469), .A2(KEYINPUT6), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n524), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n507), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n384), .A2(new_n525), .A3(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n470), .A2(KEYINPUT35), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n379), .A2(new_n507), .A3(new_n536), .A4(new_n524), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n507), .A2(new_n375), .A3(new_n378), .ZN(new_n538));
  OAI21_X1  g337(.A(KEYINPUT35), .B1(new_n538), .B2(new_n532), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n279), .B1(new_n535), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT90), .ZN(new_n542));
  XNOR2_X1  g341(.A(G57gat), .B(G64gat), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT89), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AND2_X1   g344(.A1(G71gat), .A2(G78gat), .ZN(new_n546));
  NOR2_X1   g345(.A1(G71gat), .A2(G78gat), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n546), .A2(new_n547), .ZN(new_n550));
  OR2_X1    g349(.A1(G57gat), .A2(G64gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(G57gat), .A2(G64gat), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n551), .B(new_n552), .C1(new_n546), .C2(KEYINPUT9), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n550), .B1(new_n553), .B2(KEYINPUT89), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n542), .B1(new_n549), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n545), .A2(new_n548), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n553), .A2(new_n550), .A3(KEYINPUT89), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT90), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n559), .A2(KEYINPUT21), .ZN(new_n560));
  NAND2_X1  g359(.A1(G231gat), .A2(G233gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(G127gat), .ZN(new_n563));
  XOR2_X1   g362(.A(G183gat), .B(G211gat), .Z(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n562), .B(new_n284), .ZN(new_n566));
  INV_X1    g365(.A(new_n564), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n239), .B1(new_n559), .B2(KEYINPUT21), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT91), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(G155gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n571), .B(new_n573), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n569), .A2(new_n574), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G85gat), .A2(G92gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT7), .ZN(new_n579));
  XOR2_X1   g378(.A(G99gat), .B(G106gat), .Z(new_n580));
  NOR2_X1   g379(.A1(G85gat), .A2(G92gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(G99gat), .A2(G106gat), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n581), .B1(KEYINPUT8), .B2(new_n582), .ZN(new_n583));
  AND3_X1   g382(.A1(new_n579), .A2(new_n580), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n580), .B1(new_n579), .B2(new_n583), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n262), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT94), .ZN(new_n589));
  NAND2_X1  g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT92), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT41), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n586), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n593), .B1(new_n227), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n587), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n588), .A2(KEYINPUT94), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n596), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n591), .A2(new_n592), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n600), .B(KEYINPUT93), .Z(new_n601));
  XNOR2_X1  g400(.A(G134gat), .B(G162gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n599), .B(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(KEYINPUT95), .B1(new_n577), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT95), .ZN(new_n606));
  INV_X1    g405(.A(new_n604), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n575), .A2(new_n606), .A3(new_n576), .A4(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(G230gat), .ZN(new_n609));
  INV_X1    g408(.A(G233gat), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n555), .A2(new_n558), .A3(new_n586), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT96), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT96), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n555), .A2(new_n586), .A3(new_n614), .A4(new_n558), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT10), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT97), .B1(new_n579), .B2(new_n583), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  OAI22_X1  g418(.A1(new_n619), .A2(new_n580), .B1(new_n549), .B2(new_n554), .ZN(new_n620));
  NOR3_X1   g419(.A1(new_n584), .A2(new_n585), .A3(new_n618), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n616), .A2(new_n617), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n559), .A2(KEYINPUT10), .A3(new_n594), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n611), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI211_X1 g425(.A(new_n609), .B(new_n610), .C1(new_n616), .C2(new_n623), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G120gat), .B(G148gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(G176gat), .B(G204gat), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n629), .B(new_n630), .Z(new_n631));
  NAND2_X1  g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n631), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n633), .B1(new_n626), .B2(new_n627), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n634), .A3(KEYINPUT98), .ZN(new_n635));
  OR3_X1    g434(.A1(new_n628), .A2(KEYINPUT98), .A3(new_n631), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n605), .A2(new_n608), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n541), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n639), .A2(new_n531), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(new_n229), .ZN(G1324gat));
  INV_X1    g440(.A(new_n639), .ZN(new_n642));
  INV_X1    g441(.A(new_n524), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n237), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT16), .B(G8gat), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n639), .A2(new_n524), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(KEYINPUT42), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n647), .B1(KEYINPUT42), .B2(new_n646), .ZN(G1325gat));
  OAI21_X1  g447(.A(G15gat), .B1(new_n639), .B2(new_n384), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n381), .A2(G15gat), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n649), .B1(new_n639), .B2(new_n650), .ZN(G1326gat));
  NOR2_X1   g450(.A1(new_n639), .A2(new_n507), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT43), .B(G22gat), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(G1327gat));
  INV_X1    g453(.A(new_n577), .ZN(new_n655));
  INV_X1    g454(.A(new_n637), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n655), .A2(new_n607), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n541), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n531), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n659), .A2(new_n214), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT99), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT45), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT101), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n537), .A2(new_n539), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n665), .B1(new_n537), .B2(new_n539), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n535), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(KEYINPUT102), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT102), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n535), .B(new_n670), .C1(new_n666), .C2(new_n667), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n607), .A2(KEYINPUT44), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n669), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n535), .A2(new_n540), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT44), .B1(new_n674), .B2(new_n607), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n268), .A2(new_n275), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n577), .A2(new_n677), .A3(new_n637), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT100), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(G29gat), .B1(new_n680), .B2(new_n531), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n662), .A2(new_n663), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n664), .A2(new_n681), .A3(new_n682), .ZN(G1328gat));
  NOR3_X1   g482(.A1(new_n658), .A2(G36gat), .A3(new_n524), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT46), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n680), .A2(new_n524), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n685), .B1(new_n686), .B2(new_n215), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1329gat));
  AOI21_X1  g488(.A(G43gat), .B1(new_n659), .B2(new_n379), .ZN(new_n690));
  INV_X1    g489(.A(new_n680), .ZN(new_n691));
  INV_X1    g490(.A(new_n384), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n692), .A2(G43gat), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n690), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n694), .B(KEYINPUT47), .Z(G1330gat));
  NAND2_X1  g494(.A1(new_n659), .A2(KEYINPUT104), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT104), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n507), .B1(new_n658), .B2(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(G50gat), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n533), .A2(G50gat), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n699), .B1(new_n691), .B2(new_n700), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n701), .B(KEYINPUT48), .Z(G1331gat));
  AND2_X1   g501(.A1(new_n669), .A2(new_n671), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n637), .A2(new_n677), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n605), .A2(new_n608), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n660), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(G57gat), .ZN(G1332gat));
  OAI22_X1  g508(.A1(new_n706), .A2(new_n524), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n707), .A2(new_n643), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT49), .B(G64gat), .Z(new_n712));
  OAI21_X1  g511(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT105), .ZN(G1333gat));
  INV_X1    g513(.A(G71gat), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n715), .B1(new_n706), .B2(new_n381), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT106), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n384), .A2(new_n715), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n717), .B1(new_n707), .B2(new_n718), .ZN(new_n719));
  NOR4_X1   g518(.A1(new_n706), .A2(KEYINPUT106), .A3(new_n715), .A4(new_n384), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n716), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(KEYINPUT50), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT50), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n723), .B(new_n716), .C1(new_n719), .C2(new_n720), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(G1334gat));
  NOR2_X1   g524(.A1(new_n706), .A2(new_n507), .ZN(new_n726));
  XOR2_X1   g525(.A(KEYINPUT107), .B(G78gat), .Z(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1335gat));
  INV_X1    g527(.A(KEYINPUT51), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n540), .A2(KEYINPUT101), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n537), .A2(new_n539), .A3(new_n665), .ZN(new_n731));
  AOI22_X1  g530(.A1(new_n380), .A2(new_n383), .B1(new_n533), .B2(new_n532), .ZN(new_n732));
  AOI22_X1  g531(.A1(new_n730), .A2(new_n731), .B1(new_n525), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n655), .A2(new_n607), .ZN(new_n734));
  INV_X1    g533(.A(new_n677), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n729), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT108), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n668), .A2(KEYINPUT51), .A3(new_n735), .A4(new_n734), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  OAI211_X1 g539(.A(KEYINPUT108), .B(new_n729), .C1(new_n733), .C2(new_n736), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OR4_X1    g541(.A1(G85gat), .A2(new_n742), .A3(new_n531), .A4(new_n637), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n577), .A2(new_n704), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n676), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(G85gat), .B1(new_n746), .B2(new_n531), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n743), .A2(new_n747), .ZN(G1336gat));
  OAI21_X1  g547(.A(G92gat), .B1(new_n746), .B2(new_n524), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n524), .A2(G92gat), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n740), .A2(new_n656), .A3(new_n741), .A4(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n739), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n754), .A2(new_n656), .A3(new_n751), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n749), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n753), .B1(new_n756), .B2(new_n750), .ZN(G1337gat));
  OAI21_X1  g556(.A(G99gat), .B1(new_n746), .B2(new_n384), .ZN(new_n758));
  OR3_X1    g557(.A1(new_n637), .A2(new_n381), .A3(G99gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n758), .B1(new_n742), .B2(new_n759), .ZN(G1338gat));
  INV_X1    g559(.A(KEYINPUT53), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n507), .A2(G106gat), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n740), .A2(new_n656), .A3(new_n741), .A4(new_n762), .ZN(new_n763));
  AOI211_X1 g562(.A(new_n507), .B(new_n744), .C1(new_n673), .C2(new_n675), .ZN(new_n764));
  INV_X1    g563(.A(G106gat), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n761), .B(new_n763), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n676), .A2(new_n533), .A3(new_n745), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n637), .B1(new_n737), .B2(new_n739), .ZN(new_n768));
  AOI22_X1  g567(.A1(new_n767), .A2(G106gat), .B1(new_n768), .B2(new_n762), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n766), .B1(new_n769), .B2(new_n761), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT109), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT109), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n766), .B(new_n772), .C1(new_n769), .C2(new_n761), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(G1339gat));
  AOI211_X1 g573(.A(KEYINPUT10), .B(new_n622), .C1(new_n613), .C2(new_n615), .ZN(new_n775));
  INV_X1    g574(.A(new_n625), .ZN(new_n776));
  OAI22_X1  g575(.A1(new_n775), .A2(new_n776), .B1(new_n609), .B2(new_n610), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n624), .A2(new_n611), .A3(new_n625), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n777), .A2(new_n778), .A3(KEYINPUT54), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n631), .B1(new_n626), .B2(new_n780), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  AOI22_X1  g581(.A1(new_n782), .A2(KEYINPUT55), .B1(new_n628), .B2(new_n631), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT110), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n782), .B2(KEYINPUT55), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n779), .A2(new_n781), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n786), .A2(KEYINPUT110), .A3(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n783), .A2(new_n785), .A3(new_n677), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n259), .A2(new_n263), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n208), .B1(new_n790), .B2(new_n248), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n244), .A2(new_n209), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n205), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n275), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n656), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n604), .B1(new_n789), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n783), .A2(new_n785), .A3(new_n788), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n795), .A2(new_n604), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n577), .B1(new_n797), .B2(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n605), .A2(new_n735), .A3(new_n608), .A4(new_n637), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n531), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AND4_X1   g602(.A1(new_n507), .A2(new_n803), .A3(new_n524), .A4(new_n379), .ZN(new_n804));
  XOR2_X1   g603(.A(new_n804), .B(KEYINPUT111), .Z(new_n805));
  INV_X1    g604(.A(G113gat), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n805), .A2(new_n806), .A3(new_n677), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n533), .B1(new_n801), .B2(new_n802), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n643), .A2(new_n531), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n808), .A2(new_n379), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(G113gat), .B1(new_n810), .B2(new_n279), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n807), .A2(new_n811), .ZN(G1340gat));
  INV_X1    g611(.A(G120gat), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n805), .A2(new_n813), .A3(new_n656), .ZN(new_n814));
  OAI21_X1  g613(.A(G120gat), .B1(new_n810), .B2(new_n637), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(G1341gat));
  NAND3_X1  g615(.A1(new_n804), .A2(new_n284), .A3(new_n655), .ZN(new_n817));
  OAI21_X1  g616(.A(G127gat), .B1(new_n810), .B2(new_n577), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(G1342gat));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n285), .A3(new_n604), .ZN(new_n820));
  OR2_X1    g619(.A1(new_n820), .A2(KEYINPUT112), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(KEYINPUT112), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT56), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(G134gat), .B1(new_n810), .B2(new_n607), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n821), .A2(KEYINPUT56), .A3(new_n822), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(G1343gat));
  AND2_X1   g627(.A1(new_n384), .A2(new_n809), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n533), .A2(KEYINPUT57), .ZN(new_n830));
  OR2_X1    g629(.A1(new_n798), .A2(new_n799), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n786), .A2(KEYINPUT113), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n779), .A2(new_n781), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(new_n787), .A3(new_n834), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n835), .B(new_n783), .C1(new_n277), .C2(new_n278), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n604), .B1(new_n836), .B2(new_n796), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n831), .B1(new_n837), .B2(KEYINPUT114), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT114), .ZN(new_n839));
  AOI211_X1 g638(.A(new_n839), .B(new_n604), .C1(new_n836), .C2(new_n796), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n577), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n830), .B1(new_n841), .B2(new_n802), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n801), .A2(new_n802), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT57), .B1(new_n843), .B2(new_n533), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n677), .B(new_n829), .C1(new_n842), .C2(new_n844), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n845), .A2(KEYINPUT115), .A3(G141gat), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT115), .B1(new_n845), .B2(G141gat), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n692), .A2(new_n507), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n524), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n279), .A2(G141gat), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n803), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n846), .A2(new_n847), .A3(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n279), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n857), .B(new_n829), .C1(new_n842), .C2(new_n844), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n856), .B1(new_n858), .B2(G141gat), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI211_X1 g660(.A(KEYINPUT116), .B(new_n856), .C1(new_n858), .C2(G141gat), .ZN(new_n862));
  OAI22_X1  g661(.A1(new_n854), .A2(new_n855), .B1(new_n861), .B2(new_n862), .ZN(G1344gat));
  OAI21_X1  g662(.A(KEYINPUT118), .B1(new_n837), .B2(new_n800), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT118), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n637), .A2(new_n794), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n632), .B1(new_n786), .B2(new_n787), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT88), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n677), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n867), .B1(new_n869), .B2(new_n276), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n866), .B1(new_n870), .B2(new_n835), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n831), .B(new_n865), .C1(new_n871), .C2(new_n604), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n864), .A2(new_n872), .A3(new_n577), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n638), .A2(new_n279), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT57), .B1(new_n875), .B2(new_n533), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n830), .B1(new_n801), .B2(new_n802), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n829), .A2(new_n879), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n829), .A2(new_n879), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n878), .A2(new_n656), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  AND2_X1   g681(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n803), .A2(new_n850), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n637), .A2(G148gat), .ZN(new_n885));
  AOI22_X1  g684(.A1(new_n882), .A2(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n829), .B1(new_n842), .B2(new_n844), .ZN(new_n887));
  OAI21_X1  g686(.A(G148gat), .B1(new_n887), .B2(new_n637), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n886), .A2(new_n890), .ZN(G1345gat));
  OAI21_X1  g690(.A(new_n430), .B1(new_n887), .B2(new_n577), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n884), .A2(new_n441), .A3(new_n655), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(G1346gat));
  OR3_X1    g693(.A1(new_n887), .A2(new_n442), .A3(new_n607), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(G162gat), .B1(new_n884), .B2(new_n604), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n896), .A2(new_n897), .ZN(G1347gat));
  NOR3_X1   g697(.A1(new_n381), .A2(new_n660), .A3(new_n524), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n808), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n305), .B1(new_n900), .B2(new_n857), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n660), .B1(new_n801), .B2(new_n802), .ZN(new_n902));
  AND4_X1   g701(.A1(new_n507), .A2(new_n902), .A3(new_n643), .A4(new_n379), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n735), .A2(G169gat), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n901), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT119), .ZN(G1348gat));
  AOI21_X1  g705(.A(G176gat), .B1(new_n903), .B2(new_n656), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n637), .A2(new_n306), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n900), .B2(new_n908), .ZN(G1349gat));
  INV_X1    g708(.A(KEYINPUT120), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n900), .A2(new_n655), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n577), .A2(new_n314), .ZN(new_n912));
  AOI22_X1  g711(.A1(new_n911), .A2(G183gat), .B1(new_n903), .B2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT121), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n910), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(KEYINPUT60), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT60), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n917), .B1(new_n913), .B2(new_n910), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n916), .B1(new_n915), .B2(new_n918), .ZN(G1350gat));
  NAND3_X1  g718(.A1(new_n903), .A2(new_n325), .A3(new_n604), .ZN(new_n920));
  XOR2_X1   g719(.A(new_n920), .B(KEYINPUT122), .Z(new_n921));
  AOI21_X1  g720(.A(new_n325), .B1(new_n900), .B2(new_n604), .ZN(new_n922));
  XOR2_X1   g721(.A(new_n922), .B(KEYINPUT61), .Z(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(G1351gat));
  NAND2_X1  g723(.A1(new_n848), .A2(new_n643), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT123), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n902), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(G197gat), .B1(new_n928), .B2(new_n677), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n384), .A2(new_n531), .A3(new_n643), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT124), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n878), .A2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n857), .A2(G197gat), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n929), .B1(new_n933), .B2(new_n934), .ZN(G1352gat));
  NOR3_X1   g734(.A1(new_n927), .A2(G204gat), .A3(new_n637), .ZN(new_n936));
  XNOR2_X1  g735(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n936), .B(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(G204gat), .B1(new_n932), .B2(new_n637), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1353gat));
  OAI211_X1 g739(.A(new_n655), .B(new_n931), .C1(new_n876), .C2(new_n877), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G211gat), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT63), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n941), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n944), .A2(KEYINPUT126), .A3(new_n945), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n927), .A2(G211gat), .A3(new_n577), .ZN(new_n947));
  AOI21_X1  g746(.A(KEYINPUT63), .B1(new_n941), .B2(G211gat), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT126), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n946), .A2(new_n950), .ZN(G1354gat));
  AOI21_X1  g750(.A(KEYINPUT127), .B1(new_n878), .B2(new_n931), .ZN(new_n952));
  OAI211_X1 g751(.A(KEYINPUT127), .B(new_n931), .C1(new_n876), .C2(new_n877), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(new_n604), .ZN(new_n954));
  OAI21_X1  g753(.A(G218gat), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  OR3_X1    g754(.A1(new_n927), .A2(G218gat), .A3(new_n607), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1355gat));
endmodule


