

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589;

  NOR2_X1 U322 ( .A1(n413), .A2(n412), .ZN(n492) );
  INV_X1 U323 ( .A(KEYINPUT45), .ZN(n465) );
  INV_X1 U324 ( .A(KEYINPUT5), .ZN(n353) );
  XNOR2_X1 U325 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U326 ( .A(n356), .B(n355), .ZN(n360) );
  XNOR2_X1 U327 ( .A(n378), .B(n325), .ZN(n326) );
  XNOR2_X1 U328 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U329 ( .A(n327), .B(n326), .ZN(n329) );
  XNOR2_X1 U330 ( .A(n367), .B(n366), .ZN(n369) );
  NOR2_X1 U331 ( .A1(n524), .A2(n478), .ZN(n573) );
  INV_X1 U332 ( .A(G190GAT), .ZN(n485) );
  XNOR2_X1 U333 ( .A(n452), .B(KEYINPUT38), .ZN(n509) );
  XNOR2_X1 U334 ( .A(n485), .B(KEYINPUT58), .ZN(n486) );
  XNOR2_X1 U335 ( .A(n453), .B(G43GAT), .ZN(n454) );
  XNOR2_X1 U336 ( .A(n487), .B(n486), .ZN(G1351GAT) );
  XNOR2_X1 U337 ( .A(n455), .B(n454), .ZN(G1330GAT) );
  XOR2_X1 U338 ( .A(G127GAT), .B(G176GAT), .Z(n291) );
  XNOR2_X1 U339 ( .A(KEYINPUT86), .B(KEYINPUT87), .ZN(n290) );
  XNOR2_X1 U340 ( .A(n291), .B(n290), .ZN(n295) );
  XOR2_X1 U341 ( .A(G190GAT), .B(G134GAT), .Z(n293) );
  XOR2_X1 U342 ( .A(G43GAT), .B(G99GAT), .Z(n316) );
  XOR2_X1 U343 ( .A(G113GAT), .B(KEYINPUT0), .Z(n364) );
  XNOR2_X1 U344 ( .A(n316), .B(n364), .ZN(n292) );
  XNOR2_X1 U345 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U346 ( .A(n295), .B(n294), .Z(n297) );
  NAND2_X1 U347 ( .A1(G227GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U349 ( .A(G71GAT), .B(KEYINPUT91), .Z(n299) );
  XNOR2_X1 U350 ( .A(G15GAT), .B(G120GAT), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U352 ( .A(n301), .B(n300), .Z(n310) );
  XNOR2_X1 U353 ( .A(KEYINPUT19), .B(KEYINPUT88), .ZN(n302) );
  XNOR2_X1 U354 ( .A(n302), .B(KEYINPUT18), .ZN(n303) );
  XOR2_X1 U355 ( .A(n303), .B(KEYINPUT17), .Z(n305) );
  XNOR2_X1 U356 ( .A(G169GAT), .B(G183GAT), .ZN(n304) );
  XNOR2_X1 U357 ( .A(n305), .B(n304), .ZN(n382) );
  XOR2_X1 U358 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n307) );
  XNOR2_X1 U359 ( .A(KEYINPUT85), .B(KEYINPUT20), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U361 ( .A(n382), .B(n308), .ZN(n309) );
  XNOR2_X1 U362 ( .A(n310), .B(n309), .ZN(n538) );
  XOR2_X1 U363 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n312) );
  XNOR2_X1 U364 ( .A(KEYINPUT64), .B(KEYINPUT75), .ZN(n311) );
  XNOR2_X1 U365 ( .A(n312), .B(n311), .ZN(n320) );
  XOR2_X1 U366 ( .A(KEYINPUT10), .B(KEYINPUT77), .Z(n314) );
  XNOR2_X1 U367 ( .A(G92GAT), .B(KEYINPUT65), .ZN(n313) );
  XNOR2_X1 U368 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U369 ( .A(n315), .B(G106GAT), .Z(n318) );
  XNOR2_X1 U370 ( .A(n316), .B(G218GAT), .ZN(n317) );
  XNOR2_X1 U371 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U372 ( .A(n320), .B(n319), .ZN(n331) );
  XOR2_X1 U373 ( .A(G85GAT), .B(KEYINPUT76), .Z(n322) );
  XNOR2_X1 U374 ( .A(G29GAT), .B(G134GAT), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n356) );
  INV_X1 U376 ( .A(KEYINPUT74), .ZN(n323) );
  XNOR2_X1 U377 ( .A(n356), .B(n323), .ZN(n327) );
  XNOR2_X1 U378 ( .A(G36GAT), .B(G190GAT), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n324), .B(KEYINPUT78), .ZN(n378) );
  NAND2_X1 U380 ( .A1(G232GAT), .A2(G233GAT), .ZN(n325) );
  XOR2_X1 U381 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n420) );
  XOR2_X1 U382 ( .A(G50GAT), .B(G162GAT), .Z(n386) );
  XOR2_X1 U383 ( .A(n420), .B(n386), .Z(n328) );
  XNOR2_X1 U384 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U385 ( .A(n331), .B(n330), .ZN(n561) );
  INV_X1 U386 ( .A(n561), .ZN(n488) );
  XNOR2_X1 U387 ( .A(KEYINPUT36), .B(n488), .ZN(n586) );
  XOR2_X1 U388 ( .A(KEYINPUT13), .B(KEYINPUT70), .Z(n333) );
  XNOR2_X1 U389 ( .A(G71GAT), .B(KEYINPUT71), .ZN(n332) );
  XNOR2_X1 U390 ( .A(n333), .B(n332), .ZN(n444) );
  XOR2_X1 U391 ( .A(G1GAT), .B(G127GAT), .Z(n368) );
  XNOR2_X1 U392 ( .A(n444), .B(n368), .ZN(n335) );
  AND2_X1 U393 ( .A1(G231GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U394 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n336), .B(KEYINPUT80), .ZN(n340) );
  XOR2_X1 U396 ( .A(KEYINPUT68), .B(G8GAT), .Z(n338) );
  XNOR2_X1 U397 ( .A(G15GAT), .B(G22GAT), .ZN(n337) );
  XNOR2_X1 U398 ( .A(n338), .B(n337), .ZN(n424) );
  XOR2_X1 U399 ( .A(n424), .B(KEYINPUT79), .Z(n339) );
  XNOR2_X1 U400 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U401 ( .A(G78GAT), .B(G155GAT), .Z(n342) );
  XNOR2_X1 U402 ( .A(G183GAT), .B(G211GAT), .ZN(n341) );
  XOR2_X1 U403 ( .A(n342), .B(n341), .Z(n343) );
  XNOR2_X1 U404 ( .A(n344), .B(n343), .ZN(n352) );
  XOR2_X1 U405 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n346) );
  XNOR2_X1 U406 ( .A(KEYINPUT12), .B(KEYINPUT83), .ZN(n345) );
  XNOR2_X1 U407 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U408 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n348) );
  XNOR2_X1 U409 ( .A(G57GAT), .B(G64GAT), .ZN(n347) );
  XNOR2_X1 U410 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U411 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n352), .B(n351), .ZN(n558) );
  NAND2_X1 U413 ( .A1(G225GAT), .A2(G233GAT), .ZN(n354) );
  XOR2_X1 U414 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n358) );
  XNOR2_X1 U415 ( .A(G162GAT), .B(KEYINPUT6), .ZN(n357) );
  XNOR2_X1 U416 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U417 ( .A(n360), .B(n359), .Z(n367) );
  XOR2_X1 U418 ( .A(G155GAT), .B(KEYINPUT2), .Z(n362) );
  XNOR2_X1 U419 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n362), .B(n361), .ZN(n390) );
  XNOR2_X1 U421 ( .A(G120GAT), .B(G148GAT), .ZN(n363) );
  XNOR2_X1 U422 ( .A(n363), .B(G57GAT), .ZN(n435) );
  XNOR2_X1 U423 ( .A(n390), .B(n435), .ZN(n365) );
  XOR2_X1 U424 ( .A(n369), .B(n368), .Z(n410) );
  XNOR2_X1 U425 ( .A(KEYINPUT96), .B(n410), .ZN(n524) );
  XOR2_X1 U426 ( .A(G8GAT), .B(KEYINPUT97), .Z(n371) );
  NAND2_X1 U427 ( .A1(G226GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U428 ( .A(n371), .B(n370), .ZN(n374) );
  XOR2_X1 U429 ( .A(G64GAT), .B(G92GAT), .Z(n373) );
  XNOR2_X1 U430 ( .A(G176GAT), .B(G204GAT), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n373), .B(n372), .ZN(n443) );
  XOR2_X1 U432 ( .A(n374), .B(n443), .Z(n381) );
  XOR2_X1 U433 ( .A(KEYINPUT93), .B(G218GAT), .Z(n376) );
  XNOR2_X1 U434 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n375) );
  XNOR2_X1 U435 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U436 ( .A(G197GAT), .B(n377), .ZN(n399) );
  INV_X1 U437 ( .A(n399), .ZN(n379) );
  XNOR2_X1 U438 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U439 ( .A(n381), .B(n380), .ZN(n383) );
  XNOR2_X1 U440 ( .A(n383), .B(n382), .ZN(n527) );
  XNOR2_X1 U441 ( .A(n527), .B(KEYINPUT27), .ZN(n407) );
  NAND2_X1 U442 ( .A1(n524), .A2(n407), .ZN(n535) );
  NOR2_X1 U443 ( .A1(n538), .A2(n535), .ZN(n400) );
  XOR2_X1 U444 ( .A(KEYINPUT22), .B(KEYINPUT95), .Z(n385) );
  XNOR2_X1 U445 ( .A(G148GAT), .B(KEYINPUT23), .ZN(n384) );
  XNOR2_X1 U446 ( .A(n385), .B(n384), .ZN(n397) );
  XOR2_X1 U447 ( .A(KEYINPUT24), .B(KEYINPUT94), .Z(n388) );
  XOR2_X1 U448 ( .A(G106GAT), .B(G78GAT), .Z(n447) );
  XNOR2_X1 U449 ( .A(n386), .B(n447), .ZN(n387) );
  XNOR2_X1 U450 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U451 ( .A(n389), .B(KEYINPUT92), .Z(n395) );
  XOR2_X1 U452 ( .A(n390), .B(G204GAT), .Z(n392) );
  NAND2_X1 U453 ( .A1(G228GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U454 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U455 ( .A(G22GAT), .B(n393), .ZN(n394) );
  XNOR2_X1 U456 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U457 ( .A(n397), .B(n396), .Z(n398) );
  XNOR2_X1 U458 ( .A(n399), .B(n398), .ZN(n479) );
  XNOR2_X1 U459 ( .A(n479), .B(KEYINPUT28), .ZN(n537) );
  NAND2_X1 U460 ( .A1(n400), .A2(n537), .ZN(n401) );
  XOR2_X1 U461 ( .A(KEYINPUT98), .B(n401), .Z(n413) );
  NAND2_X1 U462 ( .A1(n527), .A2(n538), .ZN(n402) );
  NAND2_X1 U463 ( .A1(n402), .A2(n479), .ZN(n403) );
  XNOR2_X1 U464 ( .A(n403), .B(KEYINPUT100), .ZN(n404) );
  XNOR2_X1 U465 ( .A(KEYINPUT25), .B(n404), .ZN(n409) );
  NOR2_X1 U466 ( .A1(n538), .A2(n479), .ZN(n405) );
  XOR2_X1 U467 ( .A(KEYINPUT99), .B(n405), .Z(n406) );
  XNOR2_X1 U468 ( .A(KEYINPUT26), .B(n406), .ZN(n572) );
  AND2_X1 U469 ( .A1(n572), .A2(n407), .ZN(n408) );
  NOR2_X1 U470 ( .A1(n409), .A2(n408), .ZN(n411) );
  NOR2_X1 U471 ( .A1(n411), .A2(n410), .ZN(n412) );
  NOR2_X1 U472 ( .A1(n558), .A2(n492), .ZN(n414) );
  XOR2_X1 U473 ( .A(KEYINPUT106), .B(n414), .Z(n415) );
  NOR2_X1 U474 ( .A1(n586), .A2(n415), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n416), .B(KEYINPUT37), .ZN(n522) );
  XOR2_X1 U476 ( .A(G36GAT), .B(G43GAT), .Z(n418) );
  XNOR2_X1 U477 ( .A(G50GAT), .B(G29GAT), .ZN(n417) );
  XNOR2_X1 U478 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U479 ( .A(n420), .B(n419), .Z(n422) );
  NAND2_X1 U480 ( .A1(G229GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U481 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U482 ( .A(n423), .B(KEYINPUT66), .Z(n426) );
  XNOR2_X1 U483 ( .A(n424), .B(KEYINPUT29), .ZN(n425) );
  XNOR2_X1 U484 ( .A(n426), .B(n425), .ZN(n434) );
  XOR2_X1 U485 ( .A(G141GAT), .B(G197GAT), .Z(n428) );
  XNOR2_X1 U486 ( .A(G169GAT), .B(G113GAT), .ZN(n427) );
  XNOR2_X1 U487 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U488 ( .A(KEYINPUT69), .B(KEYINPUT67), .Z(n430) );
  XNOR2_X1 U489 ( .A(G1GAT), .B(KEYINPUT30), .ZN(n429) );
  XNOR2_X1 U490 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U491 ( .A(n432), .B(n431), .Z(n433) );
  XNOR2_X1 U492 ( .A(n434), .B(n433), .ZN(n574) );
  INV_X1 U493 ( .A(n574), .ZN(n552) );
  INV_X1 U494 ( .A(KEYINPUT32), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n438) );
  NAND2_X1 U496 ( .A1(G230GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U498 ( .A(KEYINPUT73), .B(KEYINPUT33), .Z(n440) );
  XNOR2_X1 U499 ( .A(KEYINPUT72), .B(KEYINPUT31), .ZN(n439) );
  XOR2_X1 U500 ( .A(n440), .B(n439), .Z(n441) );
  XNOR2_X1 U501 ( .A(n442), .B(n441), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U503 ( .A(n446), .B(n445), .ZN(n451) );
  XNOR2_X1 U504 ( .A(G99GAT), .B(G85GAT), .ZN(n449) );
  INV_X1 U505 ( .A(n447), .ZN(n448) );
  XNOR2_X1 U506 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U507 ( .A(n451), .B(n450), .ZN(n580) );
  NAND2_X1 U508 ( .A1(n552), .A2(n580), .ZN(n494) );
  NOR2_X1 U509 ( .A1(n522), .A2(n494), .ZN(n452) );
  NAND2_X1 U510 ( .A1(n538), .A2(n509), .ZN(n455) );
  XOR2_X1 U511 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n453) );
  INV_X1 U512 ( .A(n558), .ZN(n583) );
  INV_X1 U513 ( .A(KEYINPUT54), .ZN(n477) );
  INV_X1 U514 ( .A(KEYINPUT47), .ZN(n464) );
  XOR2_X1 U515 ( .A(KEYINPUT112), .B(KEYINPUT46), .Z(n458) );
  INV_X1 U516 ( .A(KEYINPUT41), .ZN(n456) );
  XNOR2_X1 U517 ( .A(n580), .B(n456), .ZN(n566) );
  INV_X1 U518 ( .A(n566), .ZN(n554) );
  NAND2_X1 U519 ( .A1(n552), .A2(n554), .ZN(n457) );
  XNOR2_X1 U520 ( .A(n458), .B(n457), .ZN(n459) );
  NOR2_X1 U521 ( .A1(n459), .A2(n558), .ZN(n460) );
  XNOR2_X1 U522 ( .A(n460), .B(KEYINPUT113), .ZN(n461) );
  NOR2_X1 U523 ( .A1(n461), .A2(n561), .ZN(n462) );
  XNOR2_X1 U524 ( .A(n462), .B(KEYINPUT114), .ZN(n463) );
  XNOR2_X1 U525 ( .A(n464), .B(n463), .ZN(n473) );
  INV_X1 U526 ( .A(n580), .ZN(n468) );
  NOR2_X1 U527 ( .A1(n586), .A2(n583), .ZN(n466) );
  XNOR2_X1 U528 ( .A(n466), .B(n465), .ZN(n467) );
  NOR2_X1 U529 ( .A1(n468), .A2(n467), .ZN(n469) );
  XNOR2_X1 U530 ( .A(n469), .B(KEYINPUT115), .ZN(n470) );
  NOR2_X1 U531 ( .A1(n470), .A2(n552), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n471), .B(KEYINPUT116), .ZN(n472) );
  NOR2_X1 U533 ( .A1(n473), .A2(n472), .ZN(n474) );
  XNOR2_X1 U534 ( .A(KEYINPUT48), .B(n474), .ZN(n534) );
  XNOR2_X1 U535 ( .A(KEYINPUT121), .B(n527), .ZN(n475) );
  NOR2_X1 U536 ( .A1(n534), .A2(n475), .ZN(n476) );
  XNOR2_X1 U537 ( .A(n477), .B(n476), .ZN(n478) );
  NAND2_X1 U538 ( .A1(n573), .A2(n479), .ZN(n480) );
  XNOR2_X1 U539 ( .A(KEYINPUT55), .B(n480), .ZN(n481) );
  NAND2_X1 U540 ( .A1(n481), .A2(n538), .ZN(n565) );
  NOR2_X1 U541 ( .A1(n583), .A2(n565), .ZN(n484) );
  INV_X1 U542 ( .A(G183GAT), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n482), .B(KEYINPUT124), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(G1350GAT) );
  NOR2_X1 U545 ( .A1(n488), .A2(n565), .ZN(n487) );
  XOR2_X1 U546 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n496) );
  NAND2_X1 U547 ( .A1(n488), .A2(n558), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n489), .B(KEYINPUT16), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n490), .B(KEYINPUT84), .ZN(n491) );
  NOR2_X1 U550 ( .A1(n492), .A2(n491), .ZN(n493) );
  XNOR2_X1 U551 ( .A(KEYINPUT101), .B(n493), .ZN(n512) );
  NOR2_X1 U552 ( .A1(n494), .A2(n512), .ZN(n503) );
  NAND2_X1 U553 ( .A1(n503), .A2(n524), .ZN(n495) );
  XNOR2_X1 U554 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U555 ( .A(G1GAT), .B(n497), .Z(G1324GAT) );
  XOR2_X1 U556 ( .A(G8GAT), .B(KEYINPUT103), .Z(n499) );
  NAND2_X1 U557 ( .A1(n503), .A2(n527), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n499), .B(n498), .ZN(G1325GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT104), .B(KEYINPUT35), .Z(n501) );
  NAND2_X1 U560 ( .A1(n503), .A2(n538), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U562 ( .A(G15GAT), .B(n502), .ZN(G1326GAT) );
  XOR2_X1 U563 ( .A(G22GAT), .B(KEYINPUT105), .Z(n505) );
  INV_X1 U564 ( .A(n537), .ZN(n530) );
  NAND2_X1 U565 ( .A1(n503), .A2(n530), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n505), .B(n504), .ZN(G1327GAT) );
  XOR2_X1 U567 ( .A(G29GAT), .B(KEYINPUT39), .Z(n507) );
  NAND2_X1 U568 ( .A1(n524), .A2(n509), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n507), .B(n506), .ZN(G1328GAT) );
  NAND2_X1 U570 ( .A1(n509), .A2(n527), .ZN(n508) );
  XNOR2_X1 U571 ( .A(n508), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U572 ( .A1(n530), .A2(n509), .ZN(n510) );
  XNOR2_X1 U573 ( .A(G50GAT), .B(n510), .ZN(G1331GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n514) );
  NAND2_X1 U575 ( .A1(n554), .A2(n574), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n511), .B(KEYINPUT108), .ZN(n523) );
  NOR2_X1 U577 ( .A1(n523), .A2(n512), .ZN(n519) );
  NAND2_X1 U578 ( .A1(n519), .A2(n524), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U580 ( .A(G57GAT), .B(n515), .ZN(G1332GAT) );
  NAND2_X1 U581 ( .A1(n527), .A2(n519), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n516), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U583 ( .A1(n519), .A2(n538), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n517), .B(KEYINPUT110), .ZN(n518) );
  XNOR2_X1 U585 ( .A(G71GAT), .B(n518), .ZN(G1334GAT) );
  XOR2_X1 U586 ( .A(G78GAT), .B(KEYINPUT43), .Z(n521) );
  NAND2_X1 U587 ( .A1(n519), .A2(n530), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(G1335GAT) );
  XOR2_X1 U589 ( .A(G85GAT), .B(KEYINPUT111), .Z(n526) );
  NOR2_X1 U590 ( .A1(n523), .A2(n522), .ZN(n531) );
  NAND2_X1 U591 ( .A1(n531), .A2(n524), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(G1336GAT) );
  NAND2_X1 U593 ( .A1(n527), .A2(n531), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n528), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U595 ( .A1(n531), .A2(n538), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n529), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U597 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n532), .B(KEYINPUT44), .ZN(n533) );
  XNOR2_X1 U599 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  NOR2_X1 U600 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n536), .B(KEYINPUT117), .ZN(n550) );
  NAND2_X1 U602 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U603 ( .A1(n550), .A2(n539), .ZN(n547) );
  NAND2_X1 U604 ( .A1(n547), .A2(n552), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n540), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT49), .B(KEYINPUT118), .Z(n542) );
  NAND2_X1 U607 ( .A1(n547), .A2(n554), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U609 ( .A(G120GAT), .B(n543), .ZN(G1341GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT119), .B(KEYINPUT50), .Z(n545) );
  NAND2_X1 U611 ( .A1(n547), .A2(n558), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  XOR2_X1 U614 ( .A(G134GAT), .B(KEYINPUT51), .Z(n549) );
  NAND2_X1 U615 ( .A1(n547), .A2(n561), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(G1343GAT) );
  INV_X1 U617 ( .A(n572), .ZN(n551) );
  NOR2_X1 U618 ( .A1(n551), .A2(n550), .ZN(n562) );
  NAND2_X1 U619 ( .A1(n552), .A2(n562), .ZN(n553) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(n553), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n556) );
  NAND2_X1 U622 ( .A1(n562), .A2(n554), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(n557), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n562), .A2(n558), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(KEYINPUT120), .ZN(n560) );
  XNOR2_X1 U627 ( .A(G155GAT), .B(n560), .ZN(G1346GAT) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U630 ( .A1(n574), .A2(n565), .ZN(n564) );
  XOR2_X1 U631 ( .A(G169GAT), .B(n564), .Z(G1348GAT) );
  NOR2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n568) );
  XNOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(KEYINPUT122), .B(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1349GAT) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n585) );
  NOR2_X1 U639 ( .A1(n574), .A2(n585), .ZN(n579) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n576) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(KEYINPUT125), .B(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n585), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NOR2_X1 U648 ( .A1(n583), .A2(n585), .ZN(n584) );
  XOR2_X1 U649 ( .A(G211GAT), .B(n584), .Z(G1354GAT) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n588) );
  XNOR2_X1 U651 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

