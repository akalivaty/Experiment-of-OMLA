

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584;

  NOR2_X1 U325 ( .A1(n464), .A2(n463), .ZN(n477) );
  NOR2_X1 U326 ( .A1(n517), .A2(n521), .ZN(n447) );
  XOR2_X1 U327 ( .A(n393), .B(n428), .Z(n510) );
  XNOR2_X1 U328 ( .A(n450), .B(KEYINPUT92), .ZN(n464) );
  XNOR2_X1 U329 ( .A(n385), .B(n293), .ZN(n386) );
  NOR2_X1 U330 ( .A1(n466), .A2(n582), .ZN(n468) );
  XNOR2_X1 U331 ( .A(n439), .B(n438), .ZN(n523) );
  XNOR2_X1 U332 ( .A(n387), .B(n386), .ZN(n388) );
  AND2_X1 U333 ( .A1(G226GAT), .A2(G233GAT), .ZN(n293) );
  XOR2_X1 U334 ( .A(KEYINPUT3), .B(G162GAT), .Z(n294) );
  AND2_X1 U335 ( .A1(G232GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U336 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n348) );
  XNOR2_X1 U337 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U338 ( .A(G190GAT), .B(KEYINPUT80), .Z(n379) );
  XNOR2_X1 U339 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n394) );
  XNOR2_X1 U340 ( .A(n316), .B(n295), .ZN(n317) );
  XNOR2_X1 U341 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U342 ( .A(n395), .B(n394), .ZN(n415) );
  XNOR2_X1 U343 ( .A(n318), .B(n317), .ZN(n322) );
  XNOR2_X1 U344 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U345 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U346 ( .A(n470), .B(KEYINPUT101), .ZN(n493) );
  XNOR2_X1 U347 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U348 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U349 ( .A(n445), .B(n444), .ZN(G1349GAT) );
  XNOR2_X1 U350 ( .A(n474), .B(n473), .ZN(G1330GAT) );
  XOR2_X1 U351 ( .A(KEYINPUT76), .B(KEYINPUT13), .Z(n297) );
  XNOR2_X1 U352 ( .A(G148GAT), .B(KEYINPUT33), .ZN(n296) );
  XNOR2_X1 U353 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U354 ( .A(KEYINPUT77), .B(KEYINPUT31), .Z(n299) );
  XNOR2_X1 U355 ( .A(KEYINPUT32), .B(KEYINPUT75), .ZN(n298) );
  XNOR2_X1 U356 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n301), .B(n300), .ZN(n311) );
  XNOR2_X1 U358 ( .A(G106GAT), .B(G78GAT), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n302), .B(G204GAT), .ZN(n416) );
  XOR2_X1 U360 ( .A(n416), .B(KEYINPUT74), .Z(n304) );
  NAND2_X1 U361 ( .A1(G230GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U362 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U363 ( .A(G92GAT), .B(G64GAT), .Z(n380) );
  XOR2_X1 U364 ( .A(G85GAT), .B(G57GAT), .Z(n396) );
  XOR2_X1 U365 ( .A(n380), .B(n396), .Z(n306) );
  XNOR2_X1 U366 ( .A(G176GAT), .B(G120GAT), .ZN(n305) );
  XNOR2_X1 U367 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U368 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U369 ( .A(G99GAT), .B(G71GAT), .ZN(n435) );
  XNOR2_X1 U370 ( .A(n309), .B(n435), .ZN(n310) );
  XNOR2_X1 U371 ( .A(n311), .B(n310), .ZN(n575) );
  XOR2_X1 U372 ( .A(n379), .B(G85GAT), .Z(n313) );
  XNOR2_X1 U373 ( .A(G43GAT), .B(G218GAT), .ZN(n312) );
  XNOR2_X1 U374 ( .A(n313), .B(n312), .ZN(n318) );
  XOR2_X1 U375 ( .A(G92GAT), .B(G162GAT), .Z(n315) );
  XNOR2_X1 U376 ( .A(G134GAT), .B(G99GAT), .ZN(n314) );
  XNOR2_X1 U377 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U378 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n320) );
  XNOR2_X1 U379 ( .A(G29GAT), .B(G106GAT), .ZN(n319) );
  XNOR2_X1 U380 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U381 ( .A(n322), .B(n321), .ZN(n330) );
  XOR2_X1 U382 ( .A(KEYINPUT7), .B(KEYINPUT71), .Z(n324) );
  XNOR2_X1 U383 ( .A(G50GAT), .B(G36GAT), .ZN(n323) );
  XNOR2_X1 U384 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U385 ( .A(KEYINPUT8), .B(n325), .Z(n358) );
  XOR2_X1 U386 ( .A(KEYINPUT9), .B(KEYINPUT79), .Z(n327) );
  XNOR2_X1 U387 ( .A(KEYINPUT66), .B(KEYINPUT78), .ZN(n326) );
  XNOR2_X1 U388 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U389 ( .A(n358), .B(n328), .ZN(n329) );
  XNOR2_X1 U390 ( .A(n330), .B(n329), .ZN(n561) );
  XOR2_X1 U391 ( .A(KEYINPUT36), .B(n561), .Z(n582) );
  XOR2_X1 U392 ( .A(G8GAT), .B(KEYINPUT72), .Z(n351) );
  XOR2_X1 U393 ( .A(G71GAT), .B(G127GAT), .Z(n332) );
  XNOR2_X1 U394 ( .A(G15GAT), .B(G183GAT), .ZN(n331) );
  XNOR2_X1 U395 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U396 ( .A(n351), .B(n333), .Z(n335) );
  NAND2_X1 U397 ( .A1(G231GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U398 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U399 ( .A(KEYINPUT15), .B(KEYINPUT81), .Z(n337) );
  XNOR2_X1 U400 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n336) );
  XNOR2_X1 U401 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U402 ( .A(n339), .B(n338), .Z(n347) );
  XOR2_X1 U403 ( .A(G78GAT), .B(G155GAT), .Z(n341) );
  XNOR2_X1 U404 ( .A(G22GAT), .B(G211GAT), .ZN(n340) );
  XNOR2_X1 U405 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U406 ( .A(KEYINPUT13), .B(G64GAT), .Z(n343) );
  XNOR2_X1 U407 ( .A(G1GAT), .B(G57GAT), .ZN(n342) );
  XNOR2_X1 U408 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U409 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U410 ( .A(n347), .B(n346), .Z(n579) );
  INV_X1 U411 ( .A(n579), .ZN(n533) );
  NOR2_X1 U412 ( .A1(n582), .A2(n533), .ZN(n349) );
  NOR2_X1 U413 ( .A1(n575), .A2(n350), .ZN(n366) );
  XOR2_X1 U414 ( .A(G29GAT), .B(G1GAT), .Z(n397) );
  XOR2_X1 U415 ( .A(n397), .B(n351), .Z(n353) );
  NAND2_X1 U416 ( .A1(G229GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U417 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U418 ( .A(G141GAT), .B(G22GAT), .Z(n417) );
  XOR2_X1 U419 ( .A(n354), .B(n417), .Z(n360) );
  XOR2_X1 U420 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n356) );
  XNOR2_X1 U421 ( .A(G197GAT), .B(KEYINPUT69), .ZN(n355) );
  XNOR2_X1 U422 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U423 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U424 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U425 ( .A(n361), .B(KEYINPUT70), .Z(n365) );
  XOR2_X1 U426 ( .A(G15GAT), .B(G113GAT), .Z(n363) );
  XNOR2_X1 U427 ( .A(G169GAT), .B(G43GAT), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n363), .B(n362), .ZN(n431) );
  XNOR2_X1 U429 ( .A(n431), .B(KEYINPUT29), .ZN(n364) );
  XOR2_X1 U430 ( .A(n365), .B(n364), .Z(n543) );
  XOR2_X1 U431 ( .A(n543), .B(KEYINPUT73), .Z(n557) );
  INV_X1 U432 ( .A(n557), .ZN(n524) );
  NAND2_X1 U433 ( .A1(n366), .A2(n524), .ZN(n373) );
  INV_X1 U434 ( .A(n561), .ZN(n536) );
  NAND2_X1 U435 ( .A1(n536), .A2(n533), .ZN(n370) );
  INV_X1 U436 ( .A(n543), .ZN(n567) );
  XNOR2_X1 U437 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n367) );
  XOR2_X1 U438 ( .A(n367), .B(n575), .Z(n547) );
  INV_X1 U439 ( .A(n547), .ZN(n527) );
  NOR2_X1 U440 ( .A1(n567), .A2(n527), .ZN(n368) );
  XNOR2_X1 U441 ( .A(n368), .B(KEYINPUT46), .ZN(n369) );
  NOR2_X1 U442 ( .A1(n370), .A2(n369), .ZN(n371) );
  XNOR2_X1 U443 ( .A(n371), .B(KEYINPUT47), .ZN(n372) );
  NAND2_X1 U444 ( .A1(n373), .A2(n372), .ZN(n374) );
  XNOR2_X1 U445 ( .A(KEYINPUT48), .B(n374), .ZN(n519) );
  XOR2_X1 U446 ( .A(G176GAT), .B(KEYINPUT83), .Z(n376) );
  XNOR2_X1 U447 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n375) );
  XNOR2_X1 U448 ( .A(n376), .B(n375), .ZN(n378) );
  XOR2_X1 U449 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n377) );
  XOR2_X1 U450 ( .A(n378), .B(n377), .Z(n437) );
  INV_X1 U451 ( .A(n437), .ZN(n389) );
  XOR2_X1 U452 ( .A(n380), .B(n379), .Z(n382) );
  XNOR2_X1 U453 ( .A(G169GAT), .B(G36GAT), .ZN(n381) );
  XNOR2_X1 U454 ( .A(n382), .B(n381), .ZN(n387) );
  XOR2_X1 U455 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n384) );
  XNOR2_X1 U456 ( .A(G8GAT), .B(G204GAT), .ZN(n383) );
  XNOR2_X1 U457 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U458 ( .A(n389), .B(n388), .Z(n393) );
  XOR2_X1 U459 ( .A(KEYINPUT85), .B(G218GAT), .Z(n391) );
  XNOR2_X1 U460 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n390) );
  XNOR2_X1 U461 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U462 ( .A(G197GAT), .B(n392), .Z(n428) );
  NAND2_X1 U463 ( .A1(n519), .A2(n510), .ZN(n395) );
  XOR2_X1 U464 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n399) );
  XNOR2_X1 U465 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U466 ( .A(n399), .B(n398), .ZN(n402) );
  XNOR2_X1 U467 ( .A(G155GAT), .B(G148GAT), .ZN(n400) );
  XNOR2_X1 U468 ( .A(n294), .B(n400), .ZN(n401) );
  XOR2_X1 U469 ( .A(KEYINPUT2), .B(n401), .Z(n424) );
  XNOR2_X1 U470 ( .A(n402), .B(n424), .ZN(n403) );
  INV_X1 U471 ( .A(n403), .ZN(n405) );
  XNOR2_X1 U472 ( .A(G113GAT), .B(G141GAT), .ZN(n404) );
  XNOR2_X1 U473 ( .A(n405), .B(n404), .ZN(n409) );
  XOR2_X1 U474 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n407) );
  NAND2_X1 U475 ( .A1(G225GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U476 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U477 ( .A(n409), .B(n408), .Z(n414) );
  XOR2_X1 U478 ( .A(KEYINPUT0), .B(G134GAT), .Z(n411) );
  XNOR2_X1 U479 ( .A(G127GAT), .B(G120GAT), .ZN(n410) );
  XNOR2_X1 U480 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U481 ( .A(KEYINPUT82), .B(n412), .Z(n433) );
  XNOR2_X1 U482 ( .A(n433), .B(KEYINPUT87), .ZN(n413) );
  XNOR2_X1 U483 ( .A(n414), .B(n413), .ZN(n460) );
  XOR2_X2 U484 ( .A(KEYINPUT88), .B(n460), .Z(n508) );
  NOR2_X1 U485 ( .A1(n415), .A2(n508), .ZN(n566) );
  XOR2_X1 U486 ( .A(KEYINPUT24), .B(n416), .Z(n419) );
  XNOR2_X1 U487 ( .A(G50GAT), .B(n417), .ZN(n418) );
  XNOR2_X1 U488 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U489 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n421) );
  NAND2_X1 U490 ( .A1(G228GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U491 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U492 ( .A(n423), .B(n422), .Z(n426) );
  XNOR2_X1 U493 ( .A(n424), .B(KEYINPUT86), .ZN(n425) );
  XNOR2_X1 U494 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U495 ( .A(n428), .B(n427), .ZN(n454) );
  NAND2_X1 U496 ( .A1(n566), .A2(n454), .ZN(n429) );
  XNOR2_X1 U497 ( .A(KEYINPUT55), .B(n429), .ZN(n440) );
  XOR2_X1 U498 ( .A(KEYINPUT20), .B(G190GAT), .Z(n430) );
  XNOR2_X1 U499 ( .A(n435), .B(n434), .ZN(n439) );
  AND2_X1 U500 ( .A1(G227GAT), .A2(G233GAT), .ZN(n436) );
  NAND2_X1 U501 ( .A1(n440), .A2(n523), .ZN(n441) );
  XNOR2_X1 U502 ( .A(KEYINPUT121), .B(n441), .ZN(n562) );
  NAND2_X1 U503 ( .A1(n562), .A2(n547), .ZN(n445) );
  XOR2_X1 U504 ( .A(G176GAT), .B(KEYINPUT56), .Z(n443) );
  XOR2_X1 U505 ( .A(KEYINPUT123), .B(KEYINPUT57), .Z(n442) );
  XNOR2_X1 U506 ( .A(n523), .B(KEYINPUT84), .ZN(n449) );
  XNOR2_X1 U507 ( .A(KEYINPUT27), .B(n510), .ZN(n457) );
  NAND2_X1 U508 ( .A1(n508), .A2(n457), .ZN(n517) );
  XNOR2_X1 U509 ( .A(KEYINPUT67), .B(KEYINPUT28), .ZN(n446) );
  XNOR2_X1 U510 ( .A(n446), .B(n454), .ZN(n521) );
  XNOR2_X1 U511 ( .A(n447), .B(KEYINPUT91), .ZN(n448) );
  NOR2_X1 U512 ( .A1(n449), .A2(n448), .ZN(n450) );
  NAND2_X1 U513 ( .A1(n510), .A2(n523), .ZN(n451) );
  NAND2_X1 U514 ( .A1(n451), .A2(n454), .ZN(n452) );
  XNOR2_X1 U515 ( .A(n452), .B(KEYINPUT93), .ZN(n453) );
  XNOR2_X1 U516 ( .A(KEYINPUT25), .B(n453), .ZN(n459) );
  NOR2_X1 U517 ( .A1(n454), .A2(n523), .ZN(n455) );
  XOR2_X1 U518 ( .A(n455), .B(KEYINPUT26), .Z(n565) );
  INV_X1 U519 ( .A(n565), .ZN(n456) );
  NAND2_X1 U520 ( .A1(n457), .A2(n456), .ZN(n458) );
  NAND2_X1 U521 ( .A1(n459), .A2(n458), .ZN(n461) );
  NAND2_X1 U522 ( .A1(n461), .A2(n460), .ZN(n462) );
  XOR2_X1 U523 ( .A(KEYINPUT94), .B(n462), .Z(n463) );
  NOR2_X1 U524 ( .A1(n477), .A2(n579), .ZN(n465) );
  XNOR2_X1 U525 ( .A(n465), .B(KEYINPUT99), .ZN(n466) );
  XOR2_X1 U526 ( .A(KEYINPUT37), .B(KEYINPUT100), .Z(n467) );
  XNOR2_X1 U527 ( .A(n468), .B(n467), .ZN(n506) );
  NOR2_X1 U528 ( .A1(n524), .A2(n575), .ZN(n478) );
  NAND2_X1 U529 ( .A1(n506), .A2(n478), .ZN(n469) );
  XNOR2_X1 U530 ( .A(n469), .B(KEYINPUT38), .ZN(n470) );
  NAND2_X1 U531 ( .A1(n523), .A2(n493), .ZN(n474) );
  XOR2_X1 U532 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n472) );
  XNOR2_X1 U533 ( .A(G43GAT), .B(KEYINPUT102), .ZN(n471) );
  NOR2_X1 U534 ( .A1(n533), .A2(n561), .ZN(n475) );
  XOR2_X1 U535 ( .A(KEYINPUT16), .B(n475), .Z(n476) );
  NOR2_X1 U536 ( .A1(n477), .A2(n476), .ZN(n496) );
  AND2_X1 U537 ( .A1(n478), .A2(n496), .ZN(n487) );
  NAND2_X1 U538 ( .A1(n487), .A2(n508), .ZN(n482) );
  XOR2_X1 U539 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n480) );
  XNOR2_X1 U540 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n479) );
  XNOR2_X1 U541 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n482), .B(n481), .ZN(G1324GAT) );
  XOR2_X1 U543 ( .A(G8GAT), .B(KEYINPUT97), .Z(n484) );
  NAND2_X1 U544 ( .A1(n487), .A2(n510), .ZN(n483) );
  XNOR2_X1 U545 ( .A(n484), .B(n483), .ZN(G1325GAT) );
  XOR2_X1 U546 ( .A(G15GAT), .B(KEYINPUT35), .Z(n486) );
  NAND2_X1 U547 ( .A1(n487), .A2(n523), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n486), .B(n485), .ZN(G1326GAT) );
  NAND2_X1 U549 ( .A1(n521), .A2(n487), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n488), .B(KEYINPUT98), .ZN(n489) );
  XNOR2_X1 U551 ( .A(G22GAT), .B(n489), .ZN(G1327GAT) );
  NAND2_X1 U552 ( .A1(n508), .A2(n493), .ZN(n491) );
  XOR2_X1 U553 ( .A(G29GAT), .B(KEYINPUT39), .Z(n490) );
  XNOR2_X1 U554 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  NAND2_X1 U555 ( .A1(n493), .A2(n510), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n492), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U557 ( .A1(n493), .A2(n521), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n494), .B(KEYINPUT104), .ZN(n495) );
  XNOR2_X1 U559 ( .A(G50GAT), .B(n495), .ZN(G1331GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT42), .B(KEYINPUT105), .Z(n498) );
  NOR2_X1 U561 ( .A1(n543), .A2(n527), .ZN(n505) );
  AND2_X1 U562 ( .A1(n505), .A2(n496), .ZN(n502) );
  NAND2_X1 U563 ( .A1(n502), .A2(n508), .ZN(n497) );
  XNOR2_X1 U564 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(n499), .ZN(G1332GAT) );
  NAND2_X1 U566 ( .A1(n510), .A2(n502), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n500), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U568 ( .A1(n502), .A2(n523), .ZN(n501) );
  XNOR2_X1 U569 ( .A(n501), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U570 ( .A(G78GAT), .B(KEYINPUT43), .Z(n504) );
  NAND2_X1 U571 ( .A1(n502), .A2(n521), .ZN(n503) );
  XNOR2_X1 U572 ( .A(n504), .B(n503), .ZN(G1335GAT) );
  NAND2_X1 U573 ( .A1(n506), .A2(n505), .ZN(n507) );
  XOR2_X1 U574 ( .A(KEYINPUT106), .B(n507), .Z(n513) );
  NAND2_X1 U575 ( .A1(n508), .A2(n513), .ZN(n509) );
  XNOR2_X1 U576 ( .A(G85GAT), .B(n509), .ZN(G1336GAT) );
  NAND2_X1 U577 ( .A1(n513), .A2(n510), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n511), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U579 ( .A1(n513), .A2(n523), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n512), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT44), .B(KEYINPUT107), .Z(n515) );
  NAND2_X1 U582 ( .A1(n513), .A2(n521), .ZN(n514) );
  XNOR2_X1 U583 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U584 ( .A(G106GAT), .B(n516), .ZN(G1339GAT) );
  INV_X1 U585 ( .A(n517), .ZN(n518) );
  NAND2_X1 U586 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U587 ( .A(KEYINPUT108), .B(n520), .ZN(n542) );
  NOR2_X1 U588 ( .A1(n542), .A2(n521), .ZN(n522) );
  NAND2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n537) );
  NOR2_X1 U590 ( .A1(n524), .A2(n537), .ZN(n526) );
  XNOR2_X1 U591 ( .A(G113GAT), .B(KEYINPUT109), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(G1340GAT) );
  NOR2_X1 U593 ( .A1(n527), .A2(n537), .ZN(n529) );
  XNOR2_X1 U594 ( .A(KEYINPUT110), .B(KEYINPUT49), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U596 ( .A(G120GAT), .B(n530), .ZN(G1341GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n532) );
  XNOR2_X1 U598 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(n535) );
  NOR2_X1 U600 ( .A1(n533), .A2(n537), .ZN(n534) );
  XOR2_X1 U601 ( .A(n535), .B(n534), .Z(G1342GAT) );
  NOR2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n541) );
  XOR2_X1 U603 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n539) );
  XNOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT114), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(G1343GAT) );
  NOR2_X1 U607 ( .A1(n565), .A2(n542), .ZN(n554) );
  NAND2_X1 U608 ( .A1(n554), .A2(n543), .ZN(n544) );
  XNOR2_X1 U609 ( .A(G141GAT), .B(n544), .ZN(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT117), .B(KEYINPUT116), .Z(n546) );
  XNOR2_X1 U611 ( .A(KEYINPUT115), .B(KEYINPUT53), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n551) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n549) );
  NAND2_X1 U614 ( .A1(n547), .A2(n554), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(G1345GAT) );
  NAND2_X1 U617 ( .A1(n579), .A2(n554), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n552), .B(KEYINPUT118), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G155GAT), .B(n553), .ZN(G1346GAT) );
  XOR2_X1 U620 ( .A(G162GAT), .B(KEYINPUT119), .Z(n556) );
  NAND2_X1 U621 ( .A1(n554), .A2(n561), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1347GAT) );
  XNOR2_X1 U623 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n559) );
  NAND2_X1 U624 ( .A1(n562), .A2(n557), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1348GAT) );
  NAND2_X1 U626 ( .A1(n579), .A2(n562), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U628 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n564) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1351GAT) );
  NAND2_X1 U631 ( .A1(n566), .A2(n456), .ZN(n581) );
  NOR2_X1 U632 ( .A1(n581), .A2(n567), .ZN(n574) );
  XOR2_X1 U633 ( .A(KEYINPUT124), .B(KEYINPUT126), .Z(n569) );
  XNOR2_X1 U634 ( .A(KEYINPUT59), .B(KEYINPUT60), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XOR2_X1 U636 ( .A(n570), .B(KEYINPUT127), .Z(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  INV_X1 U641 ( .A(n581), .ZN(n578) );
  NAND2_X1 U642 ( .A1(n578), .A2(n575), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U647 ( .A(KEYINPUT62), .B(n583), .Z(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

