//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 0 0 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(G469), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT83), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT65), .B1(new_n193), .B2(G143), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(new_n191), .A3(G146), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n192), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n193), .A2(G143), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(KEYINPUT1), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n190), .B1(new_n197), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n194), .A2(new_n196), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(new_n199), .ZN(new_n203));
  INV_X1    g017(.A(new_n200), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(KEYINPUT83), .A3(new_n204), .ZN(new_n205));
  AND3_X1   g019(.A1(new_n197), .A2(KEYINPUT82), .A3(new_n200), .ZN(new_n206));
  AOI21_X1  g020(.A(KEYINPUT82), .B1(new_n197), .B2(new_n200), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n201), .B(new_n205), .C1(new_n206), .C2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT80), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(KEYINPUT3), .ZN(new_n210));
  INV_X1    g024(.A(G104), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G107), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(KEYINPUT3), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n210), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(G107), .ZN(new_n215));
  INV_X1    g029(.A(G107), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G104), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT80), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n215), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G101), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n216), .A2(G104), .ZN(new_n223));
  OAI21_X1  g037(.A(G101), .B1(new_n212), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT81), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT81), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n226), .B(G101), .C1(new_n212), .C2(new_n223), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n221), .A2(new_n222), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(KEYINPUT10), .B1(new_n208), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(G101), .B1(new_n214), .B2(new_n220), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n223), .B1(new_n212), .B2(new_n210), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n218), .A2(KEYINPUT80), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n219), .B1(new_n233), .B2(new_n217), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n232), .A2(new_n222), .A3(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n231), .A2(KEYINPUT4), .A3(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT64), .B1(new_n193), .B2(G143), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT64), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(new_n191), .A3(G146), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(new_n199), .ZN(new_n241));
  NAND2_X1  g055(.A1(KEYINPUT0), .A2(G128), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(KEYINPUT0), .A2(G128), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n241), .A2(new_n245), .B1(new_n197), .B2(new_n243), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n247), .B(G101), .C1(new_n214), .C2(new_n220), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n236), .A2(new_n246), .A3(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n202), .A2(new_n200), .A3(new_n199), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n192), .B1(new_n237), .B2(new_n239), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n250), .B1(new_n251), .B2(new_n200), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n225), .A2(new_n227), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n252), .A2(new_n253), .A3(KEYINPUT10), .A4(new_n235), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G137), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT11), .B1(new_n257), .B2(G134), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(G134), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT66), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n257), .ZN(new_n262));
  NAND2_X1  g076(.A1(KEYINPUT66), .A2(G137), .ZN(new_n263));
  AND2_X1   g077(.A1(KEYINPUT11), .A2(G134), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G131), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n260), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n266), .B1(new_n260), .B2(new_n265), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n230), .A2(new_n256), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n260), .A2(new_n265), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G131), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n260), .A2(new_n265), .A3(new_n266), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n274), .B1(new_n229), .B2(new_n255), .ZN(new_n275));
  XNOR2_X1  g089(.A(G110), .B(G140), .ZN(new_n276));
  INV_X1    g090(.A(G227), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n277), .A2(G953), .ZN(new_n278));
  XOR2_X1   g092(.A(new_n276), .B(new_n278), .Z(new_n279));
  NAND3_X1  g093(.A1(new_n270), .A2(new_n275), .A3(new_n279), .ZN(new_n280));
  NOR3_X1   g094(.A1(new_n229), .A2(new_n255), .A3(new_n274), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n253), .A2(new_n235), .ZN(new_n282));
  AOI21_X1  g096(.A(KEYINPUT83), .B1(new_n203), .B2(new_n204), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n197), .A2(new_n190), .A3(new_n200), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT82), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n250), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n197), .A2(KEYINPUT82), .A3(new_n200), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n282), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n228), .A2(new_n252), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n274), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT12), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n208), .A2(new_n228), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n251), .A2(new_n200), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n282), .A2(new_n297), .A3(new_n250), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n269), .B1(new_n295), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT12), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n281), .B1(new_n294), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n280), .B1(new_n301), .B2(new_n279), .ZN(new_n302));
  INV_X1    g116(.A(G902), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n189), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  XOR2_X1   g118(.A(KEYINPUT71), .B(G902), .Z(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n299), .A2(KEYINPUT12), .ZN(new_n307));
  AOI211_X1 g121(.A(new_n293), .B(new_n269), .C1(new_n295), .C2(new_n298), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n270), .B(new_n279), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n279), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n269), .B1(new_n230), .B2(new_n256), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n310), .B1(new_n311), .B2(new_n281), .ZN(new_n312));
  AOI211_X1 g126(.A(G469), .B(new_n306), .C1(new_n309), .C2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n188), .B1(new_n304), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT84), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G116), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G122), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(G122), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n318), .B1(new_n319), .B2(KEYINPUT14), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT95), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI211_X1 g136(.A(KEYINPUT95), .B(new_n318), .C1(new_n319), .C2(KEYINPUT14), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n322), .B(new_n323), .C1(KEYINPUT14), .C2(new_n318), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G107), .ZN(new_n325));
  INV_X1    g139(.A(new_n319), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT93), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n318), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G122), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n329), .A2(G116), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT93), .B1(new_n319), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(G107), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT94), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n327), .B1(new_n326), .B2(new_n318), .ZN(new_n335));
  NOR3_X1   g149(.A1(new_n319), .A2(new_n330), .A3(KEYINPUT93), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n216), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT94), .ZN(new_n338));
  XNOR2_X1  g152(.A(G128), .B(G143), .ZN(new_n339));
  INV_X1    g153(.A(G134), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n339), .B(new_n340), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n325), .A2(new_n334), .A3(new_n338), .A4(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT13), .B1(new_n198), .B2(G143), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n343), .A2(new_n340), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(new_n339), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n335), .A2(new_n336), .A3(new_n216), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n345), .B1(new_n346), .B2(new_n332), .ZN(new_n347));
  INV_X1    g161(.A(G217), .ZN(new_n348));
  NOR3_X1   g162(.A1(new_n187), .A2(new_n348), .A3(G953), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n342), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n349), .B1(new_n342), .B2(new_n347), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n305), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G478), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n354), .A2(KEYINPUT15), .ZN(new_n355));
  OR3_X1    g169(.A1(new_n353), .A2(KEYINPUT97), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT97), .B1(new_n353), .B2(new_n355), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n342), .A2(new_n347), .ZN(new_n358));
  INV_X1    g172(.A(new_n349), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n306), .B1(new_n360), .B2(new_n350), .ZN(new_n361));
  INV_X1    g175(.A(new_n355), .ZN(new_n362));
  NOR3_X1   g176(.A1(new_n361), .A2(KEYINPUT96), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT96), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(new_n353), .B2(new_n355), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n356), .B(new_n357), .C1(new_n363), .C2(new_n365), .ZN(new_n366));
  OR2_X1    g180(.A1(KEYINPUT69), .A2(G237), .ZN(new_n367));
  NAND2_X1  g181(.A1(KEYINPUT69), .A2(G237), .ZN(new_n368));
  AOI21_X1  g182(.A(G953), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(G143), .A3(G214), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(G143), .B1(new_n369), .B2(G214), .ZN(new_n372));
  OAI21_X1  g186(.A(G131), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n372), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(new_n266), .A3(new_n370), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT17), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n373), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G140), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(KEYINPUT75), .A3(G125), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(G125), .ZN(new_n380));
  INV_X1    g194(.A(G125), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G140), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  OAI211_X1 g197(.A(KEYINPUT16), .B(new_n379), .C1(new_n383), .C2(KEYINPUT75), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT16), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G146), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n384), .A2(new_n193), .A3(new_n386), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n377), .B(new_n391), .C1(new_n376), .C2(new_n373), .ZN(new_n392));
  XNOR2_X1  g206(.A(G113), .B(G122), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(new_n211), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT18), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n374), .B(new_n370), .C1(new_n395), .C2(new_n266), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n383), .A2(G146), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n379), .B1(new_n383), .B2(KEYINPUT75), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n398), .B1(new_n399), .B2(new_n193), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n396), .B(new_n400), .C1(new_n373), .C2(new_n395), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n392), .A2(new_n394), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n394), .B1(new_n392), .B2(new_n401), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n303), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G475), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n373), .A2(new_n375), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT19), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n380), .A2(new_n382), .A3(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n409), .B1(new_n399), .B2(new_n408), .ZN(new_n410));
  OR2_X1    g224(.A1(new_n410), .A2(G146), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n407), .A2(new_n388), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n394), .B1(new_n412), .B2(new_n401), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n266), .B1(new_n374), .B2(new_n370), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n390), .B1(KEYINPUT17), .B2(new_n414), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n396), .A2(new_n400), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(KEYINPUT18), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n415), .A2(new_n377), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n413), .B1(new_n418), .B2(new_n394), .ZN(new_n419));
  NOR2_X1   g233(.A1(G475), .A2(G902), .ZN(new_n420));
  XOR2_X1   g234(.A(new_n420), .B(KEYINPUT92), .Z(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n419), .A2(KEYINPUT20), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT20), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n412), .A2(new_n401), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n402), .B1(new_n425), .B2(new_n394), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n424), .B1(new_n426), .B2(new_n421), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n406), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(G234), .A2(G237), .ZN(new_n429));
  INV_X1    g243(.A(G953), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n429), .A2(G952), .A3(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(G898), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(KEYINPUT98), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n306), .A2(G953), .A3(new_n429), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n431), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NOR3_X1   g250(.A1(new_n366), .A2(new_n428), .A3(new_n436), .ZN(new_n437));
  OAI211_X1 g251(.A(KEYINPUT84), .B(new_n188), .C1(new_n304), .C2(new_n313), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n316), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(G214), .B1(G237), .B2(G902), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT86), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n441), .B1(new_n252), .B2(G125), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n297), .A2(KEYINPUT86), .A3(new_n381), .A4(new_n250), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n246), .A2(new_n381), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G224), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(G953), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT7), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n447), .A2(KEYINPUT89), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT89), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n445), .B1(new_n442), .B2(new_n443), .ZN(new_n454));
  INV_X1    g268(.A(new_n451), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(G110), .B(G122), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n458), .B(KEYINPUT8), .ZN(new_n459));
  XNOR2_X1  g273(.A(G116), .B(G119), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT5), .ZN(new_n461));
  INV_X1    g275(.A(G113), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n317), .A2(G119), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT5), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n466), .A2(KEYINPUT88), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n466), .A2(KEYINPUT88), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n461), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT68), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT2), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n471), .A3(new_n462), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n472), .A2(new_n473), .B1(KEYINPUT2), .B2(G113), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n460), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n469), .A2(new_n475), .A3(new_n228), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n461), .A2(new_n465), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n228), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n459), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n454), .A2(new_n455), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n474), .B(new_n460), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n236), .A2(new_n481), .A3(new_n248), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n253), .A2(new_n475), .A3(new_n235), .A4(new_n477), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n483), .A3(new_n458), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n479), .A2(new_n480), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n303), .B1(new_n457), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n482), .A2(new_n483), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT85), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT85), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n482), .A2(new_n483), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n458), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n484), .ZN(new_n492));
  OAI21_X1  g306(.A(KEYINPUT6), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n458), .ZN(new_n494));
  INV_X1    g308(.A(new_n490), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n489), .B1(new_n482), .B2(new_n483), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT6), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n493), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n454), .A2(KEYINPUT87), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT87), .ZN(new_n502));
  AOI211_X1 g316(.A(new_n502), .B(new_n445), .C1(new_n442), .C2(new_n443), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n449), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n447), .A2(new_n502), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n454), .A2(KEYINPUT87), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n450), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n486), .B1(new_n500), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(G210), .B1(G237), .B2(G902), .ZN(new_n511));
  OAI21_X1  g325(.A(KEYINPUT90), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n498), .B1(new_n497), .B2(new_n484), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n491), .A2(KEYINPUT6), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n504), .B(new_n507), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n485), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n452), .A2(new_n456), .ZN(new_n517));
  AOI21_X1  g331(.A(G902), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n515), .A2(new_n511), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT91), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT90), .ZN(new_n521));
  INV_X1    g335(.A(new_n511), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n508), .B1(new_n493), .B2(new_n499), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n521), .B(new_n522), .C1(new_n523), .C2(new_n486), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT91), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n515), .A2(new_n525), .A3(new_n511), .A4(new_n518), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n512), .A2(new_n520), .A3(new_n524), .A4(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n439), .A2(KEYINPUT99), .A3(new_n440), .A4(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(G472), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n369), .A2(G210), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT27), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT27), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n369), .A2(new_n532), .A3(G210), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  XOR2_X1   g348(.A(KEYINPUT26), .B(G101), .Z(new_n535));
  NOR2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n534), .A2(new_n535), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n481), .ZN(new_n540));
  INV_X1    g354(.A(new_n245), .ZN(new_n541));
  OAI22_X1  g355(.A1(new_n203), .A2(new_n242), .B1(new_n541), .B2(new_n251), .ZN(new_n542));
  OAI21_X1  g356(.A(KEYINPUT67), .B1(new_n269), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT67), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n274), .A2(new_n544), .A3(new_n246), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT30), .ZN(new_n546));
  INV_X1    g360(.A(new_n263), .ZN(new_n547));
  NOR2_X1   g361(.A1(KEYINPUT66), .A2(G137), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n340), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n259), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(G131), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n197), .A2(new_n200), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n273), .B(new_n551), .C1(new_n552), .C2(new_n296), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n543), .A2(new_n545), .A3(new_n546), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n241), .A2(new_n245), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n197), .A2(new_n243), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n555), .B(new_n556), .C1(new_n267), .C2(new_n268), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT30), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n540), .B1(new_n554), .B2(new_n559), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n540), .A2(new_n553), .A3(new_n557), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n539), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT29), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n561), .A2(KEYINPUT28), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n543), .A2(new_n553), .A3(new_n545), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n561), .B1(new_n566), .B2(new_n481), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT28), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n565), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT70), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n537), .A2(new_n538), .A3(new_n570), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n534), .A2(new_n535), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT70), .B1(new_n572), .B2(new_n536), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n562), .B(new_n563), .C1(new_n569), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n558), .A2(new_n481), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n540), .A2(new_n553), .A3(new_n557), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n568), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(new_n564), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n539), .A2(new_n563), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n306), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n529), .B1(new_n575), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n554), .A2(new_n559), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n481), .ZN(new_n585));
  INV_X1    g399(.A(new_n539), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n577), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT31), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n569), .A2(new_n574), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n560), .A2(new_n561), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT31), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n591), .A3(new_n586), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n588), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT32), .ZN(new_n594));
  NOR2_X1   g408(.A1(G472), .A2(G902), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n594), .B1(new_n593), .B2(new_n595), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n583), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT72), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n348), .B1(new_n305), .B2(G234), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(G110), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT73), .ZN(new_n603));
  INV_X1    g417(.A(G119), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(G128), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(KEYINPUT23), .B1(new_n198), .B2(G119), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n603), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n198), .B(G119), .C1(KEYINPUT73), .C2(KEYINPUT23), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n602), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT74), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n198), .A2(G119), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n605), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT24), .B(G110), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  AOI22_X1  g430(.A1(new_n610), .A2(new_n611), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n390), .B(new_n617), .C1(new_n611), .C2(new_n610), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n397), .B1(new_n387), .B2(G146), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT76), .B1(new_n614), .B2(new_n616), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n608), .A2(new_n602), .A3(new_n609), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT76), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n613), .A2(new_n615), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n620), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT77), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(KEYINPUT77), .B1(new_n619), .B2(new_n624), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n618), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(KEYINPUT78), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT22), .B(G137), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n430), .A2(G221), .A3(G234), .ZN(new_n632));
  XOR2_X1   g446(.A(new_n631), .B(new_n632), .Z(new_n633));
  INV_X1    g447(.A(KEYINPUT78), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n618), .B(new_n634), .C1(new_n627), .C2(new_n628), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n630), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  OR2_X1    g450(.A1(new_n627), .A2(new_n628), .ZN(new_n637));
  INV_X1    g451(.A(new_n633), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n637), .A2(new_n634), .A3(new_n638), .A4(new_n618), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n306), .B1(new_n636), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT25), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n601), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n642), .B1(new_n641), .B2(new_n640), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n636), .A2(new_n639), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n644), .A2(KEYINPUT79), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n600), .A2(G902), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n644), .A2(KEYINPUT79), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n643), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n591), .B1(new_n590), .B2(new_n586), .ZN(new_n650));
  INV_X1    g464(.A(new_n574), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n266), .B1(new_n549), .B2(new_n259), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n267), .A2(new_n652), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n557), .A2(KEYINPUT67), .B1(new_n252), .B2(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n540), .B1(new_n654), .B2(new_n545), .ZN(new_n655));
  OAI21_X1  g469(.A(KEYINPUT28), .B1(new_n655), .B2(new_n561), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n651), .B1(new_n656), .B2(new_n565), .ZN(new_n657));
  NOR4_X1   g471(.A1(new_n560), .A2(KEYINPUT31), .A3(new_n561), .A4(new_n539), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n650), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n595), .ZN(new_n660));
  OAI21_X1  g474(.A(KEYINPUT32), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT72), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n663), .A2(new_n664), .A3(new_n583), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n599), .A2(new_n649), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT99), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n527), .A2(new_n440), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n316), .A2(new_n437), .A3(new_n438), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n528), .A2(new_n666), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT100), .B(G101), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G3));
  NAND2_X1  g487(.A1(new_n593), .A2(new_n305), .ZN(new_n674));
  OR2_X1    g488(.A1(new_n674), .A2(KEYINPUT101), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(KEYINPUT101), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n529), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n659), .A2(new_n660), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n316), .A2(new_n438), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n643), .A2(new_n648), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n440), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n522), .B1(new_n523), .B2(new_n486), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n684), .B1(new_n685), .B2(new_n519), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n361), .A2(new_n354), .ZN(new_n687));
  OAI21_X1  g501(.A(KEYINPUT33), .B1(new_n351), .B2(new_n352), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT33), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n360), .A2(new_n689), .A3(new_n350), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n306), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n687), .B1(new_n691), .B2(new_n354), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n428), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n694), .A2(new_n436), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n683), .A2(new_n686), .A3(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(new_n696), .B(KEYINPUT102), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT103), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT34), .B(G104), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G6));
  OAI21_X1  g514(.A(KEYINPUT20), .B1(new_n419), .B2(new_n422), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n426), .A2(new_n424), .A3(new_n421), .ZN(new_n702));
  AOI22_X1  g516(.A1(new_n701), .A2(new_n702), .B1(new_n405), .B2(G475), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n366), .A2(new_n703), .ZN(new_n704));
  OR3_X1    g518(.A1(new_n704), .A2(KEYINPUT104), .A3(new_n436), .ZN(new_n705));
  OAI21_X1  g519(.A(KEYINPUT104), .B1(new_n704), .B2(new_n436), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n683), .A2(new_n686), .A3(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT35), .B(G107), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G9));
  NOR2_X1   g524(.A1(new_n638), .A2(KEYINPUT36), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT105), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n629), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n646), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n644), .A2(new_n641), .A3(new_n305), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n600), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n640), .A2(new_n641), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n714), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n677), .A2(new_n719), .A3(new_n678), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n528), .A2(new_n670), .A3(new_n720), .ZN(new_n721));
  XOR2_X1   g535(.A(KEYINPUT37), .B(G110), .Z(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G12));
  AND3_X1   g537(.A1(new_n316), .A2(new_n438), .A3(new_n686), .ZN(new_n724));
  INV_X1    g538(.A(G900), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n431), .B1(new_n435), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n704), .A2(new_n726), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n727), .A2(new_n718), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n724), .A2(new_n728), .A3(new_n599), .A4(new_n665), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G128), .ZN(G30));
  XNOR2_X1  g544(.A(new_n527), .B(KEYINPUT106), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT38), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(new_n733));
  XOR2_X1   g547(.A(new_n726), .B(KEYINPUT39), .Z(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n680), .A2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(KEYINPUT40), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n737), .A2(KEYINPUT40), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n576), .A2(new_n577), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n574), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n587), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n529), .B1(new_n742), .B2(new_n303), .ZN(new_n743));
  XOR2_X1   g557(.A(new_n743), .B(KEYINPUT107), .Z(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n663), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n363), .A2(new_n365), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n356), .A2(new_n357), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n703), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n745), .A2(new_n440), .A3(new_n719), .A4(new_n748), .ZN(new_n749));
  OR4_X1    g563(.A1(new_n733), .A2(new_n738), .A3(new_n739), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G143), .ZN(G45));
  NOR3_X1   g565(.A1(new_n703), .A2(new_n692), .A3(new_n726), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n718), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n724), .A2(new_n599), .A3(new_n665), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G146), .ZN(G48));
  AOI21_X1  g569(.A(new_n664), .B1(new_n663), .B2(new_n583), .ZN(new_n756));
  AOI211_X1 g570(.A(KEYINPUT72), .B(new_n582), .C1(new_n661), .C2(new_n662), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n309), .A2(new_n312), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n305), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(G469), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT108), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n759), .A2(new_n189), .A3(new_n305), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n760), .A2(KEYINPUT108), .A3(G469), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n188), .A3(new_n686), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n758), .A2(new_n649), .A3(new_n768), .A4(new_n695), .ZN(new_n769));
  XNOR2_X1  g583(.A(KEYINPUT41), .B(G113), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(G15));
  NAND4_X1  g585(.A1(new_n758), .A2(new_n707), .A3(new_n768), .A4(new_n649), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G116), .ZN(G18));
  AND2_X1   g587(.A1(new_n437), .A2(new_n718), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n758), .A2(new_n768), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G119), .ZN(G21));
  NAND2_X1  g590(.A1(new_n766), .A2(new_n188), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n574), .B1(new_n578), .B2(new_n564), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n588), .A2(new_n779), .A3(KEYINPUT109), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n592), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT109), .B1(new_n588), .B2(new_n779), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n595), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n674), .A2(G472), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n681), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n436), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n686), .A2(new_n748), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n778), .A2(new_n786), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G122), .ZN(G24));
  NAND4_X1  g604(.A1(new_n718), .A2(new_n752), .A3(new_n784), .A4(new_n783), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n767), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(KEYINPUT110), .B(G125), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n792), .B(new_n793), .ZN(G27));
  NOR3_X1   g608(.A1(new_n527), .A2(new_n684), .A3(new_n314), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n681), .B1(new_n583), .B2(new_n663), .ZN(new_n796));
  INV_X1    g610(.A(new_n752), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT42), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n795), .A2(new_n796), .A3(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n666), .A2(KEYINPUT111), .A3(new_n752), .A4(new_n795), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n798), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n599), .A2(new_n649), .A3(new_n665), .ZN(new_n803));
  INV_X1    g617(.A(new_n524), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n515), .A2(new_n518), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n521), .B1(new_n805), .B2(new_n522), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n520), .A2(new_n526), .ZN(new_n808));
  INV_X1    g622(.A(new_n314), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n807), .A2(new_n808), .A3(new_n440), .A4(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n803), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT111), .B1(new_n811), .B2(new_n752), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n800), .B1(new_n802), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G131), .ZN(G33));
  NAND3_X1  g628(.A1(new_n666), .A2(new_n727), .A3(new_n795), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G134), .ZN(G36));
  XNOR2_X1  g630(.A(new_n302), .B(KEYINPUT45), .ZN(new_n817));
  OAI21_X1  g631(.A(G469), .B1(new_n817), .B2(G902), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n818), .A2(KEYINPUT46), .ZN(new_n819));
  OR3_X1    g633(.A1(new_n819), .A2(KEYINPUT112), .A3(new_n313), .ZN(new_n820));
  OAI21_X1  g634(.A(KEYINPUT112), .B1(new_n819), .B2(new_n313), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n820), .B(new_n821), .C1(KEYINPUT46), .C2(new_n818), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n822), .A2(new_n188), .A3(new_n734), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n693), .A2(new_n703), .ZN(new_n824));
  XOR2_X1   g638(.A(new_n824), .B(KEYINPUT43), .Z(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n718), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT44), .ZN(new_n827));
  OR3_X1    g641(.A1(new_n826), .A2(new_n827), .A3(new_n679), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n527), .A2(new_n684), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n827), .B1(new_n826), .B2(new_n679), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n823), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(G137), .ZN(G39));
  NAND3_X1  g647(.A1(new_n829), .A2(new_n681), .A3(new_n752), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(new_n758), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n822), .A2(KEYINPUT47), .A3(new_n188), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT47), .B1(new_n822), .B2(new_n188), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n835), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(G140), .ZN(G42));
  AND3_X1   g654(.A1(new_n778), .A2(new_n829), .A3(new_n431), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n841), .A2(new_n796), .A3(new_n825), .ZN(new_n842));
  XOR2_X1   g656(.A(new_n842), .B(KEYINPUT48), .Z(new_n843));
  INV_X1    g657(.A(G952), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n825), .A2(new_n431), .A3(new_n786), .ZN(new_n845));
  AOI211_X1 g659(.A(new_n844), .B(G953), .C1(new_n845), .C2(new_n768), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n745), .A2(new_n681), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n841), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n846), .B1(new_n694), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n843), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n188), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n766), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n837), .A2(new_n838), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n845), .A2(new_n829), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(KEYINPUT118), .Z(new_n856));
  NOR2_X1   g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n841), .A2(new_n703), .A3(new_n692), .A4(new_n847), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n719), .A2(new_n785), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n841), .A2(new_n859), .A3(new_n825), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT120), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n845), .A2(new_n684), .A3(new_n778), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT50), .B1(new_n733), .B2(new_n863), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n733), .A2(new_n863), .A3(KEYINPUT50), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n862), .B(KEYINPUT51), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n850), .B1(new_n857), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(KEYINPUT119), .B1(new_n854), .B2(new_n856), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n865), .A2(new_n864), .ZN(new_n869));
  INV_X1    g683(.A(new_n838), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n870), .A2(new_n836), .A3(new_n852), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n872));
  INV_X1    g686(.A(new_n856), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n861), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n868), .A2(new_n869), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT51), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n867), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT53), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n694), .A2(new_n704), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n668), .A2(new_n436), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n881), .A2(new_n679), .A3(new_n682), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n671), .A2(new_n721), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n791), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n795), .A2(new_n884), .ZN(new_n885));
  OR3_X1    g699(.A1(new_n366), .A2(new_n428), .A3(new_n726), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n680), .A2(new_n719), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n887), .A2(new_n758), .A3(new_n829), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n815), .A2(new_n885), .A3(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n883), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n772), .A2(new_n769), .A3(new_n775), .A4(new_n789), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n890), .A2(new_n813), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n316), .A2(new_n438), .A3(new_n686), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n894), .A2(new_n756), .A3(new_n757), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n792), .B1(new_n895), .B2(new_n728), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n718), .A2(new_n314), .A3(new_n726), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(new_n745), .A3(new_n788), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n896), .A2(KEYINPUT52), .A3(new_n754), .A4(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n768), .A2(new_n884), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n729), .A2(new_n754), .A3(new_n900), .A4(new_n898), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT114), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT52), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n899), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n901), .A2(KEYINPUT114), .A3(new_n903), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n879), .B1(new_n893), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n899), .A2(new_n904), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n890), .A2(new_n909), .A3(new_n813), .A4(new_n892), .ZN(new_n910));
  OAI22_X1  g724(.A1(new_n908), .A2(KEYINPUT115), .B1(new_n879), .B2(new_n910), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n908), .A2(KEYINPUT115), .ZN(new_n912));
  OAI21_X1  g726(.A(KEYINPUT54), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n905), .A2(new_n906), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n883), .A2(new_n889), .A3(new_n879), .ZN(new_n915));
  INV_X1    g729(.A(new_n800), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n803), .A2(new_n810), .A3(new_n797), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT42), .B1(new_n917), .B2(KEYINPUT111), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n758), .A2(new_n795), .A3(new_n649), .A4(new_n752), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT111), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n916), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(KEYINPUT116), .B1(new_n922), .B2(new_n891), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT116), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n813), .A2(new_n924), .A3(new_n892), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n914), .A2(new_n915), .A3(new_n923), .A4(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT54), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n910), .A2(new_n879), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT117), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n929), .A2(new_n930), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n878), .B(new_n913), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n844), .A2(new_n430), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n766), .B(KEYINPUT49), .Z(new_n936));
  NOR4_X1   g750(.A1(new_n936), .A2(new_n684), .A3(new_n851), .A4(new_n824), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n733), .A2(new_n847), .A3(new_n937), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT113), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n935), .A2(new_n939), .ZN(G75));
  XNOR2_X1  g754(.A(new_n500), .B(KEYINPUT121), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT55), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n915), .A2(new_n905), .A3(new_n906), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n921), .A2(new_n798), .A3(new_n801), .ZN(new_n945));
  AOI211_X1 g759(.A(KEYINPUT116), .B(new_n891), .C1(new_n945), .C2(new_n800), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n924), .B1(new_n813), .B2(new_n892), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n944), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n910), .A2(new_n879), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n306), .B(new_n522), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT56), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n950), .A2(new_n951), .A3(new_n508), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n508), .B1(new_n950), .B2(new_n951), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n943), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n950), .A2(new_n951), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n509), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n950), .A2(new_n951), .A3(new_n508), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n956), .A2(new_n957), .A3(new_n942), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n430), .A2(G952), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n954), .A2(new_n958), .A3(new_n960), .ZN(G51));
  AOI211_X1 g775(.A(KEYINPUT122), .B(new_n927), .C1(new_n926), .C2(new_n928), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n926), .A2(new_n928), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(KEYINPUT54), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT122), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n929), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n962), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(G469), .A2(G902), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT57), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n759), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n948), .A2(new_n949), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n971), .A2(new_n305), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n817), .A2(G469), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT123), .Z(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n959), .B1(new_n970), .B2(new_n975), .ZN(G54));
  NAND3_X1  g790(.A1(new_n972), .A2(KEYINPUT58), .A3(G475), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n419), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n960), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n977), .A2(new_n419), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(new_n980), .ZN(G60));
  NAND2_X1  g795(.A1(new_n688), .A2(new_n690), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n913), .B1(new_n931), .B2(new_n932), .ZN(new_n983));
  NAND2_X1  g797(.A1(G478), .A2(G902), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT59), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n982), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n982), .A2(new_n985), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n960), .B1(new_n967), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n986), .A2(new_n988), .ZN(G63));
  XNOR2_X1  g803(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n348), .A2(new_n303), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n963), .A2(new_n713), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n993), .A2(KEYINPUT125), .A3(new_n960), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(KEYINPUT61), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n645), .A2(new_n647), .ZN(new_n996));
  INV_X1    g810(.A(new_n992), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n996), .B1(new_n971), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n998), .A2(new_n993), .A3(new_n960), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n995), .B(new_n999), .ZN(G66));
  OAI21_X1  g814(.A(G953), .B1(new_n434), .B2(new_n448), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n883), .A2(new_n891), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1001), .B1(new_n1002), .B2(G953), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n941), .B1(G898), .B2(new_n430), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1003), .B(new_n1004), .ZN(G69));
  XNOR2_X1  g819(.A(new_n584), .B(new_n410), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(new_n880), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n666), .A2(new_n736), .A3(new_n829), .A4(new_n1008), .ZN(new_n1009));
  AND3_X1   g823(.A1(new_n839), .A2(new_n832), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n896), .A2(new_n754), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(KEYINPUT62), .B1(new_n750), .B2(new_n1012), .ZN(new_n1013));
  AND3_X1   g827(.A1(new_n750), .A2(KEYINPUT62), .A3(new_n1012), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1010), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1007), .B1(new_n1015), .B2(new_n430), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n796), .A2(new_n788), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1012), .B1(new_n823), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n815), .B1(new_n823), .B2(new_n831), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1020), .A2(new_n813), .A3(new_n839), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1021), .A2(new_n430), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n430), .A2(G900), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1006), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n1016), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(G953), .B1(new_n277), .B2(new_n725), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n1027), .B(KEYINPUT126), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1026), .B(new_n1028), .ZN(G72));
  NAND2_X1  g843(.A1(G472), .A2(G902), .ZN(new_n1030));
  XOR2_X1   g844(.A(new_n1030), .B(KEYINPUT63), .Z(new_n1031));
  OR2_X1    g845(.A1(new_n883), .A2(new_n891), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1031), .B1(new_n1015), .B2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n590), .A2(new_n539), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n959), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n1020), .A2(new_n813), .A3(new_n839), .A4(new_n1002), .ZN(new_n1036));
  AND3_X1   g850(.A1(new_n1036), .A2(KEYINPUT127), .A3(new_n1031), .ZN(new_n1037));
  AOI21_X1  g851(.A(KEYINPUT127), .B1(new_n1036), .B2(new_n1031), .ZN(new_n1038));
  OAI211_X1 g852(.A(new_n539), .B(new_n590), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n587), .A2(new_n562), .ZN(new_n1040));
  OAI211_X1 g854(.A(new_n1031), .B(new_n1040), .C1(new_n911), .C2(new_n912), .ZN(new_n1041));
  AND3_X1   g855(.A1(new_n1035), .A2(new_n1039), .A3(new_n1041), .ZN(G57));
endmodule


