

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749;

  XNOR2_X1 U376 ( .A(n386), .B(n357), .ZN(n364) );
  INV_X1 U377 ( .A(n385), .ZN(n357) );
  OR2_X1 U378 ( .A1(n600), .A2(n601), .ZN(n404) );
  XNOR2_X1 U379 ( .A(n582), .B(n581), .ZN(n744) );
  XNOR2_X1 U380 ( .A(n577), .B(KEYINPUT33), .ZN(n695) );
  AND2_X1 U381 ( .A1(n602), .A2(n597), .ZN(n577) );
  AND2_X1 U382 ( .A1(n355), .A2(n647), .ZN(n560) );
  INV_X1 U383 ( .A(n535), .ZN(n356) );
  NOR2_X1 U384 ( .A1(n675), .A2(n539), .ZN(n607) );
  XNOR2_X1 U385 ( .A(n479), .B(n478), .ZN(n540) );
  AND2_X1 U386 ( .A1(n419), .A2(n418), .ZN(n417) );
  XNOR2_X1 U387 ( .A(n428), .B(n486), .ZN(n732) );
  XNOR2_X1 U388 ( .A(n400), .B(n399), .ZN(n403) );
  INV_X2 U389 ( .A(G953), .ZN(n736) );
  XNOR2_X2 U390 ( .A(n354), .B(n368), .ZN(n530) );
  NAND2_X1 U391 ( .A1(n367), .A2(n361), .ZN(n354) );
  AND2_X1 U392 ( .A1(n597), .A2(n356), .ZN(n355) );
  NAND2_X2 U393 ( .A1(n376), .A2(n665), .ZN(n562) );
  OR2_X2 U394 ( .A1(n584), .A2(n535), .ZN(n536) );
  INV_X2 U395 ( .A(n606), .ZN(n603) );
  NAND2_X1 U396 ( .A1(n358), .A2(n643), .ZN(n559) );
  NAND2_X1 U397 ( .A1(n549), .A2(n550), .ZN(n358) );
  NAND2_X2 U398 ( .A1(n384), .A2(n411), .ZN(n382) );
  NOR2_X1 U399 ( .A1(G953), .A2(G237), .ZN(n469) );
  AND2_X2 U400 ( .A1(n412), .A2(n410), .ZN(n384) );
  AND2_X2 U401 ( .A1(n414), .A2(n413), .ZN(n391) );
  XNOR2_X2 U402 ( .A(n377), .B(n453), .ZN(n516) );
  XNOR2_X2 U403 ( .A(n377), .B(n499), .ZN(n708) );
  NOR2_X1 U404 ( .A1(n564), .A2(n676), .ZN(n653) );
  INV_X1 U405 ( .A(KEYINPUT4), .ZN(n399) );
  NOR2_X1 U406 ( .A1(n565), .A2(n653), .ZN(n566) );
  XNOR2_X1 U407 ( .A(n465), .B(G140), .ZN(n428) );
  XNOR2_X1 U408 ( .A(n450), .B(G128), .ZN(n455) );
  XOR2_X1 U409 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n465) );
  BUF_X1 U410 ( .A(n722), .Z(n359) );
  XNOR2_X1 U411 ( .A(n576), .B(n439), .ZN(n360) );
  XNOR2_X1 U412 ( .A(n576), .B(n439), .ZN(n606) );
  XNOR2_X2 U413 ( .A(G101), .B(G110), .ZN(n480) );
  XNOR2_X1 U414 ( .A(n607), .B(KEYINPUT108), .ZN(n381) );
  NAND2_X1 U415 ( .A1(G214), .A2(n518), .ZN(n665) );
  INV_X1 U416 ( .A(KEYINPUT73), .ZN(n521) );
  INV_X1 U417 ( .A(n392), .ZN(n601) );
  INV_X1 U418 ( .A(KEYINPUT98), .ZN(n409) );
  NAND2_X1 U419 ( .A1(G469), .A2(n416), .ZN(n415) );
  INV_X1 U420 ( .A(G902), .ZN(n416) );
  NAND2_X1 U421 ( .A1(n420), .A2(G902), .ZN(n418) );
  XNOR2_X1 U422 ( .A(n568), .B(KEYINPUT84), .ZN(n569) );
  XNOR2_X1 U423 ( .A(G116), .B(G113), .ZN(n445) );
  XNOR2_X1 U424 ( .A(G137), .B(G134), .ZN(n451) );
  XOR2_X1 U425 ( .A(KEYINPUT70), .B(G131), .Z(n452) );
  INV_X1 U426 ( .A(KEYINPUT67), .ZN(n385) );
  XNOR2_X1 U427 ( .A(n511), .B(n510), .ZN(n678) );
  NOR2_X1 U428 ( .A1(n719), .A2(G902), .ZN(n511) );
  XNOR2_X1 U429 ( .A(n505), .B(KEYINPUT24), .ZN(n431) );
  XNOR2_X1 U430 ( .A(G119), .B(G110), .ZN(n505) );
  XNOR2_X1 U431 ( .A(KEYINPUT81), .B(KEYINPUT8), .ZN(n458) );
  XNOR2_X1 U432 ( .A(G113), .B(G131), .ZN(n472) );
  INV_X1 U433 ( .A(KEYINPUT112), .ZN(n388) );
  XOR2_X1 U434 ( .A(n519), .B(KEYINPUT30), .Z(n361) );
  INV_X1 U435 ( .A(n522), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n492), .B(n494), .ZN(n441) );
  XNOR2_X1 U437 ( .A(G478), .B(n464), .ZN(n552) );
  XNOR2_X1 U438 ( .A(n440), .B(KEYINPUT0), .ZN(n439) );
  INV_X1 U439 ( .A(KEYINPUT66), .ZN(n440) );
  XNOR2_X1 U440 ( .A(n427), .B(n370), .ZN(n426) );
  INV_X1 U441 ( .A(KEYINPUT86), .ZN(n598) );
  OR2_X1 U442 ( .A1(KEYINPUT47), .A2(n645), .ZN(n549) );
  INV_X1 U443 ( .A(G143), .ZN(n450) );
  OR2_X1 U444 ( .A1(G237), .A2(G902), .ZN(n518) );
  XOR2_X1 U445 ( .A(G101), .B(KEYINPUT5), .Z(n448) );
  XOR2_X1 U446 ( .A(G122), .B(G134), .Z(n461) );
  XNOR2_X1 U447 ( .A(n455), .B(n394), .ZN(n456) );
  XNOR2_X1 U448 ( .A(G116), .B(G107), .ZN(n394) );
  XNOR2_X1 U449 ( .A(G143), .B(G104), .ZN(n466) );
  XOR2_X1 U450 ( .A(KEYINPUT100), .B(G122), .Z(n467) );
  XNOR2_X1 U451 ( .A(n389), .B(n471), .ZN(n473) );
  XOR2_X1 U452 ( .A(KEYINPUT12), .B(KEYINPUT99), .Z(n471) );
  XNOR2_X1 U453 ( .A(n470), .B(n390), .ZN(n389) );
  INV_X1 U454 ( .A(KEYINPUT11), .ZN(n390) );
  XNOR2_X1 U455 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n484) );
  XNOR2_X1 U456 ( .A(n486), .B(n374), .ZN(n373) );
  AND2_X1 U457 ( .A1(n736), .A2(G224), .ZN(n374) );
  NAND2_X1 U458 ( .A1(G234), .A2(G237), .ZN(n512) );
  INV_X1 U459 ( .A(KEYINPUT76), .ZN(n398) );
  INV_X1 U460 ( .A(n655), .ZN(n395) );
  XNOR2_X1 U461 ( .A(n432), .B(n446), .ZN(n482) );
  XNOR2_X1 U462 ( .A(n445), .B(n444), .ZN(n432) );
  INV_X1 U463 ( .A(KEYINPUT3), .ZN(n444) );
  XNOR2_X1 U464 ( .A(G902), .B(KEYINPUT15), .ZN(n491) );
  XNOR2_X1 U465 ( .A(n588), .B(n589), .ZN(n593) );
  BUF_X1 U466 ( .A(n678), .Z(n392) );
  NOR2_X1 U467 ( .A1(G902), .A2(n712), .ZN(n479) );
  XNOR2_X1 U468 ( .A(n682), .B(n369), .ZN(n597) );
  NAND2_X1 U469 ( .A1(n593), .A2(n676), .ZN(n596) );
  XNOR2_X1 U470 ( .A(n433), .B(n482), .ZN(n728) );
  XNOR2_X1 U471 ( .A(n496), .B(n483), .ZN(n433) );
  XOR2_X1 U472 ( .A(G122), .B(KEYINPUT16), .Z(n483) );
  XNOR2_X1 U473 ( .A(n429), .B(n732), .ZN(n719) );
  XNOR2_X1 U474 ( .A(n623), .B(KEYINPUT122), .ZN(n625) );
  XNOR2_X1 U475 ( .A(n712), .B(n443), .ZN(n713) );
  XNOR2_X1 U476 ( .A(n531), .B(KEYINPUT40), .ZN(n532) );
  INV_X1 U477 ( .A(KEYINPUT111), .ZN(n531) );
  INV_X1 U478 ( .A(KEYINPUT36), .ZN(n393) );
  INV_X1 U479 ( .A(KEYINPUT35), .ZN(n581) );
  NAND2_X1 U480 ( .A1(n361), .A2(n365), .ZN(n554) );
  NOR2_X1 U481 ( .A1(n682), .A2(n608), .ZN(n632) );
  NAND2_X1 U482 ( .A1(n426), .A2(n436), .ZN(n425) );
  INV_X1 U483 ( .A(KEYINPUT56), .ZN(n434) );
  NAND2_X1 U484 ( .A1(n437), .A2(n436), .ZN(n435) );
  XNOR2_X1 U485 ( .A(n438), .B(n371), .ZN(n437) );
  INV_X1 U486 ( .A(n404), .ZN(n629) );
  XOR2_X1 U487 ( .A(KEYINPUT87), .B(n612), .Z(n362) );
  AND2_X1 U488 ( .A1(n613), .A2(KEYINPUT44), .ZN(n363) );
  AND2_X1 U489 ( .A1(n381), .A2(n378), .ZN(n365) );
  NOR2_X1 U490 ( .A1(n529), .A2(n376), .ZN(n366) );
  INV_X1 U491 ( .A(G469), .ZN(n420) );
  AND2_X1 U492 ( .A1(n381), .A2(n379), .ZN(n367) );
  XOR2_X1 U493 ( .A(n521), .B(KEYINPUT39), .Z(n368) );
  XOR2_X1 U494 ( .A(KEYINPUT104), .B(KEYINPUT6), .Z(n369) );
  INV_X1 U495 ( .A(KEYINPUT1), .ZN(n413) );
  XOR2_X1 U496 ( .A(n454), .B(n516), .Z(n370) );
  XOR2_X1 U497 ( .A(n704), .B(n703), .Z(n371) );
  NOR2_X1 U498 ( .A1(G952), .A2(n736), .ZN(n721) );
  INV_X1 U499 ( .A(n721), .ZN(n436) );
  XOR2_X1 U500 ( .A(n622), .B(KEYINPUT88), .Z(n372) );
  INV_X2 U501 ( .A(G125), .ZN(n375) );
  XNOR2_X1 U502 ( .A(n487), .B(n373), .ZN(n489) );
  XNOR2_X2 U503 ( .A(n375), .B(G146), .ZN(n486) );
  XNOR2_X1 U504 ( .A(n376), .B(n495), .ZN(n666) );
  NAND2_X1 U505 ( .A1(n555), .A2(n376), .ZN(n643) );
  XNOR2_X2 U506 ( .A(n493), .B(n441), .ZN(n376) );
  XNOR2_X2 U507 ( .A(n733), .B(G146), .ZN(n377) );
  OR2_X2 U508 ( .A1(n708), .A2(n415), .ZN(n414) );
  NOR2_X1 U509 ( .A1(n520), .A2(n522), .ZN(n379) );
  XNOR2_X2 U510 ( .A(n382), .B(n398), .ZN(n602) );
  NAND2_X1 U511 ( .A1(n383), .A2(KEYINPUT1), .ZN(n411) );
  NAND2_X1 U512 ( .A1(n417), .A2(n414), .ZN(n383) );
  NAND2_X1 U513 ( .A1(n391), .A2(n417), .ZN(n412) );
  XNOR2_X1 U514 ( .A(n560), .B(n388), .ZN(n561) );
  INV_X1 U515 ( .A(n534), .ZN(n682) );
  XOR2_X2 U516 ( .A(G104), .B(G107), .Z(n481) );
  NAND2_X1 U517 ( .A1(n744), .A2(n583), .ZN(n386) );
  NOR2_X1 U518 ( .A1(n695), .A2(n603), .ZN(n578) );
  NAND2_X1 U519 ( .A1(n702), .A2(n618), .ZN(n493) );
  XNOR2_X1 U520 ( .A(n728), .B(n490), .ZN(n702) );
  INV_X1 U521 ( .A(n366), .ZN(n422) );
  AND2_X2 U522 ( .A1(n396), .A2(n395), .ZN(n734) );
  OR2_X2 U523 ( .A1(n559), .A2(n558), .ZN(n565) );
  NOR2_X2 U524 ( .A1(n542), .A2(n694), .ZN(n543) );
  NAND2_X1 U525 ( .A1(n602), .A2(n682), .ZN(n685) );
  XNOR2_X1 U526 ( .A(n624), .B(n625), .ZN(n626) );
  AND2_X4 U527 ( .A1(n621), .A2(n620), .ZN(n717) );
  XNOR2_X1 U528 ( .A(n387), .B(n532), .ZN(n748) );
  NOR2_X1 U529 ( .A1(n530), .A2(n547), .ZN(n387) );
  NAND2_X2 U530 ( .A1(n722), .A2(n734), .ZN(n656) );
  XNOR2_X2 U531 ( .A(n656), .B(n617), .ZN(n621) );
  XNOR2_X2 U532 ( .A(n481), .B(n480), .ZN(n496) );
  XNOR2_X1 U533 ( .A(n421), .B(KEYINPUT83), .ZN(n396) );
  XNOR2_X1 U534 ( .A(n517), .B(G472), .ZN(n534) );
  XNOR2_X1 U535 ( .A(n488), .B(n489), .ZN(n490) );
  XNOR2_X1 U536 ( .A(n563), .B(n393), .ZN(n564) );
  NAND2_X1 U537 ( .A1(n364), .A2(n362), .ZN(n616) );
  NAND2_X1 U538 ( .A1(n574), .A2(n575), .ZN(n576) );
  XNOR2_X2 U539 ( .A(n562), .B(KEYINPUT19), .ZN(n574) );
  NAND2_X1 U540 ( .A1(n717), .A2(G478), .ZN(n624) );
  XNOR2_X2 U541 ( .A(n397), .B(KEYINPUT45), .ZN(n722) );
  NAND2_X1 U542 ( .A1(n615), .A2(n616), .ZN(n397) );
  AND2_X2 U543 ( .A1(n405), .A2(n404), .ZN(n611) );
  XNOR2_X1 U544 ( .A(n504), .B(n431), .ZN(n430) );
  XNOR2_X1 U545 ( .A(n430), .B(n507), .ZN(n429) );
  XNOR2_X2 U546 ( .A(KEYINPUT65), .B(KEYINPUT68), .ZN(n400) );
  NAND2_X1 U547 ( .A1(n401), .A2(n662), .ZN(n664) );
  NAND2_X1 U548 ( .A1(n659), .A2(KEYINPUT82), .ZN(n401) );
  NOR2_X1 U549 ( .A1(n596), .A2(n597), .ZN(n599) );
  XNOR2_X1 U550 ( .A(n402), .B(n716), .ZN(G60) );
  NOR2_X2 U551 ( .A1(n715), .A2(n721), .ZN(n402) );
  NAND2_X1 U552 ( .A1(n360), .A2(n587), .ZN(n588) );
  XNOR2_X2 U553 ( .A(n488), .B(n442), .ZN(n733) );
  XNOR2_X2 U554 ( .A(n403), .B(n455), .ZN(n488) );
  XNOR2_X1 U555 ( .A(n406), .B(n610), .ZN(n405) );
  NAND2_X1 U556 ( .A1(n408), .A2(n407), .ZN(n406) );
  INV_X1 U557 ( .A(n671), .ZN(n407) );
  XNOR2_X1 U558 ( .A(n609), .B(n409), .ZN(n408) );
  INV_X1 U559 ( .A(n675), .ZN(n410) );
  NAND2_X1 U560 ( .A1(n411), .A2(n412), .ZN(n676) );
  NAND2_X1 U561 ( .A1(n417), .A2(n414), .ZN(n539) );
  NAND2_X1 U562 ( .A1(n708), .A2(n420), .ZN(n419) );
  NOR2_X1 U563 ( .A1(n614), .A2(n363), .ZN(n615) );
  NOR2_X2 U564 ( .A1(n603), .A2(n685), .ZN(n605) );
  NAND2_X1 U565 ( .A1(n423), .A2(n422), .ZN(n421) );
  XNOR2_X1 U566 ( .A(n424), .B(n569), .ZN(n423) );
  NAND2_X1 U567 ( .A1(n566), .A2(n567), .ZN(n424) );
  XNOR2_X1 U568 ( .A(n425), .B(n372), .ZN(G57) );
  NAND2_X1 U569 ( .A1(n717), .A2(G472), .ZN(n427) );
  NAND2_X1 U570 ( .A1(n678), .A2(n679), .ZN(n675) );
  XNOR2_X1 U571 ( .A(n435), .B(n434), .ZN(G51) );
  NAND2_X1 U572 ( .A1(n717), .A2(G210), .ZN(n438) );
  XOR2_X1 U573 ( .A(n452), .B(n451), .Z(n442) );
  XNOR2_X1 U574 ( .A(KEYINPUT59), .B(KEYINPUT91), .ZN(n443) );
  INV_X1 U575 ( .A(KEYINPUT103), .ZN(n610) );
  XNOR2_X1 U576 ( .A(n656), .B(KEYINPUT77), .ZN(n657) );
  INV_X1 U577 ( .A(G475), .ZN(n476) );
  INV_X1 U578 ( .A(n676), .ZN(n527) );
  XNOR2_X1 U579 ( .A(n477), .B(n476), .ZN(n478) );
  INV_X1 U580 ( .A(KEYINPUT63), .ZN(n622) );
  XNOR2_X1 U581 ( .A(n714), .B(n713), .ZN(n715) );
  INV_X1 U582 ( .A(KEYINPUT123), .ZN(n627) );
  XNOR2_X1 U583 ( .A(KEYINPUT62), .B(KEYINPUT90), .ZN(n454) );
  XOR2_X1 U584 ( .A(KEYINPUT72), .B(G119), .Z(n446) );
  NAND2_X1 U585 ( .A1(n469), .A2(G210), .ZN(n447) );
  XNOR2_X1 U586 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U587 ( .A(n482), .B(n449), .ZN(n453) );
  XNOR2_X1 U588 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n457) );
  XNOR2_X1 U589 ( .A(n457), .B(n456), .ZN(n463) );
  NAND2_X1 U590 ( .A1(n736), .A2(G234), .ZN(n459) );
  XNOR2_X1 U591 ( .A(n459), .B(n458), .ZN(n506) );
  NAND2_X1 U592 ( .A1(G217), .A2(n506), .ZN(n460) );
  XNOR2_X1 U593 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U594 ( .A(n463), .B(n462), .ZN(n623) );
  NOR2_X1 U595 ( .A1(G902), .A2(n623), .ZN(n464) );
  XNOR2_X1 U596 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U597 ( .A(n732), .B(n468), .ZN(n475) );
  NAND2_X1 U598 ( .A1(G214), .A2(n469), .ZN(n470) );
  XNOR2_X1 U599 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U600 ( .A(n475), .B(n474), .ZN(n712) );
  XNOR2_X1 U601 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n477) );
  NOR2_X1 U602 ( .A1(n552), .A2(n540), .ZN(n650) );
  INV_X1 U603 ( .A(n650), .ZN(n637) );
  INV_X1 U604 ( .A(KEYINPUT38), .ZN(n495) );
  XOR2_X1 U605 ( .A(KEYINPUT93), .B(KEYINPUT78), .Z(n485) );
  XNOR2_X1 U606 ( .A(n485), .B(n484), .ZN(n487) );
  XNOR2_X1 U607 ( .A(n491), .B(KEYINPUT92), .ZN(n618) );
  NAND2_X1 U608 ( .A1(G210), .A2(n518), .ZN(n492) );
  XNOR2_X1 U609 ( .A(KEYINPUT94), .B(KEYINPUT79), .ZN(n494) );
  INV_X1 U610 ( .A(n666), .ZN(n520) );
  XOR2_X1 U611 ( .A(n496), .B(G140), .Z(n498) );
  NAND2_X1 U612 ( .A1(G227), .A2(n736), .ZN(n497) );
  XNOR2_X1 U613 ( .A(n498), .B(n497), .ZN(n499) );
  NAND2_X1 U614 ( .A1(n618), .A2(G234), .ZN(n500) );
  XNOR2_X1 U615 ( .A(KEYINPUT20), .B(n500), .ZN(n508) );
  NAND2_X1 U616 ( .A1(n508), .A2(G221), .ZN(n501) );
  XNOR2_X1 U617 ( .A(KEYINPUT21), .B(n501), .ZN(n586) );
  INV_X1 U618 ( .A(n586), .ZN(n679) );
  XOR2_X1 U619 ( .A(KEYINPUT23), .B(KEYINPUT96), .Z(n503) );
  XNOR2_X1 U620 ( .A(G128), .B(G137), .ZN(n502) );
  XNOR2_X1 U621 ( .A(n503), .B(n502), .ZN(n504) );
  NAND2_X1 U622 ( .A1(G221), .A2(n506), .ZN(n507) );
  NAND2_X1 U623 ( .A1(G217), .A2(n508), .ZN(n509) );
  XNOR2_X1 U624 ( .A(n509), .B(KEYINPUT25), .ZN(n510) );
  XNOR2_X1 U625 ( .A(KEYINPUT14), .B(n512), .ZN(n514) );
  AND2_X1 U626 ( .A1(G953), .A2(n514), .ZN(n513) );
  NAND2_X1 U627 ( .A1(G902), .A2(n513), .ZN(n570) );
  NOR2_X1 U628 ( .A1(G900), .A2(n570), .ZN(n515) );
  NAND2_X1 U629 ( .A1(G952), .A2(n514), .ZN(n693) );
  NOR2_X1 U630 ( .A1(G953), .A2(n693), .ZN(n572) );
  NOR2_X1 U631 ( .A1(n515), .A2(n572), .ZN(n522) );
  NOR2_X1 U632 ( .A1(G902), .A2(n516), .ZN(n517) );
  NAND2_X1 U633 ( .A1(n682), .A2(n665), .ZN(n519) );
  NOR2_X1 U634 ( .A1(n637), .A2(n530), .ZN(n655) );
  NOR2_X1 U635 ( .A1(n522), .A2(n678), .ZN(n523) );
  NAND2_X1 U636 ( .A1(n523), .A2(n679), .ZN(n535) );
  NAND2_X1 U637 ( .A1(n552), .A2(n540), .ZN(n524) );
  XNOR2_X2 U638 ( .A(n524), .B(KEYINPUT102), .ZN(n547) );
  XNOR2_X2 U639 ( .A(n547), .B(KEYINPUT107), .ZN(n647) );
  NAND2_X1 U640 ( .A1(n560), .A2(n665), .ZN(n526) );
  NOR2_X1 U641 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U642 ( .A(n528), .B(KEYINPUT43), .ZN(n529) );
  XNOR2_X1 U643 ( .A(KEYINPUT28), .B(KEYINPUT110), .ZN(n533) );
  XNOR2_X1 U644 ( .A(n533), .B(KEYINPUT109), .ZN(n537) );
  BUF_X1 U645 ( .A(n534), .Z(n584) );
  XOR2_X1 U646 ( .A(n537), .B(n536), .Z(n538) );
  NOR2_X1 U647 ( .A1(n539), .A2(n538), .ZN(n548) );
  INV_X1 U648 ( .A(n548), .ZN(n542) );
  INV_X1 U649 ( .A(n540), .ZN(n551) );
  NAND2_X1 U650 ( .A1(n552), .A2(n551), .ZN(n669) );
  NAND2_X1 U651 ( .A1(n666), .A2(n665), .ZN(n670) );
  NOR2_X1 U652 ( .A1(n669), .A2(n670), .ZN(n541) );
  XNOR2_X1 U653 ( .A(n541), .B(KEYINPUT41), .ZN(n694) );
  XNOR2_X1 U654 ( .A(n543), .B(KEYINPUT42), .ZN(n747) );
  NOR2_X1 U655 ( .A1(n748), .A2(n747), .ZN(n546) );
  XOR2_X1 U656 ( .A(KEYINPUT46), .B(KEYINPUT85), .Z(n544) );
  XNOR2_X1 U657 ( .A(KEYINPUT64), .B(n544), .ZN(n545) );
  XNOR2_X1 U658 ( .A(n546), .B(n545), .ZN(n567) );
  AND2_X1 U659 ( .A1(n547), .A2(n637), .ZN(n671) );
  XNOR2_X1 U660 ( .A(KEYINPUT47), .B(n671), .ZN(n550) );
  NAND2_X1 U661 ( .A1(n548), .A2(n574), .ZN(n638) );
  INV_X1 U662 ( .A(n638), .ZN(n645) );
  NOR2_X1 U663 ( .A1(n552), .A2(n551), .ZN(n579) );
  INV_X1 U664 ( .A(n579), .ZN(n553) );
  NOR2_X1 U665 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U666 ( .A1(n638), .A2(KEYINPUT47), .ZN(n557) );
  XOR2_X1 U667 ( .A(KEYINPUT80), .B(n557), .Z(n558) );
  NOR2_X1 U668 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U669 ( .A(KEYINPUT48), .B(KEYINPUT71), .ZN(n568) );
  NOR2_X1 U670 ( .A1(G898), .A2(n570), .ZN(n571) );
  NOR2_X1 U671 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U672 ( .A(KEYINPUT95), .B(n573), .ZN(n575) );
  XNOR2_X1 U673 ( .A(n578), .B(KEYINPUT34), .ZN(n580) );
  NAND2_X1 U674 ( .A1(n580), .A2(n579), .ZN(n582) );
  INV_X1 U675 ( .A(KEYINPUT44), .ZN(n583) );
  NAND2_X1 U676 ( .A1(n601), .A2(n584), .ZN(n591) );
  XNOR2_X1 U677 ( .A(KEYINPUT75), .B(KEYINPUT22), .ZN(n585) );
  XNOR2_X1 U678 ( .A(n585), .B(KEYINPUT74), .ZN(n589) );
  NOR2_X1 U679 ( .A1(n669), .A2(n586), .ZN(n587) );
  XNOR2_X1 U680 ( .A(KEYINPUT106), .B(n596), .ZN(n590) );
  NOR2_X1 U681 ( .A1(n591), .A2(n590), .ZN(n636) );
  NOR2_X1 U682 ( .A1(n676), .A2(n597), .ZN(n592) );
  NAND2_X1 U683 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U684 ( .A1(n594), .A2(n392), .ZN(n595) );
  XNOR2_X1 U685 ( .A(n595), .B(KEYINPUT32), .ZN(n746) );
  NOR2_X1 U686 ( .A1(n636), .A2(n746), .ZN(n612) );
  XNOR2_X1 U687 ( .A(n599), .B(n598), .ZN(n600) );
  XNOR2_X1 U688 ( .A(KEYINPUT31), .B(KEYINPUT97), .ZN(n604) );
  XNOR2_X1 U689 ( .A(n605), .B(n604), .ZN(n651) );
  NAND2_X1 U690 ( .A1(n607), .A2(n360), .ZN(n608) );
  NOR2_X1 U691 ( .A1(n651), .A2(n632), .ZN(n609) );
  XNOR2_X1 U692 ( .A(n611), .B(KEYINPUT105), .ZN(n614) );
  NAND2_X1 U693 ( .A1(n744), .A2(n612), .ZN(n613) );
  INV_X1 U694 ( .A(KEYINPUT2), .ZN(n658) );
  NOR2_X1 U695 ( .A1(KEYINPUT77), .A2(n658), .ZN(n617) );
  AND2_X1 U696 ( .A1(KEYINPUT77), .A2(n658), .ZN(n619) );
  NOR2_X1 U697 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X2 U698 ( .A1(n626), .A2(n721), .ZN(n628) );
  XNOR2_X1 U699 ( .A(n628), .B(n627), .ZN(G63) );
  XOR2_X1 U700 ( .A(G101), .B(n629), .Z(G3) );
  XOR2_X1 U701 ( .A(G104), .B(KEYINPUT113), .Z(n631) );
  NAND2_X1 U702 ( .A1(n632), .A2(n647), .ZN(n630) );
  XNOR2_X1 U703 ( .A(n631), .B(n630), .ZN(G6) );
  XOR2_X1 U704 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n634) );
  NAND2_X1 U705 ( .A1(n632), .A2(n650), .ZN(n633) );
  XNOR2_X1 U706 ( .A(n634), .B(n633), .ZN(n635) );
  XNOR2_X1 U707 ( .A(G107), .B(n635), .ZN(G9) );
  XOR2_X1 U708 ( .A(n636), .B(G110), .Z(G12) );
  NOR2_X1 U709 ( .A1(n638), .A2(n637), .ZN(n642) );
  XOR2_X1 U710 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n640) );
  XNOR2_X1 U711 ( .A(G128), .B(KEYINPUT115), .ZN(n639) );
  XNOR2_X1 U712 ( .A(n640), .B(n639), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n642), .B(n641), .ZN(G30) );
  XNOR2_X1 U714 ( .A(G143), .B(KEYINPUT116), .ZN(n644) );
  XNOR2_X1 U715 ( .A(n644), .B(n643), .ZN(G45) );
  NAND2_X1 U716 ( .A1(n647), .A2(n645), .ZN(n646) );
  XNOR2_X1 U717 ( .A(n646), .B(G146), .ZN(G48) );
  XOR2_X1 U718 ( .A(G113), .B(KEYINPUT117), .Z(n649) );
  NAND2_X1 U719 ( .A1(n651), .A2(n647), .ZN(n648) );
  XNOR2_X1 U720 ( .A(n649), .B(n648), .ZN(G15) );
  NAND2_X1 U721 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U722 ( .A(n652), .B(G116), .ZN(G18) );
  XNOR2_X1 U723 ( .A(n653), .B(G125), .ZN(n654) );
  XNOR2_X1 U724 ( .A(n654), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U725 ( .A(G134), .B(n655), .Z(G36) );
  XOR2_X1 U726 ( .A(G140), .B(n366), .Z(G42) );
  NOR2_X1 U727 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U728 ( .A(KEYINPUT82), .B(n734), .ZN(n661) );
  NOR2_X1 U729 ( .A1(KEYINPUT77), .A2(KEYINPUT2), .ZN(n660) );
  NAND2_X1 U730 ( .A1(n661), .A2(n660), .ZN(n662) );
  OR2_X1 U731 ( .A1(n359), .A2(KEYINPUT2), .ZN(n663) );
  NAND2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n699) );
  NOR2_X1 U733 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U734 ( .A(n667), .B(KEYINPUT118), .ZN(n668) );
  NOR2_X1 U735 ( .A1(n669), .A2(n668), .ZN(n673) );
  NOR2_X1 U736 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U737 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U738 ( .A1(n674), .A2(n695), .ZN(n690) );
  NAND2_X1 U739 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U740 ( .A(n677), .B(KEYINPUT50), .ZN(n684) );
  NOR2_X1 U741 ( .A1(n679), .A2(n392), .ZN(n680) );
  XOR2_X1 U742 ( .A(KEYINPUT49), .B(n680), .Z(n681) );
  NOR2_X1 U743 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U744 ( .A1(n684), .A2(n683), .ZN(n686) );
  NAND2_X1 U745 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U746 ( .A(KEYINPUT51), .B(n687), .ZN(n688) );
  NOR2_X1 U747 ( .A1(n694), .A2(n688), .ZN(n689) );
  NOR2_X1 U748 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U749 ( .A(n691), .B(KEYINPUT52), .ZN(n692) );
  NOR2_X1 U750 ( .A1(n693), .A2(n692), .ZN(n697) );
  NOR2_X1 U751 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U752 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U753 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U754 ( .A1(n700), .A2(G953), .ZN(n701) );
  XNOR2_X1 U755 ( .A(n701), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U756 ( .A(KEYINPUT89), .B(KEYINPUT55), .Z(n704) );
  XNOR2_X1 U757 ( .A(n702), .B(KEYINPUT54), .ZN(n703) );
  XOR2_X1 U758 ( .A(KEYINPUT120), .B(KEYINPUT119), .Z(n706) );
  XNOR2_X1 U759 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n705) );
  XNOR2_X1 U760 ( .A(n706), .B(n705), .ZN(n707) );
  XOR2_X1 U761 ( .A(n708), .B(n707), .Z(n710) );
  NAND2_X1 U762 ( .A1(n717), .A2(G469), .ZN(n709) );
  XNOR2_X1 U763 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U764 ( .A1(n721), .A2(n711), .ZN(G54) );
  NAND2_X1 U765 ( .A1(n717), .A2(G475), .ZN(n714) );
  XOR2_X1 U766 ( .A(KEYINPUT60), .B(KEYINPUT121), .Z(n716) );
  NAND2_X1 U767 ( .A1(G217), .A2(n717), .ZN(n718) );
  XNOR2_X1 U768 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U769 ( .A1(n721), .A2(n720), .ZN(G66) );
  NAND2_X1 U770 ( .A1(n736), .A2(n359), .ZN(n726) );
  NAND2_X1 U771 ( .A1(G953), .A2(G224), .ZN(n723) );
  XNOR2_X1 U772 ( .A(KEYINPUT61), .B(n723), .ZN(n724) );
  NAND2_X1 U773 ( .A1(n724), .A2(G898), .ZN(n725) );
  NAND2_X1 U774 ( .A1(n726), .A2(n725), .ZN(n730) );
  NOR2_X1 U775 ( .A1(G898), .A2(n736), .ZN(n727) );
  NOR2_X1 U776 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U777 ( .A(n730), .B(n729), .ZN(n731) );
  XNOR2_X1 U778 ( .A(KEYINPUT124), .B(n731), .ZN(G69) );
  XOR2_X1 U779 ( .A(n733), .B(n732), .Z(n739) );
  XNOR2_X1 U780 ( .A(n739), .B(n734), .ZN(n735) );
  XNOR2_X1 U781 ( .A(n735), .B(KEYINPUT125), .ZN(n737) );
  NAND2_X1 U782 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U783 ( .A(n738), .B(KEYINPUT126), .ZN(n743) );
  XNOR2_X1 U784 ( .A(G227), .B(n739), .ZN(n740) );
  NAND2_X1 U785 ( .A1(n740), .A2(G900), .ZN(n741) );
  NAND2_X1 U786 ( .A1(n741), .A2(G953), .ZN(n742) );
  NAND2_X1 U787 ( .A1(n743), .A2(n742), .ZN(G72) );
  INV_X1 U788 ( .A(n744), .ZN(n745) );
  XOR2_X1 U789 ( .A(G122), .B(n745), .Z(G24) );
  XOR2_X1 U790 ( .A(G119), .B(n746), .Z(G21) );
  XOR2_X1 U791 ( .A(n747), .B(G137), .Z(G39) );
  XNOR2_X1 U792 ( .A(G131), .B(KEYINPUT127), .ZN(n749) );
  XNOR2_X1 U793 ( .A(n749), .B(n748), .ZN(G33) );
endmodule

