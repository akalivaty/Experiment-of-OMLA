

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X4 U559 ( .A1(n537), .A2(n536), .ZN(G160) );
  NOR2_X1 U560 ( .A1(n699), .A2(n761), .ZN(n706) );
  INV_X1 U561 ( .A(KEYINPUT102), .ZN(n731) );
  XNOR2_X1 U562 ( .A(n731), .B(KEYINPUT31), .ZN(n732) );
  XNOR2_X1 U563 ( .A(n733), .B(n732), .ZN(n734) );
  OR2_X1 U564 ( .A1(n699), .A2(n761), .ZN(n738) );
  NOR2_X1 U565 ( .A1(G1966), .A2(n737), .ZN(n756) );
  XNOR2_X1 U566 ( .A(KEYINPUT104), .B(KEYINPUT32), .ZN(n746) );
  XNOR2_X1 U567 ( .A(n747), .B(n746), .ZN(n837) );
  NOR2_X1 U568 ( .A1(G651), .A2(n652), .ZN(n647) );
  INV_X1 U569 ( .A(KEYINPUT23), .ZN(n525) );
  INV_X1 U570 ( .A(G2104), .ZN(n530) );
  NOR2_X1 U571 ( .A1(n530), .A2(G2105), .ZN(n523) );
  XNOR2_X2 U572 ( .A(n523), .B(KEYINPUT64), .ZN(n899) );
  NAND2_X1 U573 ( .A1(G101), .A2(n899), .ZN(n524) );
  XNOR2_X1 U574 ( .A(n525), .B(n524), .ZN(n527) );
  INV_X1 U575 ( .A(G2105), .ZN(n529) );
  NOR2_X1 U576 ( .A1(G2104), .A2(n529), .ZN(n895) );
  NAND2_X1 U577 ( .A1(n895), .A2(G125), .ZN(n526) );
  NAND2_X1 U578 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U579 ( .A(n528), .B(KEYINPUT65), .ZN(n532) );
  NOR2_X1 U580 ( .A1(n530), .A2(n529), .ZN(n894) );
  NAND2_X1 U581 ( .A1(G113), .A2(n894), .ZN(n531) );
  NAND2_X1 U582 ( .A1(n532), .A2(n531), .ZN(n537) );
  NOR2_X1 U583 ( .A1(G2104), .A2(G2105), .ZN(n533) );
  XOR2_X1 U584 ( .A(KEYINPUT17), .B(n533), .Z(n534) );
  XNOR2_X2 U585 ( .A(KEYINPUT66), .B(n534), .ZN(n898) );
  NAND2_X1 U586 ( .A1(G137), .A2(n898), .ZN(n535) );
  XNOR2_X1 U587 ( .A(KEYINPUT67), .B(n535), .ZN(n536) );
  INV_X1 U588 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U589 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  INV_X1 U590 ( .A(G82), .ZN(G220) );
  INV_X1 U591 ( .A(G132), .ZN(G219) );
  NAND2_X1 U592 ( .A1(G69), .A2(G120), .ZN(n538) );
  NOR2_X1 U593 ( .A1(G237), .A2(n538), .ZN(n539) );
  NAND2_X1 U594 ( .A1(G108), .A2(n539), .ZN(n857) );
  NAND2_X1 U595 ( .A1(n857), .A2(G567), .ZN(n544) );
  NOR2_X1 U596 ( .A1(G220), .A2(G219), .ZN(n540) );
  XOR2_X1 U597 ( .A(KEYINPUT22), .B(n540), .Z(n541) );
  NOR2_X1 U598 ( .A1(G218), .A2(n541), .ZN(n542) );
  NAND2_X1 U599 ( .A1(G96), .A2(n542), .ZN(n858) );
  NAND2_X1 U600 ( .A1(n858), .A2(G2106), .ZN(n543) );
  AND2_X1 U601 ( .A1(n544), .A2(n543), .ZN(G319) );
  NOR2_X1 U602 ( .A1(G543), .A2(G651), .ZN(n637) );
  NAND2_X1 U603 ( .A1(n637), .A2(G90), .ZN(n546) );
  XOR2_X1 U604 ( .A(G543), .B(KEYINPUT0), .Z(n652) );
  XOR2_X1 U605 ( .A(KEYINPUT68), .B(G651), .Z(n550) );
  NOR2_X1 U606 ( .A1(n652), .A2(n550), .ZN(n638) );
  NAND2_X1 U607 ( .A1(G77), .A2(n638), .ZN(n545) );
  NAND2_X1 U608 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U609 ( .A(n547), .B(KEYINPUT9), .ZN(n549) );
  NAND2_X1 U610 ( .A1(G52), .A2(n647), .ZN(n548) );
  NAND2_X1 U611 ( .A1(n549), .A2(n548), .ZN(n554) );
  NOR2_X1 U612 ( .A1(G543), .A2(n550), .ZN(n551) );
  XOR2_X2 U613 ( .A(KEYINPUT1), .B(n551), .Z(n655) );
  NAND2_X1 U614 ( .A1(n655), .A2(G64), .ZN(n552) );
  XOR2_X1 U615 ( .A(KEYINPUT70), .B(n552), .Z(n553) );
  NOR2_X1 U616 ( .A1(n554), .A2(n553), .ZN(G171) );
  AND2_X1 U617 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U618 ( .A1(n894), .A2(G111), .ZN(n556) );
  NAND2_X1 U619 ( .A1(G135), .A2(n898), .ZN(n555) );
  NAND2_X1 U620 ( .A1(n556), .A2(n555), .ZN(n559) );
  NAND2_X1 U621 ( .A1(n895), .A2(G123), .ZN(n557) );
  XOR2_X1 U622 ( .A(KEYINPUT18), .B(n557), .Z(n558) );
  NOR2_X1 U623 ( .A1(n559), .A2(n558), .ZN(n561) );
  NAND2_X1 U624 ( .A1(G99), .A2(n899), .ZN(n560) );
  NAND2_X1 U625 ( .A1(n561), .A2(n560), .ZN(n941) );
  XNOR2_X1 U626 ( .A(G2096), .B(n941), .ZN(n562) );
  OR2_X1 U627 ( .A1(G2100), .A2(n562), .ZN(G156) );
  NAND2_X1 U628 ( .A1(G50), .A2(n647), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(KEYINPUT84), .ZN(n565) );
  NAND2_X1 U630 ( .A1(G75), .A2(n638), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n569) );
  NAND2_X1 U632 ( .A1(n637), .A2(G88), .ZN(n567) );
  NAND2_X1 U633 ( .A1(G62), .A2(n655), .ZN(n566) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(G166) );
  INV_X1 U636 ( .A(G166), .ZN(G303) );
  NAND2_X1 U637 ( .A1(n637), .A2(G89), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n570), .B(KEYINPUT4), .ZN(n572) );
  NAND2_X1 U639 ( .A1(G76), .A2(n638), .ZN(n571) );
  NAND2_X1 U640 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n573), .B(KEYINPUT5), .ZN(n578) );
  NAND2_X1 U642 ( .A1(G51), .A2(n647), .ZN(n575) );
  NAND2_X1 U643 ( .A1(G63), .A2(n655), .ZN(n574) );
  NAND2_X1 U644 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U645 ( .A(KEYINPUT6), .B(n576), .Z(n577) );
  NAND2_X1 U646 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U647 ( .A(n579), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U648 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U649 ( .A1(G7), .A2(G661), .ZN(n580) );
  XOR2_X1 U650 ( .A(n580), .B(KEYINPUT10), .Z(n853) );
  NAND2_X1 U651 ( .A1(n853), .A2(G567), .ZN(n581) );
  XOR2_X1 U652 ( .A(KEYINPUT11), .B(n581), .Z(G234) );
  NAND2_X1 U653 ( .A1(G81), .A2(n637), .ZN(n582) );
  XNOR2_X1 U654 ( .A(n582), .B(KEYINPUT12), .ZN(n583) );
  XNOR2_X1 U655 ( .A(n583), .B(KEYINPUT72), .ZN(n585) );
  NAND2_X1 U656 ( .A1(G68), .A2(n638), .ZN(n584) );
  NAND2_X1 U657 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U658 ( .A(n586), .B(KEYINPUT13), .ZN(n588) );
  NAND2_X1 U659 ( .A1(G43), .A2(n647), .ZN(n587) );
  NAND2_X1 U660 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n655), .A2(G56), .ZN(n589) );
  XOR2_X1 U662 ( .A(KEYINPUT14), .B(n589), .Z(n590) );
  NOR2_X1 U663 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U664 ( .A(KEYINPUT73), .B(n592), .Z(n999) );
  NAND2_X1 U665 ( .A1(n999), .A2(G860), .ZN(G153) );
  XOR2_X1 U666 ( .A(G171), .B(KEYINPUT74), .Z(G301) );
  NAND2_X1 U667 ( .A1(G868), .A2(G301), .ZN(n601) );
  NAND2_X1 U668 ( .A1(n637), .A2(G92), .ZN(n594) );
  NAND2_X1 U669 ( .A1(G79), .A2(n638), .ZN(n593) );
  NAND2_X1 U670 ( .A1(n594), .A2(n593), .ZN(n598) );
  NAND2_X1 U671 ( .A1(G54), .A2(n647), .ZN(n596) );
  NAND2_X1 U672 ( .A1(G66), .A2(n655), .ZN(n595) );
  NAND2_X1 U673 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U674 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U675 ( .A(KEYINPUT15), .B(n599), .ZN(n1000) );
  INV_X1 U676 ( .A(G868), .ZN(n668) );
  NAND2_X1 U677 ( .A1(n1000), .A2(n668), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n601), .A2(n600), .ZN(G284) );
  NAND2_X1 U679 ( .A1(n647), .A2(G53), .ZN(n603) );
  NAND2_X1 U680 ( .A1(G78), .A2(n638), .ZN(n602) );
  NAND2_X1 U681 ( .A1(n603), .A2(n602), .ZN(n606) );
  NAND2_X1 U682 ( .A1(G91), .A2(n637), .ZN(n604) );
  XNOR2_X1 U683 ( .A(KEYINPUT71), .B(n604), .ZN(n605) );
  NOR2_X1 U684 ( .A1(n606), .A2(n605), .ZN(n608) );
  NAND2_X1 U685 ( .A1(G65), .A2(n655), .ZN(n607) );
  NAND2_X1 U686 ( .A1(n608), .A2(n607), .ZN(G299) );
  XOR2_X1 U687 ( .A(KEYINPUT75), .B(n668), .Z(n609) );
  NOR2_X1 U688 ( .A1(G286), .A2(n609), .ZN(n612) );
  NOR2_X1 U689 ( .A1(G868), .A2(G299), .ZN(n610) );
  XNOR2_X1 U690 ( .A(n610), .B(KEYINPUT76), .ZN(n611) );
  NOR2_X1 U691 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U692 ( .A(KEYINPUT77), .B(n613), .Z(G297) );
  INV_X1 U693 ( .A(G559), .ZN(n617) );
  NOR2_X1 U694 ( .A1(G860), .A2(n617), .ZN(n614) );
  NOR2_X1 U695 ( .A1(n1000), .A2(n614), .ZN(n615) );
  XOR2_X1 U696 ( .A(n615), .B(KEYINPUT16), .Z(n616) );
  XNOR2_X1 U697 ( .A(KEYINPUT78), .B(n616), .ZN(G148) );
  INV_X1 U698 ( .A(n1000), .ZN(n697) );
  NAND2_X1 U699 ( .A1(n617), .A2(n697), .ZN(n618) );
  NAND2_X1 U700 ( .A1(n618), .A2(G868), .ZN(n620) );
  INV_X1 U701 ( .A(n999), .ZN(n694) );
  NAND2_X1 U702 ( .A1(n694), .A2(n668), .ZN(n619) );
  NAND2_X1 U703 ( .A1(n620), .A2(n619), .ZN(G282) );
  NAND2_X1 U704 ( .A1(n697), .A2(G559), .ZN(n665) );
  XOR2_X1 U705 ( .A(n999), .B(n665), .Z(n621) );
  NOR2_X1 U706 ( .A1(n621), .A2(G860), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n637), .A2(G93), .ZN(n623) );
  NAND2_X1 U708 ( .A1(G80), .A2(n638), .ZN(n622) );
  NAND2_X1 U709 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U710 ( .A1(G55), .A2(n647), .ZN(n625) );
  NAND2_X1 U711 ( .A1(G67), .A2(n655), .ZN(n624) );
  NAND2_X1 U712 ( .A1(n625), .A2(n624), .ZN(n626) );
  OR2_X1 U713 ( .A1(n627), .A2(n626), .ZN(n667) );
  XOR2_X1 U714 ( .A(n628), .B(n667), .Z(G145) );
  NAND2_X1 U715 ( .A1(G48), .A2(n647), .ZN(n630) );
  NAND2_X1 U716 ( .A1(G86), .A2(n637), .ZN(n629) );
  NAND2_X1 U717 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U718 ( .A1(n638), .A2(G73), .ZN(n631) );
  XNOR2_X1 U719 ( .A(n631), .B(KEYINPUT83), .ZN(n632) );
  XNOR2_X1 U720 ( .A(n632), .B(KEYINPUT2), .ZN(n633) );
  NOR2_X1 U721 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U722 ( .A1(G61), .A2(n655), .ZN(n635) );
  NAND2_X1 U723 ( .A1(n636), .A2(n635), .ZN(G305) );
  NAND2_X1 U724 ( .A1(n637), .A2(G85), .ZN(n640) );
  NAND2_X1 U725 ( .A1(G72), .A2(n638), .ZN(n639) );
  NAND2_X1 U726 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U727 ( .A(KEYINPUT69), .B(n641), .ZN(n645) );
  NAND2_X1 U728 ( .A1(n655), .A2(G60), .ZN(n643) );
  NAND2_X1 U729 ( .A1(G47), .A2(n647), .ZN(n642) );
  AND2_X1 U730 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U731 ( .A1(n645), .A2(n644), .ZN(G290) );
  NAND2_X1 U732 ( .A1(G651), .A2(G74), .ZN(n646) );
  XNOR2_X1 U733 ( .A(KEYINPUT80), .B(n646), .ZN(n650) );
  NAND2_X1 U734 ( .A1(n647), .A2(G49), .ZN(n648) );
  XOR2_X1 U735 ( .A(KEYINPUT79), .B(n648), .Z(n649) );
  NAND2_X1 U736 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U737 ( .A(KEYINPUT81), .B(n651), .ZN(n657) );
  NAND2_X1 U738 ( .A1(G87), .A2(n652), .ZN(n653) );
  XOR2_X1 U739 ( .A(KEYINPUT82), .B(n653), .Z(n654) );
  NOR2_X1 U740 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U741 ( .A1(n657), .A2(n656), .ZN(G288) );
  XNOR2_X1 U742 ( .A(KEYINPUT19), .B(KEYINPUT85), .ZN(n659) );
  XOR2_X1 U743 ( .A(G305), .B(G303), .Z(n658) );
  XNOR2_X1 U744 ( .A(n659), .B(n658), .ZN(n660) );
  XOR2_X1 U745 ( .A(n660), .B(n667), .Z(n662) );
  XOR2_X1 U746 ( .A(G290), .B(G299), .Z(n661) );
  XNOR2_X1 U747 ( .A(n662), .B(n661), .ZN(n663) );
  XOR2_X1 U748 ( .A(n663), .B(G288), .Z(n664) );
  XOR2_X1 U749 ( .A(n999), .B(n664), .Z(n918) );
  XNOR2_X1 U750 ( .A(n665), .B(n918), .ZN(n666) );
  NAND2_X1 U751 ( .A1(n666), .A2(G868), .ZN(n670) );
  NAND2_X1 U752 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U753 ( .A1(n670), .A2(n669), .ZN(G295) );
  NAND2_X1 U754 ( .A1(G2084), .A2(G2078), .ZN(n671) );
  XOR2_X1 U755 ( .A(KEYINPUT20), .B(n671), .Z(n672) );
  NAND2_X1 U756 ( .A1(G2090), .A2(n672), .ZN(n673) );
  XNOR2_X1 U757 ( .A(KEYINPUT21), .B(n673), .ZN(n674) );
  NAND2_X1 U758 ( .A1(n674), .A2(G2072), .ZN(G158) );
  NAND2_X1 U759 ( .A1(G661), .A2(G483), .ZN(n675) );
  XOR2_X1 U760 ( .A(KEYINPUT86), .B(n675), .Z(n676) );
  NAND2_X1 U761 ( .A1(n676), .A2(G319), .ZN(n677) );
  XNOR2_X1 U762 ( .A(n677), .B(KEYINPUT87), .ZN(n856) );
  NAND2_X1 U763 ( .A1(G36), .A2(n856), .ZN(n678) );
  XNOR2_X1 U764 ( .A(n678), .B(KEYINPUT88), .ZN(G176) );
  NAND2_X1 U765 ( .A1(G138), .A2(n898), .ZN(n680) );
  NAND2_X1 U766 ( .A1(G102), .A2(n899), .ZN(n679) );
  NAND2_X1 U767 ( .A1(n680), .A2(n679), .ZN(n684) );
  NAND2_X1 U768 ( .A1(G114), .A2(n894), .ZN(n682) );
  NAND2_X1 U769 ( .A1(G126), .A2(n895), .ZN(n681) );
  NAND2_X1 U770 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U771 ( .A1(n684), .A2(n683), .ZN(G164) );
  XNOR2_X1 U772 ( .A(KEYINPUT29), .B(KEYINPUT99), .ZN(n718) );
  NOR2_X1 U773 ( .A1(G164), .A2(G1384), .ZN(n762) );
  INV_X1 U774 ( .A(n762), .ZN(n699) );
  NAND2_X1 U775 ( .A1(G160), .A2(G40), .ZN(n761) );
  NAND2_X1 U776 ( .A1(G1996), .A2(n706), .ZN(n685) );
  XNOR2_X1 U777 ( .A(KEYINPUT26), .B(n685), .ZN(n687) );
  INV_X1 U778 ( .A(G1341), .ZN(n998) );
  NOR2_X1 U779 ( .A1(n706), .A2(n998), .ZN(n686) );
  NAND2_X1 U780 ( .A1(KEYINPUT26), .A2(n686), .ZN(n690) );
  NAND2_X1 U781 ( .A1(n687), .A2(n690), .ZN(n689) );
  INV_X1 U782 ( .A(KEYINPUT97), .ZN(n688) );
  NAND2_X1 U783 ( .A1(n689), .A2(n688), .ZN(n692) );
  NAND2_X1 U784 ( .A1(n690), .A2(KEYINPUT97), .ZN(n691) );
  NAND2_X1 U785 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U786 ( .A1(n694), .A2(n693), .ZN(n698) );
  NOR2_X1 U787 ( .A1(n698), .A2(n697), .ZN(n696) );
  INV_X1 U788 ( .A(KEYINPUT98), .ZN(n695) );
  XNOR2_X1 U789 ( .A(n696), .B(n695), .ZN(n705) );
  NAND2_X1 U790 ( .A1(n698), .A2(n697), .ZN(n703) );
  NOR2_X1 U791 ( .A1(n706), .A2(G1348), .ZN(n701) );
  NOR2_X1 U792 ( .A1(G2067), .A2(n738), .ZN(n700) );
  NOR2_X1 U793 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U794 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U795 ( .A1(n705), .A2(n704), .ZN(n711) );
  INV_X1 U796 ( .A(G299), .ZN(n713) );
  NAND2_X1 U797 ( .A1(n706), .A2(G2072), .ZN(n707) );
  XNOR2_X1 U798 ( .A(n707), .B(KEYINPUT27), .ZN(n709) );
  AND2_X1 U799 ( .A1(G1956), .A2(n738), .ZN(n708) );
  NOR2_X1 U800 ( .A1(n709), .A2(n708), .ZN(n712) );
  NAND2_X1 U801 ( .A1(n713), .A2(n712), .ZN(n710) );
  NAND2_X1 U802 ( .A1(n711), .A2(n710), .ZN(n716) );
  NOR2_X1 U803 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U804 ( .A(n714), .B(KEYINPUT28), .Z(n715) );
  NAND2_X1 U805 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U806 ( .A(n718), .B(n717), .ZN(n722) );
  XNOR2_X1 U807 ( .A(G2078), .B(KEYINPUT25), .ZN(n965) );
  NOR2_X1 U808 ( .A1(n738), .A2(n965), .ZN(n720) );
  AND2_X1 U809 ( .A1(n738), .A2(G1961), .ZN(n719) );
  NOR2_X1 U810 ( .A1(n720), .A2(n719), .ZN(n728) );
  NAND2_X1 U811 ( .A1(n728), .A2(G171), .ZN(n721) );
  NAND2_X1 U812 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U813 ( .A(n723), .B(KEYINPUT100), .ZN(n735) );
  NAND2_X1 U814 ( .A1(G8), .A2(n738), .ZN(n737) );
  NOR2_X1 U815 ( .A1(G2084), .A2(n738), .ZN(n757) );
  NOR2_X1 U816 ( .A1(n756), .A2(n757), .ZN(n724) );
  NAND2_X1 U817 ( .A1(G8), .A2(n724), .ZN(n725) );
  XNOR2_X1 U818 ( .A(KEYINPUT101), .B(n725), .ZN(n726) );
  XOR2_X1 U819 ( .A(KEYINPUT30), .B(n726), .Z(n727) );
  NOR2_X1 U820 ( .A1(G168), .A2(n727), .ZN(n730) );
  NOR2_X1 U821 ( .A1(G171), .A2(n728), .ZN(n729) );
  NOR2_X1 U822 ( .A1(n730), .A2(n729), .ZN(n733) );
  NAND2_X1 U823 ( .A1(n735), .A2(n734), .ZN(n754) );
  AND2_X1 U824 ( .A1(G286), .A2(G8), .ZN(n736) );
  NAND2_X1 U825 ( .A1(n754), .A2(n736), .ZN(n745) );
  INV_X1 U826 ( .A(G8), .ZN(n743) );
  INV_X1 U827 ( .A(n737), .ZN(n832) );
  NOR2_X1 U828 ( .A1(G1971), .A2(n737), .ZN(n740) );
  NOR2_X1 U829 ( .A1(G2090), .A2(n738), .ZN(n739) );
  NOR2_X1 U830 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U831 ( .A1(n741), .A2(G303), .ZN(n742) );
  OR2_X1 U832 ( .A1(n743), .A2(n742), .ZN(n744) );
  AND2_X1 U833 ( .A1(n745), .A2(n744), .ZN(n747) );
  INV_X1 U834 ( .A(KEYINPUT105), .ZN(n749) );
  NOR2_X1 U835 ( .A1(G1976), .A2(G288), .ZN(n1003) );
  NAND2_X1 U836 ( .A1(n1003), .A2(KEYINPUT33), .ZN(n748) );
  NAND2_X1 U837 ( .A1(n749), .A2(n748), .ZN(n751) );
  NAND2_X1 U838 ( .A1(n1003), .A2(KEYINPUT105), .ZN(n750) );
  NAND2_X1 U839 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U840 ( .A1(n737), .A2(n752), .ZN(n821) );
  INV_X1 U841 ( .A(n821), .ZN(n753) );
  AND2_X1 U842 ( .A1(n837), .A2(n753), .ZN(n797) );
  XNOR2_X1 U843 ( .A(KEYINPUT103), .B(n754), .ZN(n755) );
  NOR2_X1 U844 ( .A1(n756), .A2(n755), .ZN(n759) );
  NAND2_X1 U845 ( .A1(n757), .A2(G8), .ZN(n758) );
  NAND2_X1 U846 ( .A1(n759), .A2(n758), .ZN(n835) );
  NAND2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n992) );
  INV_X1 U848 ( .A(n992), .ZN(n760) );
  NOR2_X1 U849 ( .A1(n760), .A2(KEYINPUT105), .ZN(n813) );
  AND2_X1 U850 ( .A1(n835), .A2(n813), .ZN(n795) );
  XOR2_X1 U851 ( .A(G1981), .B(G305), .Z(n1009) );
  NOR2_X1 U852 ( .A1(n762), .A2(n761), .ZN(n845) );
  XNOR2_X1 U853 ( .A(KEYINPUT37), .B(G2067), .ZN(n798) );
  XNOR2_X1 U854 ( .A(KEYINPUT91), .B(KEYINPUT36), .ZN(n774) );
  NAND2_X1 U855 ( .A1(G116), .A2(n894), .ZN(n764) );
  NAND2_X1 U856 ( .A1(G128), .A2(n895), .ZN(n763) );
  NAND2_X1 U857 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U858 ( .A(KEYINPUT35), .B(n765), .ZN(n772) );
  XNOR2_X1 U859 ( .A(KEYINPUT34), .B(KEYINPUT90), .ZN(n770) );
  NAND2_X1 U860 ( .A1(G104), .A2(n899), .ZN(n768) );
  NAND2_X1 U861 ( .A1(G140), .A2(n898), .ZN(n766) );
  XOR2_X1 U862 ( .A(KEYINPUT89), .B(n766), .Z(n767) );
  NAND2_X1 U863 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U864 ( .A(n770), .B(n769), .Z(n771) );
  NAND2_X1 U865 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U866 ( .A(n774), .B(n773), .ZN(n914) );
  NOR2_X1 U867 ( .A1(n798), .A2(n914), .ZN(n948) );
  NAND2_X1 U868 ( .A1(n845), .A2(n948), .ZN(n808) );
  NAND2_X1 U869 ( .A1(G131), .A2(n898), .ZN(n775) );
  XNOR2_X1 U870 ( .A(n775), .B(KEYINPUT92), .ZN(n777) );
  NAND2_X1 U871 ( .A1(G95), .A2(n899), .ZN(n776) );
  NAND2_X1 U872 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U873 ( .A(KEYINPUT93), .B(n778), .ZN(n782) );
  NAND2_X1 U874 ( .A1(G107), .A2(n894), .ZN(n780) );
  NAND2_X1 U875 ( .A1(G119), .A2(n895), .ZN(n779) );
  AND2_X1 U876 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U877 ( .A1(n782), .A2(n781), .ZN(n909) );
  AND2_X1 U878 ( .A1(n909), .A2(G1991), .ZN(n793) );
  NAND2_X1 U879 ( .A1(G105), .A2(n899), .ZN(n783) );
  XNOR2_X1 U880 ( .A(KEYINPUT38), .B(n783), .ZN(n788) );
  NAND2_X1 U881 ( .A1(G117), .A2(n894), .ZN(n785) );
  NAND2_X1 U882 ( .A1(G129), .A2(n895), .ZN(n784) );
  NAND2_X1 U883 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U884 ( .A(KEYINPUT94), .B(n786), .Z(n787) );
  NAND2_X1 U885 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U886 ( .A(n789), .B(KEYINPUT95), .ZN(n791) );
  NAND2_X1 U887 ( .A1(G141), .A2(n898), .ZN(n790) );
  NAND2_X1 U888 ( .A1(n791), .A2(n790), .ZN(n911) );
  AND2_X1 U889 ( .A1(n911), .A2(G1996), .ZN(n792) );
  NOR2_X1 U890 ( .A1(n793), .A2(n792), .ZN(n946) );
  INV_X1 U891 ( .A(n946), .ZN(n794) );
  NAND2_X1 U892 ( .A1(n794), .A2(n845), .ZN(n800) );
  AND2_X1 U893 ( .A1(n808), .A2(n800), .ZN(n840) );
  AND2_X1 U894 ( .A1(n1009), .A2(n840), .ZN(n812) );
  AND2_X1 U895 ( .A1(n795), .A2(n812), .ZN(n796) );
  NAND2_X1 U896 ( .A1(n797), .A2(n796), .ZN(n826) );
  NAND2_X1 U897 ( .A1(n798), .A2(n914), .ZN(n959) );
  NOR2_X1 U898 ( .A1(n911), .A2(G1996), .ZN(n799) );
  XNOR2_X1 U899 ( .A(n799), .B(KEYINPUT106), .ZN(n939) );
  INV_X1 U900 ( .A(n800), .ZN(n804) );
  NOR2_X1 U901 ( .A1(G1991), .A2(n909), .ZN(n801) );
  XOR2_X1 U902 ( .A(KEYINPUT107), .B(n801), .Z(n944) );
  NOR2_X1 U903 ( .A1(G1986), .A2(G290), .ZN(n802) );
  NOR2_X1 U904 ( .A1(n944), .A2(n802), .ZN(n803) );
  NOR2_X1 U905 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U906 ( .A1(n939), .A2(n805), .ZN(n806) );
  XNOR2_X1 U907 ( .A(KEYINPUT108), .B(n806), .ZN(n807) );
  XNOR2_X1 U908 ( .A(n807), .B(KEYINPUT39), .ZN(n809) );
  NAND2_X1 U909 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U910 ( .A1(n959), .A2(n810), .ZN(n811) );
  NAND2_X1 U911 ( .A1(n811), .A2(n845), .ZN(n844) );
  INV_X1 U912 ( .A(n812), .ZN(n823) );
  INV_X1 U913 ( .A(KEYINPUT33), .ZN(n819) );
  INV_X1 U914 ( .A(n813), .ZN(n817) );
  NOR2_X1 U915 ( .A1(G303), .A2(G1971), .ZN(n814) );
  NOR2_X1 U916 ( .A1(n814), .A2(n1003), .ZN(n815) );
  OR2_X1 U917 ( .A1(n737), .A2(n815), .ZN(n816) );
  OR2_X1 U918 ( .A1(n817), .A2(n816), .ZN(n818) );
  AND2_X1 U919 ( .A1(n819), .A2(n818), .ZN(n820) );
  OR2_X1 U920 ( .A1(n821), .A2(n820), .ZN(n822) );
  OR2_X1 U921 ( .A1(n823), .A2(n822), .ZN(n824) );
  AND2_X1 U922 ( .A1(n844), .A2(n824), .ZN(n825) );
  AND2_X1 U923 ( .A1(n826), .A2(n825), .ZN(n843) );
  NOR2_X1 U924 ( .A1(G1981), .A2(G305), .ZN(n827) );
  XOR2_X1 U925 ( .A(n827), .B(KEYINPUT24), .Z(n828) );
  NOR2_X1 U926 ( .A1(n737), .A2(n828), .ZN(n829) );
  XOR2_X1 U927 ( .A(n829), .B(KEYINPUT96), .Z(n834) );
  NOR2_X1 U928 ( .A1(G2090), .A2(G303), .ZN(n830) );
  NAND2_X1 U929 ( .A1(G8), .A2(n830), .ZN(n831) );
  OR2_X1 U930 ( .A1(n832), .A2(n831), .ZN(n833) );
  AND2_X1 U931 ( .A1(n834), .A2(n833), .ZN(n839) );
  AND2_X1 U932 ( .A1(n835), .A2(n737), .ZN(n836) );
  NAND2_X1 U933 ( .A1(n837), .A2(n836), .ZN(n838) );
  NAND2_X1 U934 ( .A1(n839), .A2(n838), .ZN(n841) );
  NAND2_X1 U935 ( .A1(n841), .A2(n840), .ZN(n842) );
  NAND2_X1 U936 ( .A1(n843), .A2(n842), .ZN(n849) );
  INV_X1 U937 ( .A(n844), .ZN(n847) );
  XNOR2_X1 U938 ( .A(G1986), .B(G290), .ZN(n995) );
  NAND2_X1 U939 ( .A1(n995), .A2(n845), .ZN(n846) );
  OR2_X1 U940 ( .A1(n847), .A2(n846), .ZN(n848) );
  AND2_X1 U941 ( .A1(n849), .A2(n848), .ZN(n851) );
  XOR2_X1 U942 ( .A(KEYINPUT40), .B(KEYINPUT109), .Z(n850) );
  XNOR2_X1 U943 ( .A(n851), .B(n850), .ZN(G329) );
  NAND2_X1 U944 ( .A1(n853), .A2(G2106), .ZN(n852) );
  XNOR2_X1 U945 ( .A(n852), .B(KEYINPUT112), .ZN(G217) );
  INV_X1 U946 ( .A(n853), .ZN(G223) );
  AND2_X1 U947 ( .A1(G15), .A2(G2), .ZN(n854) );
  NAND2_X1 U948 ( .A1(G661), .A2(n854), .ZN(G259) );
  NAND2_X1 U949 ( .A1(G3), .A2(G1), .ZN(n855) );
  NAND2_X1 U950 ( .A1(n856), .A2(n855), .ZN(G188) );
  XNOR2_X1 U951 ( .A(G96), .B(KEYINPUT113), .ZN(G221) );
  INV_X1 U953 ( .A(G120), .ZN(G236) );
  INV_X1 U954 ( .A(G69), .ZN(G235) );
  NOR2_X1 U955 ( .A1(n858), .A2(n857), .ZN(G325) );
  INV_X1 U956 ( .A(G325), .ZN(G261) );
  XOR2_X1 U957 ( .A(G2100), .B(G2096), .Z(n860) );
  XNOR2_X1 U958 ( .A(KEYINPUT42), .B(G2678), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U960 ( .A(KEYINPUT43), .B(G2072), .Z(n862) );
  XNOR2_X1 U961 ( .A(G2067), .B(G2090), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U963 ( .A(n864), .B(n863), .Z(n866) );
  XNOR2_X1 U964 ( .A(G2084), .B(G2078), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n866), .B(n865), .ZN(G227) );
  XNOR2_X1 U966 ( .A(G1981), .B(G2474), .ZN(n876) );
  XOR2_X1 U967 ( .A(G1956), .B(G1961), .Z(n868) );
  XNOR2_X1 U968 ( .A(G1976), .B(G1966), .ZN(n867) );
  XNOR2_X1 U969 ( .A(n868), .B(n867), .ZN(n872) );
  XOR2_X1 U970 ( .A(G1971), .B(G1986), .Z(n870) );
  XNOR2_X1 U971 ( .A(G1996), .B(G1991), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n870), .B(n869), .ZN(n871) );
  XOR2_X1 U973 ( .A(n872), .B(n871), .Z(n874) );
  XNOR2_X1 U974 ( .A(KEYINPUT114), .B(KEYINPUT41), .ZN(n873) );
  XNOR2_X1 U975 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U976 ( .A(n876), .B(n875), .ZN(G229) );
  NAND2_X1 U977 ( .A1(G124), .A2(n895), .ZN(n877) );
  XNOR2_X1 U978 ( .A(n877), .B(KEYINPUT44), .ZN(n879) );
  NAND2_X1 U979 ( .A1(n894), .A2(G112), .ZN(n878) );
  NAND2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n883) );
  NAND2_X1 U981 ( .A1(G136), .A2(n898), .ZN(n881) );
  NAND2_X1 U982 ( .A1(G100), .A2(n899), .ZN(n880) );
  NAND2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n882) );
  NOR2_X1 U984 ( .A1(n883), .A2(n882), .ZN(G162) );
  XOR2_X1 U985 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n893) );
  NAND2_X1 U986 ( .A1(G139), .A2(n898), .ZN(n885) );
  NAND2_X1 U987 ( .A1(G103), .A2(n899), .ZN(n884) );
  NAND2_X1 U988 ( .A1(n885), .A2(n884), .ZN(n891) );
  NAND2_X1 U989 ( .A1(n895), .A2(G127), .ZN(n886) );
  XOR2_X1 U990 ( .A(KEYINPUT115), .B(n886), .Z(n888) );
  NAND2_X1 U991 ( .A1(n894), .A2(G115), .ZN(n887) );
  NAND2_X1 U992 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U993 ( .A(KEYINPUT47), .B(n889), .Z(n890) );
  NOR2_X1 U994 ( .A1(n891), .A2(n890), .ZN(n952) );
  XNOR2_X1 U995 ( .A(G164), .B(n952), .ZN(n892) );
  XNOR2_X1 U996 ( .A(n893), .B(n892), .ZN(n906) );
  NAND2_X1 U997 ( .A1(G118), .A2(n894), .ZN(n897) );
  NAND2_X1 U998 ( .A1(G130), .A2(n895), .ZN(n896) );
  NAND2_X1 U999 ( .A1(n897), .A2(n896), .ZN(n904) );
  NAND2_X1 U1000 ( .A1(G142), .A2(n898), .ZN(n901) );
  NAND2_X1 U1001 ( .A1(G106), .A2(n899), .ZN(n900) );
  NAND2_X1 U1002 ( .A1(n901), .A2(n900), .ZN(n902) );
  XOR2_X1 U1003 ( .A(n902), .B(KEYINPUT45), .Z(n903) );
  NOR2_X1 U1004 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U1005 ( .A(n906), .B(n905), .Z(n907) );
  XOR2_X1 U1006 ( .A(G162), .B(n907), .Z(n908) );
  XNOR2_X1 U1007 ( .A(n941), .B(n908), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(n910), .B(n909), .ZN(n913) );
  XOR2_X1 U1009 ( .A(G160), .B(n911), .Z(n912) );
  XNOR2_X1 U1010 ( .A(n913), .B(n912), .ZN(n915) );
  XOR2_X1 U1011 ( .A(n915), .B(n914), .Z(n916) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n916), .ZN(G395) );
  XNOR2_X1 U1013 ( .A(G171), .B(n1000), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(n918), .B(n917), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(n919), .B(G286), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n920), .ZN(G397) );
  XNOR2_X1 U1017 ( .A(G2427), .B(KEYINPUT111), .ZN(n930) );
  XOR2_X1 U1018 ( .A(G2443), .B(G2438), .Z(n922) );
  XNOR2_X1 U1019 ( .A(G2430), .B(G2454), .ZN(n921) );
  XNOR2_X1 U1020 ( .A(n922), .B(n921), .ZN(n926) );
  XOR2_X1 U1021 ( .A(KEYINPUT110), .B(G2435), .Z(n924) );
  XOR2_X1 U1022 ( .A(G1348), .B(n998), .Z(n923) );
  XNOR2_X1 U1023 ( .A(n924), .B(n923), .ZN(n925) );
  XOR2_X1 U1024 ( .A(n926), .B(n925), .Z(n928) );
  XNOR2_X1 U1025 ( .A(G2451), .B(G2446), .ZN(n927) );
  XNOR2_X1 U1026 ( .A(n928), .B(n927), .ZN(n929) );
  XNOR2_X1 U1027 ( .A(n930), .B(n929), .ZN(n931) );
  NAND2_X1 U1028 ( .A1(n931), .A2(G14), .ZN(n937) );
  NAND2_X1 U1029 ( .A1(G319), .A2(n937), .ZN(n934) );
  NOR2_X1 U1030 ( .A1(G227), .A2(G229), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(KEYINPUT49), .B(n932), .ZN(n933) );
  NOR2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n936) );
  NOR2_X1 U1033 ( .A1(G395), .A2(G397), .ZN(n935) );
  NAND2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(G225) );
  INV_X1 U1035 ( .A(G225), .ZN(G308) );
  INV_X1 U1036 ( .A(G108), .ZN(G238) );
  INV_X1 U1037 ( .A(n937), .ZN(G401) );
  XNOR2_X1 U1038 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n1047) );
  XOR2_X1 U1039 ( .A(G2090), .B(G162), .Z(n938) );
  NOR2_X1 U1040 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1041 ( .A(KEYINPUT51), .B(n940), .Z(n951) );
  XNOR2_X1 U1042 ( .A(G160), .B(G2084), .ZN(n942) );
  NAND2_X1 U1043 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1044 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1047 ( .A(n949), .B(KEYINPUT116), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n957) );
  XOR2_X1 U1049 ( .A(G2072), .B(n952), .Z(n954) );
  XOR2_X1 U1050 ( .A(G164), .B(G2078), .Z(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1052 ( .A(KEYINPUT50), .B(n955), .Z(n956) );
  NOR2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(n960), .B(KEYINPUT52), .ZN(n961) );
  XNOR2_X1 U1056 ( .A(KEYINPUT117), .B(n961), .ZN(n962) );
  INV_X1 U1057 ( .A(KEYINPUT55), .ZN(n985) );
  NAND2_X1 U1058 ( .A1(n962), .A2(n985), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n963), .A2(G29), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(KEYINPUT118), .B(n964), .ZN(n1045) );
  XOR2_X1 U1061 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n977) );
  XNOR2_X1 U1062 ( .A(G27), .B(n965), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(G1996), .B(G32), .ZN(n967) );
  XNOR2_X1 U1064 ( .A(G2072), .B(G33), .ZN(n966) );
  NOR2_X1 U1065 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n971) );
  XNOR2_X1 U1067 ( .A(G26), .B(G2067), .ZN(n970) );
  NOR2_X1 U1068 ( .A1(n971), .A2(n970), .ZN(n975) );
  XOR2_X1 U1069 ( .A(G1991), .B(G25), .Z(n972) );
  NAND2_X1 U1070 ( .A1(n972), .A2(G28), .ZN(n973) );
  XNOR2_X1 U1071 ( .A(n973), .B(KEYINPUT119), .ZN(n974) );
  NAND2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1073 ( .A(n977), .B(n976), .ZN(n983) );
  XOR2_X1 U1074 ( .A(G2090), .B(G35), .Z(n981) );
  XNOR2_X1 U1075 ( .A(KEYINPUT54), .B(G34), .ZN(n978) );
  XNOR2_X1 U1076 ( .A(n978), .B(KEYINPUT121), .ZN(n979) );
  XNOR2_X1 U1077 ( .A(n979), .B(G2084), .ZN(n980) );
  NAND2_X1 U1078 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1079 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1080 ( .A(n985), .B(n984), .Z(n987) );
  INV_X1 U1081 ( .A(G29), .ZN(n986) );
  NAND2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1083 ( .A1(n988), .A2(G11), .ZN(n1043) );
  INV_X1 U1084 ( .A(G16), .ZN(n1039) );
  XOR2_X1 U1085 ( .A(n1039), .B(KEYINPUT56), .Z(n1015) );
  XOR2_X1 U1086 ( .A(G303), .B(G1971), .Z(n989) );
  XNOR2_X1 U1087 ( .A(n989), .B(KEYINPUT123), .ZN(n991) );
  XOR2_X1 U1088 ( .A(G171), .B(G1961), .Z(n990) );
  NOR2_X1 U1089 ( .A1(n991), .A2(n990), .ZN(n997) );
  XOR2_X1 U1090 ( .A(G1956), .B(G299), .Z(n993) );
  NAND2_X1 U1091 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1092 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1093 ( .A1(n997), .A2(n996), .ZN(n1007) );
  XOR2_X1 U1094 ( .A(n999), .B(n998), .Z(n1005) );
  XNOR2_X1 U1095 ( .A(G1348), .B(n1000), .ZN(n1001) );
  XNOR2_X1 U1096 ( .A(KEYINPUT122), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1097 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1098 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1099 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1100 ( .A(KEYINPUT124), .B(n1008), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(G168), .B(G1966), .ZN(n1010) );
  NAND2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1103 ( .A(KEYINPUT57), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1041) );
  XNOR2_X1 U1106 ( .A(G1986), .B(G24), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(G1976), .B(G23), .ZN(n1017) );
  XNOR2_X1 U1108 ( .A(G22), .B(G1971), .ZN(n1016) );
  NOR2_X1 U1109 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1110 ( .A(KEYINPUT125), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1111 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1112 ( .A(KEYINPUT58), .B(n1021), .ZN(n1022) );
  XNOR2_X1 U1113 ( .A(n1022), .B(KEYINPUT126), .ZN(n1034) );
  XOR2_X1 U1114 ( .A(G19), .B(G1341), .Z(n1026) );
  XNOR2_X1 U1115 ( .A(G1981), .B(G6), .ZN(n1024) );
  XNOR2_X1 U1116 ( .A(G1956), .B(G20), .ZN(n1023) );
  NOR2_X1 U1117 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1118 ( .A1(n1026), .A2(n1025), .ZN(n1029) );
  XOR2_X1 U1119 ( .A(KEYINPUT59), .B(G1348), .Z(n1027) );
  XNOR2_X1 U1120 ( .A(G4), .B(n1027), .ZN(n1028) );
  NOR2_X1 U1121 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1122 ( .A(KEYINPUT60), .B(n1030), .Z(n1032) );
  XNOR2_X1 U1123 ( .A(G1966), .B(G21), .ZN(n1031) );
  NOR2_X1 U1124 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1125 ( .A1(n1034), .A2(n1033), .ZN(n1036) );
  XNOR2_X1 U1126 ( .A(G5), .B(G1961), .ZN(n1035) );
  NOR2_X1 U1127 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XNOR2_X1 U1128 ( .A(KEYINPUT61), .B(n1037), .ZN(n1038) );
  NAND2_X1 U1129 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NAND2_X1 U1130 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  NOR2_X1 U1131 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  NAND2_X1 U1132 ( .A1(n1045), .A2(n1044), .ZN(n1046) );
  XOR2_X1 U1133 ( .A(n1047), .B(n1046), .Z(G150) );
  INV_X1 U1134 ( .A(G150), .ZN(G311) );
endmodule

