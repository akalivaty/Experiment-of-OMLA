

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757;

  INV_X1 U374 ( .A(KEYINPUT85), .ZN(n353) );
  AND2_X1 U375 ( .A1(n369), .A2(n368), .ZN(n367) );
  XNOR2_X1 U376 ( .A(KEYINPUT32), .B(n579), .ZN(n755) );
  AND2_X1 U377 ( .A1(n593), .A2(KEYINPUT34), .ZN(n381) );
  BUF_X1 U378 ( .A(G113), .Z(n352) );
  XNOR2_X1 U379 ( .A(KEYINPUT3), .B(G113), .ZN(n454) );
  AND2_X2 U380 ( .A1(n362), .A2(n361), .ZN(n371) );
  XNOR2_X2 U381 ( .A(n461), .B(n460), .ZN(n523) );
  XNOR2_X2 U382 ( .A(n607), .B(n353), .ZN(n648) );
  XNOR2_X1 U383 ( .A(n559), .B(n558), .ZN(n609) );
  INV_X1 U384 ( .A(G953), .ZN(n745) );
  XNOR2_X2 U385 ( .A(n449), .B(KEYINPUT4), .ZN(n465) );
  INV_X1 U386 ( .A(n586), .ZN(n631) );
  NOR2_X1 U387 ( .A1(n542), .A2(n631), .ZN(n513) );
  INV_X1 U388 ( .A(KEYINPUT70), .ZN(n408) );
  AND2_X2 U389 ( .A1(n659), .A2(n658), .ZN(n720) );
  NOR2_X1 U390 ( .A1(n383), .A2(n381), .ZN(n421) );
  NOR2_X2 U391 ( .A1(n526), .A2(n525), .ZN(n698) );
  NOR2_X1 U392 ( .A1(n575), .A2(n587), .ZN(n583) );
  XNOR2_X1 U393 ( .A(n516), .B(KEYINPUT104), .ZN(n526) );
  XNOR2_X1 U394 ( .A(n590), .B(n404), .ZN(n593) );
  INV_X1 U395 ( .A(n585), .ZN(n625) );
  XNOR2_X1 U396 ( .A(n472), .B(G469), .ZN(n540) );
  XNOR2_X1 U397 ( .A(n418), .B(n484), .ZN(n585) );
  XNOR2_X1 U398 ( .A(n454), .B(n408), .ZN(n407) );
  XNOR2_X1 U399 ( .A(G119), .B(G116), .ZN(n406) );
  NAND2_X2 U400 ( .A1(n580), .A2(n755), .ZN(n581) );
  XNOR2_X1 U401 ( .A(n465), .B(n464), .ZN(n487) );
  AND2_X1 U402 ( .A1(n548), .A2(n414), .ZN(n413) );
  XNOR2_X1 U403 ( .A(n530), .B(n415), .ZN(n414) );
  OR2_X1 U404 ( .A1(G902), .A2(G237), .ZN(n496) );
  XNOR2_X1 U405 ( .A(n465), .B(n451), .ZN(n360) );
  INV_X1 U406 ( .A(n450), .ZN(n451) );
  XNOR2_X1 U407 ( .A(n390), .B(n389), .ZN(n541) );
  INV_X1 U408 ( .A(G472), .ZN(n389) );
  OR2_X1 U409 ( .A1(n677), .A2(G902), .ZN(n390) );
  NOR2_X1 U410 ( .A1(n411), .A2(n409), .ZN(n549) );
  XNOR2_X1 U411 ( .A(n410), .B(KEYINPUT46), .ZN(n409) );
  XNOR2_X1 U412 ( .A(n528), .B(KEYINPUT73), .ZN(n412) );
  NAND2_X1 U413 ( .A1(n377), .A2(KEYINPUT87), .ZN(n361) );
  NAND2_X1 U414 ( .A1(n374), .A2(n373), .ZN(n372) );
  NAND2_X1 U415 ( .A1(n367), .A2(n363), .ZN(n375) );
  NAND2_X1 U416 ( .A1(n366), .A2(n364), .ZN(n363) );
  NAND2_X1 U417 ( .A1(n370), .A2(KEYINPUT44), .ZN(n368) );
  AND2_X1 U418 ( .A1(n611), .A2(n497), .ZN(n401) );
  INV_X1 U419 ( .A(n509), .ZN(n403) );
  XNOR2_X1 U420 ( .A(n417), .B(G125), .ZN(n450) );
  INV_X1 U421 ( .A(G146), .ZN(n417) );
  NAND2_X1 U422 ( .A1(n670), .A2(n652), .ZN(n461) );
  XNOR2_X1 U423 ( .A(n391), .B(n495), .ZN(n677) );
  XNOR2_X1 U424 ( .A(n487), .B(n488), .ZN(n391) );
  XNOR2_X1 U425 ( .A(n450), .B(n416), .ZN(n742) );
  INV_X1 U426 ( .A(KEYINPUT10), .ZN(n416) );
  XNOR2_X1 U427 ( .A(G128), .B(G110), .ZN(n473) );
  XOR2_X1 U428 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n474) );
  XNOR2_X1 U429 ( .A(n384), .B(n428), .ZN(n430) );
  XNOR2_X1 U430 ( .A(G116), .B(G122), .ZN(n428) );
  XNOR2_X1 U431 ( .A(n385), .B(KEYINPUT9), .ZN(n384) );
  XNOR2_X1 U432 ( .A(KEYINPUT98), .B(KEYINPUT7), .ZN(n385) );
  INV_X1 U433 ( .A(G143), .ZN(n425) );
  XNOR2_X1 U434 ( .A(n476), .B(KEYINPUT93), .ZN(n466) );
  NOR2_X1 U435 ( .A1(n542), .A2(n582), .ZN(n543) );
  NAND2_X1 U436 ( .A1(n422), .A2(n566), .ZN(n383) );
  NOR2_X1 U437 ( .A1(n609), .A2(KEYINPUT34), .ZN(n423) );
  XNOR2_X1 U438 ( .A(n387), .B(n386), .ZN(n533) );
  INV_X1 U439 ( .A(G478), .ZN(n386) );
  OR2_X1 U440 ( .A1(n717), .A2(G902), .ZN(n387) );
  INV_X1 U441 ( .A(KEYINPUT92), .ZN(n404) );
  OR2_X1 U442 ( .A1(n721), .A2(G902), .ZN(n418) );
  NAND2_X1 U443 ( .A1(n656), .A2(n655), .ZN(n659) );
  XOR2_X1 U444 ( .A(KEYINPUT89), .B(n665), .Z(n719) );
  INV_X1 U445 ( .A(KEYINPUT83), .ZN(n415) );
  NOR2_X1 U446 ( .A1(KEYINPUT47), .A2(n527), .ZN(n528) );
  NAND2_X1 U447 ( .A1(n388), .A2(n757), .ZN(n410) );
  NAND2_X1 U448 ( .A1(n599), .A2(n598), .ZN(n377) );
  INV_X1 U449 ( .A(KEYINPUT71), .ZN(n370) );
  AND2_X1 U450 ( .A1(n365), .A2(KEYINPUT71), .ZN(n364) );
  INV_X1 U451 ( .A(KEYINPUT44), .ZN(n365) );
  XOR2_X1 U452 ( .A(G146), .B(G137), .Z(n491) );
  XNOR2_X1 U453 ( .A(G140), .B(G143), .ZN(n438) );
  XNOR2_X1 U454 ( .A(n352), .B(G122), .ZN(n440) );
  NOR2_X1 U455 ( .A1(G953), .A2(G237), .ZN(n489) );
  AND2_X1 U456 ( .A1(n754), .A2(n393), .ZN(n392) );
  INV_X1 U457 ( .A(n710), .ZN(n393) );
  XNOR2_X1 U458 ( .A(n395), .B(n405), .ZN(n602) );
  INV_X1 U459 ( .A(KEYINPUT45), .ZN(n405) );
  NAND2_X1 U460 ( .A1(n372), .A2(n371), .ZN(n376) );
  XNOR2_X1 U461 ( .A(G131), .B(G134), .ZN(n464) );
  XOR2_X1 U462 ( .A(KEYINPUT14), .B(KEYINPUT91), .Z(n499) );
  XNOR2_X1 U463 ( .A(n555), .B(n463), .ZN(n610) );
  XNOR2_X1 U464 ( .A(n462), .B(KEYINPUT38), .ZN(n463) );
  NOR2_X1 U465 ( .A1(n403), .A2(n355), .ZN(n399) );
  XNOR2_X1 U466 ( .A(n359), .B(n378), .ZN(n670) );
  XNOR2_X1 U467 ( .A(n726), .B(n360), .ZN(n359) );
  XNOR2_X1 U468 ( .A(n572), .B(n573), .ZN(n575) );
  BUF_X1 U469 ( .A(n523), .Z(n555) );
  XNOR2_X1 U470 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U471 ( .A(n477), .B(n419), .ZN(n721) );
  XNOR2_X1 U472 ( .A(n478), .B(n356), .ZN(n419) );
  XNOR2_X1 U473 ( .A(n435), .B(n434), .ZN(n717) );
  XNOR2_X1 U474 ( .A(n662), .B(n661), .ZN(n663) );
  AND2_X1 U475 ( .A1(n380), .A2(n379), .ZN(n707) );
  INV_X1 U476 ( .A(n621), .ZN(n379) );
  XNOR2_X1 U477 ( .A(n546), .B(KEYINPUT36), .ZN(n380) );
  NAND2_X1 U478 ( .A1(n424), .A2(n423), .ZN(n420) );
  XNOR2_X1 U479 ( .A(n711), .B(n712), .ZN(n713) );
  XOR2_X1 U480 ( .A(G110), .B(G104), .Z(n354) );
  NOR2_X1 U481 ( .A1(n611), .A2(n497), .ZN(n355) );
  AND2_X1 U482 ( .A1(n479), .A2(G221), .ZN(n356) );
  XNOR2_X1 U483 ( .A(n487), .B(n466), .ZN(n741) );
  XNOR2_X1 U484 ( .A(KEYINPUT86), .B(KEYINPUT48), .ZN(n357) );
  AND2_X1 U485 ( .A1(KEYINPUT87), .A2(KEYINPUT44), .ZN(n358) );
  XNOR2_X2 U486 ( .A(n494), .B(n456), .ZN(n726) );
  NAND2_X1 U487 ( .A1(n581), .A2(n358), .ZN(n362) );
  INV_X1 U488 ( .A(n581), .ZN(n366) );
  NAND2_X1 U489 ( .A1(n581), .A2(n370), .ZN(n369) );
  NAND2_X1 U490 ( .A1(n581), .A2(KEYINPUT44), .ZN(n373) );
  NOR2_X1 U491 ( .A1(n377), .A2(KEYINPUT87), .ZN(n374) );
  NAND2_X1 U492 ( .A1(n376), .A2(n375), .ZN(n395) );
  XNOR2_X1 U493 ( .A(n470), .B(n457), .ZN(n378) );
  NAND2_X1 U494 ( .A1(n413), .A2(n412), .ZN(n411) );
  XNOR2_X1 U495 ( .A(n549), .B(n357), .ZN(n394) );
  NAND2_X1 U496 ( .A1(n720), .A2(G475), .ZN(n664) );
  NOR2_X2 U497 ( .A1(n625), .A2(n574), .ZN(n691) );
  NAND2_X1 U498 ( .A1(n657), .A2(n653), .ZN(n656) );
  NOR2_X2 U499 ( .A1(n602), .A2(n601), .ZN(n657) );
  NAND2_X1 U500 ( .A1(n720), .A2(G217), .ZN(n723) );
  XNOR2_X1 U501 ( .A(n382), .B(KEYINPUT123), .ZN(G66) );
  NAND2_X1 U502 ( .A1(n725), .A2(n724), .ZN(n382) );
  NAND2_X1 U503 ( .A1(n557), .A2(n587), .ZN(n559) );
  INV_X1 U504 ( .A(n533), .ZN(n517) );
  XNOR2_X1 U505 ( .A(n388), .B(G131), .ZN(G33) );
  XNOR2_X2 U506 ( .A(n522), .B(KEYINPUT40), .ZN(n388) );
  NAND2_X1 U507 ( .A1(n394), .A2(n392), .ZN(n601) );
  NAND2_X1 U508 ( .A1(n586), .A2(n401), .ZN(n400) );
  AND2_X1 U509 ( .A1(n397), .A2(n396), .ZN(n505) );
  INV_X1 U510 ( .A(n594), .ZN(n396) );
  NOR2_X1 U511 ( .A1(n402), .A2(n398), .ZN(n397) );
  NAND2_X1 U512 ( .A1(n400), .A2(n399), .ZN(n398) );
  NOR2_X1 U513 ( .A1(n586), .A2(n497), .ZN(n402) );
  XNOR2_X2 U514 ( .A(n565), .B(KEYINPUT0), .ZN(n590) );
  XNOR2_X2 U515 ( .A(n407), .B(n406), .ZN(n494) );
  NAND2_X1 U516 ( .A1(n421), .A2(n420), .ZN(n567) );
  INV_X1 U517 ( .A(n593), .ZN(n424) );
  NAND2_X1 U518 ( .A1(n609), .A2(KEYINPUT34), .ZN(n422) );
  XNOR2_X2 U519 ( .A(n426), .B(n425), .ZN(n449) );
  XNOR2_X2 U520 ( .A(G128), .B(KEYINPUT79), .ZN(n426) );
  XNOR2_X1 U521 ( .A(n545), .B(n524), .ZN(n564) );
  XNOR2_X1 U522 ( .A(n664), .B(n663), .ZN(n666) );
  XNOR2_X1 U523 ( .A(n723), .B(n722), .ZN(n725) );
  BUF_X1 U524 ( .A(n564), .Z(n525) );
  NOR2_X2 U525 ( .A1(n564), .A2(n563), .ZN(n565) );
  INV_X1 U526 ( .A(n721), .ZN(n722) );
  AND2_X1 U527 ( .A1(n745), .A2(n647), .ZN(n427) );
  INV_X1 U528 ( .A(KEYINPUT74), .ZN(n462) );
  XNOR2_X1 U529 ( .A(n455), .B(G122), .ZN(n456) );
  NOR2_X1 U530 ( .A1(n657), .A2(n604), .ZN(n600) );
  XNOR2_X1 U531 ( .A(n494), .B(n493), .ZN(n495) );
  INV_X1 U532 ( .A(n540), .ZN(n514) );
  INV_X1 U533 ( .A(KEYINPUT1), .ZN(n539) );
  BUF_X1 U534 ( .A(n602), .Z(n732) );
  XNOR2_X1 U535 ( .A(n741), .B(n471), .ZN(n711) );
  XNOR2_X1 U536 ( .A(n540), .B(n539), .ZN(n587) );
  INV_X1 U537 ( .A(KEYINPUT39), .ZN(n507) );
  XNOR2_X1 U538 ( .A(n679), .B(n678), .ZN(n680) );
  INV_X1 U539 ( .A(KEYINPUT120), .ZN(n649) );
  XNOR2_X1 U540 ( .A(n714), .B(n713), .ZN(n715) );
  XNOR2_X1 U541 ( .A(G107), .B(G134), .ZN(n429) );
  XNOR2_X1 U542 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U543 ( .A(n449), .B(n431), .ZN(n435) );
  NAND2_X1 U544 ( .A1(n745), .A2(G234), .ZN(n433) );
  XNOR2_X1 U545 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n432) );
  XNOR2_X1 U546 ( .A(n433), .B(n432), .ZN(n479) );
  NAND2_X1 U547 ( .A1(G217), .A2(n479), .ZN(n434) );
  XOR2_X1 U548 ( .A(KEYINPUT97), .B(KEYINPUT13), .Z(n437) );
  XNOR2_X1 U549 ( .A(KEYINPUT96), .B(G475), .ZN(n436) );
  XNOR2_X1 U550 ( .A(n437), .B(n436), .ZN(n448) );
  XOR2_X1 U551 ( .A(G131), .B(G104), .Z(n439) );
  XNOR2_X1 U552 ( .A(n439), .B(n438), .ZN(n443) );
  XOR2_X1 U553 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n441) );
  XNOR2_X1 U554 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U555 ( .A(n443), .B(n442), .Z(n445) );
  NAND2_X1 U556 ( .A1(n489), .A2(G214), .ZN(n444) );
  XNOR2_X1 U557 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U558 ( .A(n742), .B(n446), .ZN(n660) );
  NOR2_X1 U559 ( .A1(G902), .A2(n660), .ZN(n447) );
  XNOR2_X1 U560 ( .A(n448), .B(n447), .ZN(n531) );
  NOR2_X1 U561 ( .A1(n533), .A2(n531), .ZN(n692) );
  XOR2_X1 U562 ( .A(KEYINPUT66), .B(G101), .Z(n488) );
  XNOR2_X1 U563 ( .A(G107), .B(n354), .ZN(n727) );
  XNOR2_X1 U564 ( .A(n488), .B(n727), .ZN(n470) );
  XOR2_X1 U565 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n453) );
  NAND2_X1 U566 ( .A1(G224), .A2(n745), .ZN(n452) );
  XNOR2_X1 U567 ( .A(n453), .B(n452), .ZN(n457) );
  INV_X1 U568 ( .A(KEYINPUT16), .ZN(n455) );
  XNOR2_X1 U569 ( .A(G902), .B(KEYINPUT15), .ZN(n652) );
  XOR2_X1 U570 ( .A(KEYINPUT80), .B(KEYINPUT90), .Z(n459) );
  NAND2_X1 U571 ( .A1(G210), .A2(n496), .ZN(n458) );
  XNOR2_X1 U572 ( .A(n459), .B(n458), .ZN(n460) );
  INV_X1 U573 ( .A(n610), .ZN(n506) );
  XOR2_X1 U574 ( .A(G137), .B(G140), .Z(n476) );
  XOR2_X1 U575 ( .A(G146), .B(KEYINPUT78), .Z(n468) );
  NAND2_X1 U576 ( .A1(G227), .A2(n745), .ZN(n467) );
  XNOR2_X1 U577 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U578 ( .A(n470), .B(n469), .ZN(n471) );
  NOR2_X1 U579 ( .A1(n711), .A2(G902), .ZN(n472) );
  XNOR2_X1 U580 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U581 ( .A(n475), .B(G119), .Z(n478) );
  XNOR2_X1 U582 ( .A(n742), .B(n476), .ZN(n477) );
  XOR2_X1 U583 ( .A(KEYINPUT25), .B(KEYINPUT77), .Z(n483) );
  NAND2_X1 U584 ( .A1(n652), .A2(G234), .ZN(n480) );
  XNOR2_X1 U585 ( .A(n480), .B(KEYINPUT20), .ZN(n481) );
  XNOR2_X1 U586 ( .A(KEYINPUT94), .B(n481), .ZN(n485) );
  NAND2_X1 U587 ( .A1(G217), .A2(n485), .ZN(n482) );
  XNOR2_X1 U588 ( .A(n483), .B(n482), .ZN(n484) );
  NAND2_X1 U589 ( .A1(n485), .A2(G221), .ZN(n486) );
  XOR2_X1 U590 ( .A(n486), .B(KEYINPUT21), .Z(n626) );
  XOR2_X1 U591 ( .A(n626), .B(KEYINPUT95), .Z(n568) );
  NAND2_X1 U592 ( .A1(n625), .A2(n568), .ZN(n622) );
  OR2_X1 U593 ( .A1(n540), .A2(n622), .ZN(n594) );
  INV_X1 U594 ( .A(KEYINPUT30), .ZN(n497) );
  NAND2_X1 U595 ( .A1(n489), .A2(G210), .ZN(n490) );
  XNOR2_X1 U596 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U597 ( .A(n492), .B(KEYINPUT5), .Z(n493) );
  INV_X1 U598 ( .A(n541), .ZN(n586) );
  NAND2_X1 U599 ( .A1(G214), .A2(n496), .ZN(n611) );
  NAND2_X1 U600 ( .A1(G237), .A2(G234), .ZN(n498) );
  XNOR2_X1 U601 ( .A(n499), .B(n498), .ZN(n501) );
  NAND2_X1 U602 ( .A1(G952), .A2(n501), .ZN(n643) );
  NOR2_X1 U603 ( .A1(G953), .A2(n643), .ZN(n562) );
  AND2_X1 U604 ( .A1(G953), .A2(G902), .ZN(n500) );
  NAND2_X1 U605 ( .A1(n501), .A2(n500), .ZN(n560) );
  XOR2_X1 U606 ( .A(n560), .B(KEYINPUT101), .Z(n502) );
  NOR2_X1 U607 ( .A1(G900), .A2(n502), .ZN(n503) );
  NOR2_X1 U608 ( .A1(n562), .A2(n503), .ZN(n504) );
  XNOR2_X1 U609 ( .A(KEYINPUT81), .B(n504), .ZN(n509) );
  XNOR2_X1 U610 ( .A(n505), .B(KEYINPUT75), .ZN(n535) );
  NOR2_X1 U611 ( .A1(n506), .A2(n535), .ZN(n508) );
  XNOR2_X1 U612 ( .A(n508), .B(n507), .ZN(n521) );
  AND2_X1 U613 ( .A1(n692), .A2(n521), .ZN(n710) );
  NAND2_X1 U614 ( .A1(n626), .A2(n509), .ZN(n510) );
  XNOR2_X1 U615 ( .A(KEYINPUT69), .B(n510), .ZN(n511) );
  NAND2_X1 U616 ( .A1(n511), .A2(n585), .ZN(n512) );
  XNOR2_X1 U617 ( .A(KEYINPUT68), .B(n512), .ZN(n542) );
  XNOR2_X1 U618 ( .A(n513), .B(KEYINPUT28), .ZN(n515) );
  NAND2_X1 U619 ( .A1(n515), .A2(n514), .ZN(n516) );
  NAND2_X1 U620 ( .A1(n611), .A2(n610), .ZN(n616) );
  NOR2_X1 U621 ( .A1(n531), .A2(n517), .ZN(n569) );
  INV_X1 U622 ( .A(n569), .ZN(n613) );
  NOR2_X1 U623 ( .A1(n616), .A2(n613), .ZN(n518) );
  XNOR2_X1 U624 ( .A(KEYINPUT41), .B(n518), .ZN(n644) );
  NOR2_X1 U625 ( .A1(n526), .A2(n644), .ZN(n520) );
  XNOR2_X1 U626 ( .A(KEYINPUT105), .B(KEYINPUT42), .ZN(n519) );
  XNOR2_X1 U627 ( .A(n520), .B(n519), .ZN(n757) );
  NAND2_X1 U628 ( .A1(n533), .A2(n531), .ZN(n700) );
  INV_X1 U629 ( .A(n700), .ZN(n697) );
  NAND2_X1 U630 ( .A1(n521), .A2(n697), .ZN(n522) );
  NAND2_X1 U631 ( .A1(n523), .A2(n611), .ZN(n545) );
  XOR2_X1 U632 ( .A(KEYINPUT76), .B(KEYINPUT19), .Z(n524) );
  INV_X1 U633 ( .A(n692), .ZN(n704) );
  NAND2_X1 U634 ( .A1(n700), .A2(n704), .ZN(n596) );
  NAND2_X1 U635 ( .A1(n698), .A2(n596), .ZN(n527) );
  INV_X1 U636 ( .A(n698), .ZN(n529) );
  NAND2_X1 U637 ( .A1(KEYINPUT47), .A2(n529), .ZN(n530) );
  INV_X1 U638 ( .A(n596), .ZN(n615) );
  NAND2_X1 U639 ( .A1(KEYINPUT47), .A2(n615), .ZN(n537) );
  INV_X1 U640 ( .A(n531), .ZN(n532) );
  NOR2_X1 U641 ( .A1(n533), .A2(n532), .ZN(n566) );
  INV_X1 U642 ( .A(n566), .ZN(n534) );
  NOR2_X1 U643 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U644 ( .A1(n555), .A2(n536), .ZN(n696) );
  NAND2_X1 U645 ( .A1(n537), .A2(n696), .ZN(n538) );
  XNOR2_X1 U646 ( .A(n538), .B(KEYINPUT82), .ZN(n547) );
  INV_X1 U647 ( .A(n587), .ZN(n621) );
  XNOR2_X1 U648 ( .A(n541), .B(KEYINPUT6), .ZN(n576) );
  INV_X1 U649 ( .A(n576), .ZN(n582) );
  XNOR2_X1 U650 ( .A(KEYINPUT102), .B(n543), .ZN(n544) );
  NAND2_X1 U651 ( .A1(n544), .A2(n697), .ZN(n550) );
  NOR2_X1 U652 ( .A1(n550), .A2(n545), .ZN(n546) );
  NOR2_X1 U653 ( .A1(n547), .A2(n707), .ZN(n548) );
  INV_X1 U654 ( .A(n550), .ZN(n551) );
  NAND2_X1 U655 ( .A1(n551), .A2(n611), .ZN(n552) );
  NOR2_X1 U656 ( .A1(n587), .A2(n552), .ZN(n553) );
  XNOR2_X1 U657 ( .A(n553), .B(KEYINPUT43), .ZN(n554) );
  NOR2_X1 U658 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U659 ( .A(KEYINPUT103), .B(n556), .ZN(n754) );
  INV_X1 U660 ( .A(n622), .ZN(n588) );
  AND2_X1 U661 ( .A1(n588), .A2(n576), .ZN(n557) );
  XOR2_X1 U662 ( .A(KEYINPUT100), .B(KEYINPUT33), .Z(n558) );
  NOR2_X1 U663 ( .A1(G898), .A2(n560), .ZN(n561) );
  NOR2_X1 U664 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U665 ( .A(n567), .B(KEYINPUT35), .ZN(n752) );
  XNOR2_X1 U666 ( .A(KEYINPUT22), .B(KEYINPUT72), .ZN(n573) );
  NAND2_X1 U667 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U668 ( .A(n570), .B(KEYINPUT99), .ZN(n571) );
  NAND2_X1 U669 ( .A1(n571), .A2(n590), .ZN(n572) );
  NAND2_X1 U670 ( .A1(n583), .A2(n631), .ZN(n574) );
  NOR2_X1 U671 ( .A1(n752), .A2(n691), .ZN(n580) );
  NOR2_X1 U672 ( .A1(n576), .A2(n575), .ZN(n578) );
  NOR2_X1 U673 ( .A1(n625), .A2(n621), .ZN(n577) );
  NAND2_X1 U674 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U675 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U676 ( .A1(n585), .A2(n584), .ZN(n684) );
  INV_X1 U677 ( .A(n684), .ZN(n599) );
  AND2_X1 U678 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U679 ( .A1(n586), .A2(n589), .ZN(n634) );
  INV_X1 U680 ( .A(n590), .ZN(n591) );
  NOR2_X1 U681 ( .A1(n634), .A2(n591), .ZN(n592) );
  XNOR2_X1 U682 ( .A(n592), .B(KEYINPUT31), .ZN(n703) );
  NOR2_X1 U683 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U684 ( .A1(n595), .A2(n631), .ZN(n688) );
  NAND2_X1 U685 ( .A1(n703), .A2(n688), .ZN(n597) );
  NAND2_X1 U686 ( .A1(n597), .A2(n596), .ZN(n598) );
  INV_X1 U687 ( .A(KEYINPUT84), .ZN(n604) );
  XNOR2_X1 U688 ( .A(n600), .B(KEYINPUT2), .ZN(n606) );
  INV_X1 U689 ( .A(n601), .ZN(n743) );
  NAND2_X1 U690 ( .A1(n743), .A2(n732), .ZN(n603) );
  NAND2_X1 U691 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U692 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U693 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U694 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U695 ( .A(n614), .B(KEYINPUT118), .ZN(n618) );
  NOR2_X1 U696 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U697 ( .A1(n618), .A2(n617), .ZN(n619) );
  XOR2_X1 U698 ( .A(KEYINPUT119), .B(n619), .Z(n620) );
  NOR2_X1 U699 ( .A1(n609), .A2(n620), .ZN(n640) );
  NAND2_X1 U700 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U701 ( .A(n623), .B(KEYINPUT50), .ZN(n624) );
  XNOR2_X1 U702 ( .A(KEYINPUT115), .B(n624), .ZN(n630) );
  OR2_X1 U703 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U704 ( .A(n627), .B(KEYINPUT114), .ZN(n628) );
  XNOR2_X1 U705 ( .A(KEYINPUT49), .B(n628), .ZN(n629) );
  NOR2_X1 U706 ( .A1(n630), .A2(n629), .ZN(n632) );
  NAND2_X1 U707 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U708 ( .A(n633), .B(KEYINPUT116), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U710 ( .A(KEYINPUT51), .B(n636), .ZN(n637) );
  NOR2_X1 U711 ( .A1(n644), .A2(n637), .ZN(n638) );
  XOR2_X1 U712 ( .A(KEYINPUT117), .B(n638), .Z(n639) );
  NOR2_X1 U713 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U714 ( .A(n641), .B(KEYINPUT52), .ZN(n642) );
  NOR2_X1 U715 ( .A1(n643), .A2(n642), .ZN(n646) );
  NOR2_X1 U716 ( .A1(n609), .A2(n644), .ZN(n645) );
  NOR2_X1 U717 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U718 ( .A1(n648), .A2(n427), .ZN(n651) );
  XNOR2_X1 U719 ( .A(n649), .B(KEYINPUT53), .ZN(n650) );
  XNOR2_X1 U720 ( .A(n651), .B(n650), .ZN(G75) );
  INV_X1 U721 ( .A(n652), .ZN(n653) );
  NAND2_X1 U722 ( .A1(n653), .A2(KEYINPUT2), .ZN(n654) );
  XOR2_X1 U723 ( .A(KEYINPUT65), .B(n654), .Z(n655) );
  NAND2_X1 U724 ( .A1(KEYINPUT2), .A2(n657), .ZN(n658) );
  XNOR2_X1 U725 ( .A(n660), .B(KEYINPUT64), .ZN(n662) );
  XOR2_X1 U726 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n661) );
  NOR2_X1 U727 ( .A1(G952), .A2(n745), .ZN(n665) );
  INV_X1 U728 ( .A(n719), .ZN(n724) );
  NAND2_X1 U729 ( .A1(n666), .A2(n724), .ZN(n668) );
  XOR2_X1 U730 ( .A(KEYINPUT122), .B(KEYINPUT60), .Z(n667) );
  XNOR2_X1 U731 ( .A(n668), .B(n667), .ZN(G60) );
  NAND2_X1 U732 ( .A1(n720), .A2(G210), .ZN(n672) );
  XOR2_X1 U733 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n669) );
  XNOR2_X1 U734 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U735 ( .A(n672), .B(n671), .ZN(n673) );
  NAND2_X1 U736 ( .A1(n673), .A2(n724), .ZN(n675) );
  INV_X1 U737 ( .A(KEYINPUT56), .ZN(n674) );
  XNOR2_X1 U738 ( .A(n675), .B(n674), .ZN(G51) );
  NAND2_X1 U739 ( .A1(n720), .A2(G472), .ZN(n679) );
  XOR2_X1 U740 ( .A(KEYINPUT62), .B(KEYINPUT106), .Z(n676) );
  NAND2_X1 U741 ( .A1(n680), .A2(n724), .ZN(n683) );
  XOR2_X1 U742 ( .A(KEYINPUT63), .B(KEYINPUT107), .Z(n681) );
  XNOR2_X1 U743 ( .A(KEYINPUT88), .B(n681), .ZN(n682) );
  XNOR2_X1 U744 ( .A(n683), .B(n682), .ZN(G57) );
  XOR2_X1 U745 ( .A(n684), .B(G101), .Z(G3) );
  NOR2_X1 U746 ( .A1(n700), .A2(n688), .ZN(n685) );
  XOR2_X1 U747 ( .A(G104), .B(n685), .Z(G6) );
  XOR2_X1 U748 ( .A(KEYINPUT108), .B(KEYINPUT26), .Z(n687) );
  XNOR2_X1 U749 ( .A(G107), .B(KEYINPUT27), .ZN(n686) );
  XNOR2_X1 U750 ( .A(n687), .B(n686), .ZN(n690) );
  NOR2_X1 U751 ( .A1(n704), .A2(n688), .ZN(n689) );
  XOR2_X1 U752 ( .A(n690), .B(n689), .Z(G9) );
  XOR2_X1 U753 ( .A(n691), .B(G110), .Z(G12) );
  XOR2_X1 U754 ( .A(KEYINPUT109), .B(KEYINPUT29), .Z(n694) );
  NAND2_X1 U755 ( .A1(n698), .A2(n692), .ZN(n693) );
  XNOR2_X1 U756 ( .A(n694), .B(n693), .ZN(n695) );
  XOR2_X1 U757 ( .A(G128), .B(n695), .Z(G30) );
  XNOR2_X1 U758 ( .A(G143), .B(n696), .ZN(G45) );
  NAND2_X1 U759 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U760 ( .A(n699), .B(G146), .ZN(G48) );
  NOR2_X1 U761 ( .A1(n700), .A2(n703), .ZN(n701) );
  XOR2_X1 U762 ( .A(KEYINPUT110), .B(n701), .Z(n702) );
  XNOR2_X1 U763 ( .A(n352), .B(n702), .ZN(G15) );
  NOR2_X1 U764 ( .A1(n704), .A2(n703), .ZN(n706) );
  XNOR2_X1 U765 ( .A(G116), .B(KEYINPUT111), .ZN(n705) );
  XNOR2_X1 U766 ( .A(n706), .B(n705), .ZN(G18) );
  XNOR2_X1 U767 ( .A(n707), .B(KEYINPUT112), .ZN(n708) );
  XNOR2_X1 U768 ( .A(n708), .B(KEYINPUT37), .ZN(n709) );
  XNOR2_X1 U769 ( .A(G125), .B(n709), .ZN(G27) );
  XOR2_X1 U770 ( .A(G134), .B(n710), .Z(G36) );
  NAND2_X1 U771 ( .A1(n720), .A2(G469), .ZN(n714) );
  XOR2_X1 U772 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n712) );
  NOR2_X1 U773 ( .A1(n719), .A2(n715), .ZN(G54) );
  NAND2_X1 U774 ( .A1(G478), .A2(n720), .ZN(n716) );
  XNOR2_X1 U775 ( .A(n717), .B(n716), .ZN(n718) );
  NOR2_X1 U776 ( .A1(n719), .A2(n718), .ZN(G63) );
  XNOR2_X1 U777 ( .A(n726), .B(KEYINPUT125), .ZN(n728) );
  XNOR2_X1 U778 ( .A(n728), .B(n727), .ZN(n729) );
  XNOR2_X1 U779 ( .A(n729), .B(G101), .ZN(n731) );
  NOR2_X1 U780 ( .A1(n745), .A2(G898), .ZN(n730) );
  NOR2_X1 U781 ( .A1(n731), .A2(n730), .ZN(n740) );
  OR2_X1 U782 ( .A1(G953), .A2(n732), .ZN(n737) );
  NAND2_X1 U783 ( .A1(G224), .A2(G953), .ZN(n733) );
  XNOR2_X1 U784 ( .A(n733), .B(KEYINPUT124), .ZN(n734) );
  XNOR2_X1 U785 ( .A(KEYINPUT61), .B(n734), .ZN(n735) );
  NAND2_X1 U786 ( .A1(n735), .A2(G898), .ZN(n736) );
  NAND2_X1 U787 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U788 ( .A(n738), .B(KEYINPUT126), .ZN(n739) );
  XNOR2_X1 U789 ( .A(n740), .B(n739), .ZN(G69) );
  XNOR2_X1 U790 ( .A(n742), .B(n741), .ZN(n747) );
  INV_X1 U791 ( .A(n747), .ZN(n744) );
  XOR2_X1 U792 ( .A(n744), .B(n743), .Z(n746) );
  NAND2_X1 U793 ( .A1(n746), .A2(n745), .ZN(n751) );
  XOR2_X1 U794 ( .A(G227), .B(n747), .Z(n748) );
  NAND2_X1 U795 ( .A1(n748), .A2(G900), .ZN(n749) );
  NAND2_X1 U796 ( .A1(n749), .A2(G953), .ZN(n750) );
  NAND2_X1 U797 ( .A1(n751), .A2(n750), .ZN(G72) );
  XOR2_X1 U798 ( .A(n752), .B(G122), .Z(G24) );
  XOR2_X1 U799 ( .A(G140), .B(KEYINPUT113), .Z(n753) );
  XNOR2_X1 U800 ( .A(n754), .B(n753), .ZN(G42) );
  XOR2_X1 U801 ( .A(G119), .B(n755), .Z(n756) );
  XNOR2_X1 U802 ( .A(KEYINPUT127), .B(n756), .ZN(G21) );
  XNOR2_X1 U803 ( .A(G137), .B(n757), .ZN(G39) );
endmodule

