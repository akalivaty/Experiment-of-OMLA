//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT27), .B(G183gat), .ZN(new_n203));
  INV_X1    g002(.A(G190gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT28), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n209), .A2(KEYINPUT67), .ZN(new_n210));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n209), .ZN(new_n212));
  NOR2_X1   g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT26), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT67), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n210), .B(new_n211), .C1(new_n212), .C2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n207), .A2(new_n208), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT68), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n217), .B(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT25), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n208), .B(KEYINPUT24), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n213), .A2(KEYINPUT23), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n213), .A2(KEYINPUT23), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n213), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n227), .A2(new_n228), .A3(new_n211), .A4(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n220), .B1(new_n224), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n223), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n221), .A2(new_n235), .ZN(new_n236));
  AND3_X1   g035(.A1(new_n225), .A2(KEYINPUT25), .A3(new_n211), .ZN(new_n237));
  AND3_X1   g036(.A1(new_n236), .A2(new_n228), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AND4_X1   g039(.A1(new_n239), .A2(new_n236), .A3(new_n228), .A4(new_n237), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n231), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n219), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G120gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G113gat), .ZN(new_n245));
  INV_X1    g044(.A(G113gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G120gat), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT1), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G127gat), .B(G134gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT69), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n248), .A2(new_n249), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n243), .A2(new_n254), .ZN(new_n255));
  OR2_X1    g054(.A1(new_n217), .A2(new_n218), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n217), .A2(new_n218), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n238), .B(new_n239), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n256), .A2(new_n257), .B1(new_n258), .B2(new_n231), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(new_n253), .ZN(new_n260));
  INV_X1    g059(.A(G227gat), .ZN(new_n261));
  INV_X1    g060(.A(G233gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n255), .A2(new_n260), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT32), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n264), .A2(KEYINPUT70), .A3(KEYINPUT32), .ZN(new_n268));
  XOR2_X1   g067(.A(G15gat), .B(G43gat), .Z(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(KEYINPUT71), .ZN(new_n270));
  XNOR2_X1  g069(.A(G71gat), .B(G99gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT33), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n272), .B1(new_n264), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n267), .A2(new_n268), .A3(new_n274), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n264), .B(KEYINPUT32), .C1(new_n273), .C2(new_n272), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT34), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n255), .A2(new_n260), .ZN(new_n279));
  INV_X1    g078(.A(new_n263), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  AOI211_X1 g080(.A(KEYINPUT34), .B(new_n263), .C1(new_n255), .C2(new_n260), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n277), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G22gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(G197gat), .B(G204gat), .ZN(new_n287));
  INV_X1    g086(.A(G211gat), .ZN(new_n288));
  INV_X1    g087(.A(G218gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n287), .B1(KEYINPUT22), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G211gat), .B(G218gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT29), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT3), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(KEYINPUT76), .B(G141gat), .Z(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G148gat), .ZN(new_n298));
  INV_X1    g097(.A(G148gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G141gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301));
  OR3_X1    g100(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n298), .A2(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OR2_X1    g102(.A1(new_n299), .A2(G141gat), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT2), .B1(new_n304), .B2(new_n300), .ZN(new_n305));
  INV_X1    g104(.A(G155gat), .ZN(new_n306));
  INV_X1    g105(.A(G162gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n306), .A2(new_n307), .A3(KEYINPUT75), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT75), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n309), .B1(G155gat), .B2(G162gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(new_n310), .A3(new_n301), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n305), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n303), .A2(new_n312), .ZN(new_n313));
  OAI211_X1 g112(.A(G228gat), .B(G233gat), .C1(new_n296), .C2(new_n313), .ZN(new_n314));
  OR3_X1    g113(.A1(new_n303), .A2(KEYINPUT3), .A3(new_n312), .ZN(new_n315));
  XOR2_X1   g114(.A(KEYINPUT73), .B(KEYINPUT29), .Z(new_n316));
  AOI21_X1  g115(.A(new_n294), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G228gat), .A2(G233gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n320), .B(KEYINPUT78), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n316), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n293), .A2(new_n323), .ZN(new_n324));
  OR2_X1    g123(.A1(new_n324), .A2(KEYINPUT79), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT3), .B1(new_n324), .B2(KEYINPUT79), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n313), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n322), .B1(new_n327), .B2(new_n317), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n286), .B1(new_n319), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n319), .A2(new_n328), .A3(new_n286), .ZN(new_n331));
  XNOR2_X1  g130(.A(G78gat), .B(G106gat), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n332), .ZN(new_n334));
  INV_X1    g133(.A(new_n331), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n334), .B1(new_n335), .B2(new_n329), .ZN(new_n336));
  XOR2_X1   g135(.A(KEYINPUT31), .B(G50gat), .Z(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n333), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n333), .A2(new_n336), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(new_n337), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n275), .A2(new_n283), .A3(new_n276), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n285), .A2(new_n339), .A3(new_n341), .A4(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n344));
  NAND2_X1  g143(.A1(G226gat), .A2(G233gat), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n344), .B1(new_n259), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n345), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n243), .A2(KEYINPUT74), .A3(new_n347), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n242), .A2(new_n217), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n345), .B1(new_n349), .B2(KEYINPUT29), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n346), .A2(new_n348), .A3(new_n350), .A4(new_n294), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n323), .A2(new_n347), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n243), .A2(new_n352), .B1(new_n349), .B2(new_n347), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n293), .ZN(new_n354));
  XNOR2_X1  g153(.A(G8gat), .B(G36gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(G64gat), .B(G92gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n351), .A2(new_n354), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT30), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n358), .B1(new_n351), .B2(new_n354), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n359), .A2(KEYINPUT30), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n313), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n253), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT4), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(KEYINPUT3), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(new_n253), .A3(new_n315), .ZN(new_n370));
  NAND2_X1  g169(.A1(G225gat), .A2(G233gat), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT4), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n372), .B1(new_n253), .B2(new_n366), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n368), .A2(new_n370), .A3(new_n371), .A4(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT5), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n371), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n254), .A2(new_n313), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n378), .B1(new_n379), .B2(new_n367), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n375), .B1(new_n374), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G1gat), .B(G29gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(KEYINPUT0), .ZN(new_n383));
  XNOR2_X1  g182(.A(G57gat), .B(G85gat), .ZN(new_n384));
  XOR2_X1   g183(.A(new_n383), .B(new_n384), .Z(new_n385));
  NOR3_X1   g184(.A1(new_n377), .A2(new_n381), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n386), .A2(KEYINPUT77), .A3(KEYINPUT6), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n374), .A2(new_n380), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT5), .ZN(new_n389));
  INV_X1    g188(.A(new_n385), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(new_n390), .A3(new_n376), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n385), .B1(new_n377), .B2(new_n381), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT6), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n389), .A2(KEYINPUT6), .A3(new_n390), .A4(new_n376), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT77), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n387), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n365), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n202), .B1(new_n343), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n399), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n341), .A2(new_n339), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n275), .A2(new_n283), .A3(new_n276), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n283), .B1(new_n275), .B2(new_n276), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n401), .A2(new_n402), .A3(new_n405), .A4(KEYINPUT35), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT36), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n407), .B1(new_n405), .B2(KEYINPUT72), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n285), .A2(new_n342), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT72), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT36), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n341), .A2(new_n339), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n399), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n408), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n368), .A2(new_n370), .A3(new_n373), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n378), .ZN(new_n416));
  OR2_X1    g215(.A1(new_n416), .A2(KEYINPUT39), .ZN(new_n417));
  OR2_X1    g216(.A1(new_n379), .A2(new_n367), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n416), .B(KEYINPUT39), .C1(new_n378), .C2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n417), .A2(new_n419), .A3(new_n385), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT40), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n417), .A2(new_n419), .A3(KEYINPUT40), .A4(new_n385), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(new_n391), .A3(new_n423), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n339), .B(new_n341), .C1(new_n365), .C2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n358), .A2(KEYINPUT38), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT37), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n428), .B1(new_n353), .B2(new_n294), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n346), .A2(new_n348), .A3(new_n350), .A4(new_n293), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n427), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n351), .A2(new_n428), .A3(new_n354), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n359), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n398), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT80), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n351), .A2(new_n354), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT37), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n438), .A2(new_n357), .A3(new_n432), .ZN(new_n439));
  AOI22_X1  g238(.A1(new_n435), .A2(new_n436), .B1(KEYINPUT38), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT80), .B1(new_n398), .B2(new_n434), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n425), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n400), .B(new_n406), .C1(new_n414), .C2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT87), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT86), .B(G1gat), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT16), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(G15gat), .B(G22gat), .ZN(new_n448));
  INV_X1    g247(.A(G1gat), .ZN(new_n449));
  AND2_X1   g248(.A1(new_n449), .A2(KEYINPUT86), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(KEYINPUT86), .ZN(new_n451));
  OAI211_X1 g250(.A(KEYINPUT87), .B(KEYINPUT16), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n447), .A2(new_n448), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(G8gat), .ZN(new_n454));
  OR2_X1    g253(.A1(new_n448), .A2(G1gat), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n454), .B1(new_n453), .B2(new_n455), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(G71gat), .A2(G78gat), .ZN(new_n459));
  INV_X1    g258(.A(G71gat), .ZN(new_n460));
  INV_X1    g259(.A(G78gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT9), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(KEYINPUT90), .A2(G57gat), .ZN(new_n465));
  AND2_X1   g264(.A1(KEYINPUT91), .A2(G64gat), .ZN(new_n466));
  NOR2_X1   g265(.A1(KEYINPUT91), .A2(G64gat), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT91), .ZN(new_n469));
  INV_X1    g268(.A(G64gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AND2_X1   g270(.A1(KEYINPUT90), .A2(G57gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(KEYINPUT91), .A2(G64gat), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n464), .A2(new_n468), .A3(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G57gat), .B(G64gat), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n459), .B(new_n462), .C1(new_n476), .C2(new_n463), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT92), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n478), .B(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT21), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n458), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  XOR2_X1   g281(.A(new_n482), .B(KEYINPUT93), .Z(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G183gat), .B(G211gat), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n478), .A2(new_n481), .ZN(new_n487));
  NAND2_X1  g286(.A1(G231gat), .A2(G233gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G127gat), .B(G155gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  XOR2_X1   g290(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n491), .A2(new_n492), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n486), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n494), .A2(new_n495), .A3(new_n486), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n484), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n498), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(new_n483), .A3(new_n496), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  XOR2_X1   g301(.A(G134gat), .B(G162gat), .Z(new_n503));
  AND2_X1   g302(.A1(G232gat), .A2(G233gat), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n504), .A2(KEYINPUT41), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n503), .B(new_n505), .Z(new_n506));
  XOR2_X1   g305(.A(new_n506), .B(KEYINPUT94), .Z(new_n507));
  XNOR2_X1  g306(.A(G190gat), .B(G218gat), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G99gat), .B(G106gat), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(KEYINPUT95), .A2(KEYINPUT7), .ZN(new_n512));
  NAND2_X1  g311(.A1(G85gat), .A2(G92gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(G99gat), .A2(G106gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT8), .ZN(new_n516));
  OR2_X1    g315(.A1(G85gat), .A2(G92gat), .ZN(new_n517));
  OR2_X1    g316(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n514), .A2(new_n516), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(KEYINPUT96), .A2(G85gat), .A3(G92gat), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n520), .A2(new_n512), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n511), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT8), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n523), .B1(G99gat), .B2(G106gat), .ZN(new_n524));
  OAI22_X1  g323(.A1(KEYINPUT96), .A2(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n520), .A2(new_n512), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n526), .A2(new_n510), .A3(new_n527), .A4(new_n514), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n522), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT15), .ZN(new_n530));
  INV_X1    g329(.A(G43gat), .ZN(new_n531));
  INV_X1    g330(.A(G50gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G43gat), .A2(G50gat), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n530), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT14), .ZN(new_n536));
  INV_X1    g335(.A(G29gat), .ZN(new_n537));
  INV_X1    g336(.A(G36gat), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n539), .A2(KEYINPUT84), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G29gat), .A2(G36gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT84), .B1(new_n539), .B2(new_n540), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n535), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n533), .A2(KEYINPUT85), .A3(new_n534), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT15), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n533), .A2(KEYINPUT85), .A3(new_n530), .A4(new_n534), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n539), .A2(new_n540), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n548), .A2(new_n549), .A3(new_n550), .A4(new_n542), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n545), .A2(new_n546), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n546), .B1(new_n545), .B2(new_n551), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n529), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT97), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g356(.A(KEYINPUT97), .B(new_n529), .C1(new_n553), .C2(new_n554), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n529), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n551), .ZN(new_n561));
  AOI22_X1  g360(.A1(new_n560), .A2(new_n561), .B1(KEYINPUT41), .B2(new_n504), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n509), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n562), .ZN(new_n564));
  AOI211_X1 g363(.A(new_n564), .B(new_n508), .C1(new_n557), .C2(new_n558), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n507), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT98), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g367(.A(KEYINPUT98), .B(new_n507), .C1(new_n563), .C2(new_n565), .ZN(new_n569));
  INV_X1    g368(.A(new_n558), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n561), .A2(KEYINPUT17), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(new_n552), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT97), .B1(new_n572), .B2(new_n529), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n562), .B(new_n509), .C1(new_n570), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(new_n506), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT99), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n562), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(new_n508), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n575), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n563), .A2(KEYINPUT99), .ZN(new_n580));
  AOI22_X1  g379(.A1(new_n568), .A2(new_n569), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n502), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT83), .ZN(new_n583));
  XOR2_X1   g382(.A(G113gat), .B(G141gat), .Z(new_n584));
  XNOR2_X1  g383(.A(G169gat), .B(G197gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(KEYINPUT81), .B(KEYINPUT11), .Z(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT82), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n586), .B(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT12), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n561), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n458), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n453), .A2(new_n455), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(G8gat), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT88), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n597), .A2(new_n598), .B1(new_n571), .B2(new_n552), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n595), .A2(new_n596), .A3(KEYINPUT88), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n593), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT89), .ZN(new_n602));
  NAND2_X1  g401(.A1(G229gat), .A2(G233gat), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n601), .A2(new_n602), .A3(KEYINPUT18), .A4(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n598), .B1(new_n456), .B2(new_n457), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n572), .A2(new_n605), .A3(new_n600), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n597), .A2(new_n561), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n606), .A2(KEYINPUT18), .A3(new_n603), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT89), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n606), .A2(new_n603), .A3(new_n607), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT18), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n458), .A2(new_n592), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n607), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n603), .B(KEYINPUT13), .Z(new_n615));
  AOI22_X1  g414(.A1(new_n611), .A2(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AOI211_X1 g415(.A(new_n583), .B(new_n591), .C1(new_n610), .C2(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n608), .A2(KEYINPUT89), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n608), .A2(KEYINPUT89), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n616), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n590), .B1(new_n620), .B2(KEYINPUT83), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n560), .A2(KEYINPUT10), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n480), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT100), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n475), .A2(new_n477), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n529), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n478), .A2(new_n528), .A3(new_n522), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT10), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n626), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI211_X1 g431(.A(KEYINPUT100), .B(KEYINPUT10), .C1(new_n628), .C2(new_n629), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n625), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G230gat), .A2(G233gat), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n636), .B1(new_n630), .B2(new_n635), .ZN(new_n637));
  XOR2_X1   g436(.A(G120gat), .B(G148gat), .Z(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT101), .ZN(new_n639));
  XOR2_X1   g438(.A(G176gat), .B(G204gat), .Z(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n637), .A2(new_n641), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n582), .A2(new_n623), .A3(new_n644), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n443), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n398), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(G1gat), .ZN(G1324gat));
  INV_X1    g448(.A(new_n365), .ZN(new_n650));
  XOR2_X1   g449(.A(KEYINPUT16), .B(G8gat), .Z(new_n651));
  NAND3_X1  g450(.A1(new_n646), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT42), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n654), .B(KEYINPUT103), .Z(new_n655));
  NAND2_X1  g454(.A1(new_n652), .A2(new_n653), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n454), .B1(new_n646), .B2(new_n650), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT102), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n655), .A2(new_n656), .A3(new_n658), .ZN(G1325gat));
  INV_X1    g458(.A(new_n646), .ZN(new_n660));
  OR3_X1    g459(.A1(new_n660), .A2(G15gat), .A3(new_n409), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n408), .A2(new_n411), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(G15gat), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n661), .A2(new_n664), .ZN(G1326gat));
  NAND2_X1  g464(.A1(new_n646), .A2(new_n412), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT43), .B(G22gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(G1327gat));
  AND2_X1   g467(.A1(new_n387), .A2(new_n397), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n360), .B1(new_n432), .B2(new_n431), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n669), .A2(new_n670), .A3(new_n436), .A4(new_n394), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n439), .A2(KEYINPUT38), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n671), .A2(new_n441), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n425), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n675), .A2(new_n411), .A3(new_n408), .A4(new_n413), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n400), .A2(new_n406), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n581), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n678), .A2(KEYINPUT44), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(KEYINPUT44), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n502), .ZN(new_n682));
  INV_X1    g481(.A(new_n644), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n682), .A2(new_n622), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT104), .Z(new_n685));
  NAND2_X1  g484(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(G29gat), .B1(new_n686), .B2(new_n398), .ZN(new_n687));
  AOI211_X1 g486(.A(new_n581), .B(new_n684), .C1(new_n676), .C2(new_n677), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n688), .A2(new_n537), .A3(new_n647), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT45), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n687), .A2(new_n690), .ZN(G1328gat));
  NAND3_X1  g490(.A1(new_n688), .A2(new_n538), .A3(new_n650), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(KEYINPUT46), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT105), .ZN(new_n694));
  OAI21_X1  g493(.A(G36gat), .B1(new_n686), .B2(new_n365), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n692), .A2(KEYINPUT46), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(G1329gat));
  NAND2_X1  g496(.A1(new_n688), .A2(new_n405), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n531), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n662), .A2(G43gat), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n699), .B1(new_n686), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(KEYINPUT47), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT47), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n703), .B(new_n699), .C1(new_n686), .C2(new_n700), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(G1330gat));
  NAND2_X1  g504(.A1(new_n688), .A2(new_n412), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n532), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n412), .A2(G50gat), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n707), .B1(new_n686), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(KEYINPUT48), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT48), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n711), .B(new_n707), .C1(new_n686), .C2(new_n708), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(G1331gat));
  NOR2_X1   g512(.A1(new_n582), .A2(new_n622), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n644), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT106), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n716), .B1(new_n676), .B2(new_n677), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n647), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(G57gat), .ZN(G1332gat));
  INV_X1    g518(.A(KEYINPUT49), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n650), .B1(new_n720), .B2(new_n470), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT107), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n717), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n720), .A2(new_n470), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1333gat));
  AOI21_X1  g524(.A(G71gat), .B1(new_n717), .B2(new_n405), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n663), .A2(new_n460), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n726), .B1(new_n717), .B2(new_n727), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n728), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g528(.A1(new_n717), .A2(new_n412), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g530(.A1(new_n502), .A2(new_n622), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n644), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n681), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(G85gat), .B1(new_n735), .B2(new_n398), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n568), .A2(new_n569), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n579), .A2(new_n580), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n443), .A2(KEYINPUT51), .A3(new_n739), .A4(new_n732), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n678), .A2(KEYINPUT108), .A3(KEYINPUT51), .A4(new_n732), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n678), .A2(new_n732), .ZN(new_n745));
  AOI22_X1  g544(.A1(new_n742), .A2(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OR3_X1    g545(.A1(new_n398), .A2(G85gat), .A3(new_n683), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n736), .B1(new_n746), .B2(new_n747), .ZN(G1336gat));
  NAND4_X1  g547(.A1(new_n679), .A2(new_n680), .A3(new_n650), .A4(new_n734), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT52), .B1(new_n749), .B2(G92gat), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n742), .A2(new_n743), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n745), .A2(new_n744), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n365), .A2(G92gat), .A3(new_n683), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n751), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n755), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n746), .A2(KEYINPUT110), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n750), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n745), .A2(KEYINPUT109), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT109), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n761), .B1(new_n678), .B2(new_n732), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n744), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n757), .B1(new_n763), .B2(new_n752), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n749), .A2(G92gat), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT52), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n759), .A2(new_n766), .ZN(G1337gat));
  OAI21_X1  g566(.A(G99gat), .B1(new_n735), .B2(new_n663), .ZN(new_n768));
  OR3_X1    g567(.A1(new_n409), .A2(G99gat), .A3(new_n683), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n746), .B2(new_n769), .ZN(G1338gat));
  NOR3_X1   g569(.A1(new_n402), .A2(G106gat), .A3(new_n683), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n772), .B1(new_n763), .B2(new_n752), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n679), .A2(new_n680), .A3(new_n412), .A4(new_n734), .ZN(new_n774));
  XNOR2_X1  g573(.A(KEYINPUT111), .B(G106gat), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT53), .B1(new_n773), .B2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n776), .B(new_n779), .C1(new_n746), .C2(new_n772), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(G1339gat));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n782), .B1(new_n634), .B2(new_n635), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n480), .A2(new_n624), .ZN(new_n785));
  INV_X1    g584(.A(new_n629), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n478), .B1(new_n528), .B2(new_n522), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n631), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT100), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n630), .A2(new_n626), .A3(new_n631), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n785), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n635), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n784), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n625), .B(new_n792), .C1(new_n632), .C2(new_n633), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(KEYINPUT112), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n783), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n634), .A2(new_n782), .A3(new_n635), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n641), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n796), .A2(KEYINPUT55), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n642), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT113), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n800), .A2(KEYINPUT113), .A3(new_n642), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n796), .A2(new_n799), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n803), .A2(new_n622), .A3(new_n804), .A4(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n610), .A2(new_n616), .A3(new_n590), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n601), .A2(new_n603), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n614), .A2(new_n615), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n589), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n644), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n739), .B1(new_n808), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n804), .A2(new_n807), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT113), .B1(new_n800), .B2(new_n642), .ZN(new_n818));
  NOR4_X1   g617(.A1(new_n817), .A2(new_n818), .A3(new_n581), .A4(new_n813), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n682), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n582), .A2(new_n622), .A3(new_n644), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n650), .A2(new_n398), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n343), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(new_n623), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(new_n246), .ZN(G1340gat));
  NOR2_X1   g628(.A1(new_n827), .A2(new_n683), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(new_n244), .ZN(G1341gat));
  NOR2_X1   g630(.A1(new_n827), .A2(new_n682), .ZN(new_n832));
  XNOR2_X1  g631(.A(KEYINPUT114), .B(G127gat), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n832), .B(new_n833), .ZN(G1342gat));
  NAND3_X1  g633(.A1(new_n825), .A2(new_n826), .A3(new_n739), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n835), .A2(G134gat), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(KEYINPUT56), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(G134gat), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT115), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(G1343gat));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n823), .A2(new_n841), .A3(new_n412), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n408), .A2(new_n411), .A3(new_n824), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n637), .A2(new_n641), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n791), .A2(new_n784), .A3(new_n792), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n794), .A2(KEYINPUT112), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n798), .B1(new_n849), .B2(new_n783), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n846), .B1(new_n850), .B2(KEYINPUT55), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n620), .A2(KEYINPUT83), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n591), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n620), .A2(KEYINPUT83), .A3(new_n590), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n851), .A2(new_n853), .A3(new_n807), .A4(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n739), .B1(new_n855), .B2(new_n815), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n682), .B1(new_n819), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(KEYINPUT116), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT116), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n859), .B(new_n682), .C1(new_n819), .C2(new_n856), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n858), .A2(new_n822), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n841), .B1(new_n861), .B2(new_n412), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n845), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n297), .B1(new_n863), .B2(new_n622), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n662), .A2(new_n402), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n825), .A2(new_n865), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n866), .A2(G141gat), .A3(new_n623), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT58), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n297), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n870), .B1(new_n863), .B2(new_n622), .ZN(new_n871));
  NOR4_X1   g670(.A1(new_n845), .A2(new_n862), .A3(KEYINPUT117), .A4(new_n623), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT58), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n623), .A2(G141gat), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n874), .B1(new_n866), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT118), .B1(new_n873), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n402), .B1(new_n820), .B2(new_n822), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n843), .B1(new_n879), .B2(new_n841), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n821), .B1(new_n857), .B2(KEYINPUT116), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n402), .B1(new_n881), .B2(new_n860), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n880), .B(new_n622), .C1(new_n841), .C2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT117), .ZN(new_n884));
  INV_X1    g683(.A(new_n862), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n885), .A2(new_n870), .A3(new_n622), .A4(new_n880), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n297), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n887), .A2(new_n888), .A3(new_n876), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n868), .B1(new_n878), .B2(new_n889), .ZN(G1344gat));
  INV_X1    g689(.A(new_n866), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n299), .A3(new_n644), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n803), .A2(new_n739), .A3(new_n804), .A4(new_n807), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n804), .A2(new_n807), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n897), .A2(KEYINPUT119), .A3(new_n739), .A4(new_n803), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n813), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n682), .B1(new_n899), .B2(new_n856), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n822), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT57), .B1(new_n901), .B2(new_n412), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(KEYINPUT120), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT120), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n402), .B1(new_n900), .B2(new_n822), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(KEYINPUT57), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n879), .A2(KEYINPUT57), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n903), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n644), .A3(new_n844), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n893), .B1(new_n909), .B2(G148gat), .ZN(new_n910));
  AOI211_X1 g709(.A(KEYINPUT59), .B(new_n299), .C1(new_n863), .C2(new_n644), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n892), .B1(new_n910), .B2(new_n911), .ZN(G1345gat));
  INV_X1    g711(.A(new_n863), .ZN(new_n913));
  OAI21_X1  g712(.A(G155gat), .B1(new_n913), .B2(new_n682), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n891), .A2(new_n306), .A3(new_n502), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1346gat));
  OAI21_X1  g715(.A(G162gat), .B1(new_n913), .B2(new_n581), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n891), .A2(new_n307), .A3(new_n739), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1347gat));
  NAND2_X1  g718(.A1(new_n650), .A2(new_n398), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT122), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n921), .A2(new_n343), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(new_n823), .ZN(new_n923));
  INV_X1    g722(.A(G169gat), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n923), .A2(new_n924), .A3(new_n623), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n823), .A2(new_n398), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n926), .A2(KEYINPUT121), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n926), .A2(KEYINPUT121), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n650), .B(new_n826), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n929), .A2(new_n623), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n925), .B1(new_n930), .B2(new_n924), .ZN(G1348gat));
  OAI21_X1  g730(.A(G176gat), .B1(new_n923), .B2(new_n683), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n683), .A2(G176gat), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n929), .B2(new_n933), .ZN(G1349gat));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n935), .B1(new_n923), .B2(new_n682), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n922), .A2(KEYINPUT123), .A3(new_n502), .A4(new_n823), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(G183gat), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n502), .A2(new_n203), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n929), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g740(.A(G190gat), .B1(new_n923), .B2(new_n581), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT61), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n739), .A2(new_n204), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n929), .B2(new_n944), .ZN(G1351gat));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n946));
  XOR2_X1   g745(.A(KEYINPUT124), .B(G197gat), .Z(new_n947));
  NOR2_X1   g746(.A1(new_n921), .A2(new_n662), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(new_n907), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n950), .B1(new_n902), .B2(KEYINPUT120), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n949), .B1(new_n951), .B2(new_n906), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n947), .B1(new_n952), .B2(new_n622), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n650), .B(new_n865), .C1(new_n927), .C2(new_n928), .ZN(new_n954));
  INV_X1    g753(.A(new_n947), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n954), .A2(new_n623), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n946), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n908), .A2(new_n622), .A3(new_n948), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(new_n955), .ZN(new_n959));
  INV_X1    g758(.A(new_n956), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n959), .A2(new_n960), .A3(KEYINPUT125), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n957), .A2(new_n961), .ZN(G1352gat));
  OR2_X1    g761(.A1(new_n683), .A2(G204gat), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n954), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT62), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n908), .A2(new_n644), .A3(new_n948), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(G204gat), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n965), .A2(new_n967), .ZN(G1353gat));
  NAND3_X1  g767(.A1(new_n908), .A2(new_n502), .A3(new_n948), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n969), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n970));
  AOI21_X1  g769(.A(KEYINPUT63), .B1(new_n969), .B2(G211gat), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n502), .A2(new_n288), .ZN(new_n972));
  OAI22_X1  g771(.A1(new_n970), .A2(new_n971), .B1(new_n954), .B2(new_n972), .ZN(G1354gat));
  OAI21_X1  g772(.A(new_n289), .B1(new_n954), .B2(new_n581), .ZN(new_n974));
  OR2_X1    g773(.A1(new_n974), .A2(KEYINPUT126), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(KEYINPUT126), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n739), .A2(G218gat), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n977), .B(KEYINPUT127), .ZN(new_n978));
  AOI22_X1  g777(.A1(new_n975), .A2(new_n976), .B1(new_n952), .B2(new_n978), .ZN(G1355gat));
endmodule


