//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n554, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n806, new_n807, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XNOR2_X1  g014(.A(KEYINPUT67), .B(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT68), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  OR4_X1    g029(.A1(G237), .A2(G238), .A3(G235), .A4(G236), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(new_n459), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(new_n459), .ZN(new_n463));
  INV_X1    g038(.A(G137), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT70), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n462), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n466), .B1(new_n467), .B2(new_n459), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n469), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n465), .B1(new_n468), .B2(new_n475), .ZN(G160));
  OR2_X1    g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n459), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n459), .A2(G112), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(G136), .ZN(new_n484));
  OR3_X1    g059(.A1(new_n463), .A2(KEYINPUT71), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(KEYINPUT71), .B1(new_n463), .B2(new_n484), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(G162));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n488), .A2(new_n459), .A3(G138), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT73), .B1(new_n472), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT73), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR3_X1   g067(.A1(new_n492), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n462), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n459), .C1(new_n470), .C2(new_n471), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n490), .A2(new_n494), .B1(KEYINPUT4), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n459), .A2(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT72), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n500), .A2(new_n502), .A3(new_n503), .A4(G2104), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n479), .A2(G126), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n496), .A2(new_n507), .ZN(G164));
  AOI21_X1  g083(.A(G543), .B1(KEYINPUT74), .B2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(KEYINPUT74), .A2(KEYINPUT5), .A3(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n513));
  XOR2_X1   g088(.A(KEYINPUT6), .B(G651), .Z(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n512), .A2(G62), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT75), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n516), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n515), .A2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  INV_X1    g097(.A(KEYINPUT76), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n514), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT6), .B(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(KEYINPUT76), .ZN(new_n526));
  AND3_X1   g101(.A1(new_n524), .A2(G543), .A3(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  INV_X1    g106(.A(new_n511), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n509), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n514), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  XOR2_X1   g110(.A(KEYINPUT77), .B(G89), .Z(new_n536));
  OAI211_X1 g111(.A(new_n529), .B(new_n531), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n528), .A2(new_n537), .ZN(G168));
  NAND2_X1  g113(.A1(new_n527), .A2(G52), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n516), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n534), .A2(G90), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n539), .A2(new_n541), .A3(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  AOI22_X1  g119(.A1(new_n527), .A2(G43), .B1(G81), .B2(new_n534), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n512), .A2(G56), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n516), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n545), .B1(KEYINPUT78), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n548), .A2(KEYINPUT78), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  NAND4_X1  g131(.A1(new_n524), .A2(G53), .A3(G543), .A4(new_n526), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT9), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n533), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n561), .A2(G651), .B1(new_n534), .B2(G91), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(G299));
  INV_X1    g138(.A(G168), .ZN(G286));
  NAND2_X1  g139(.A1(new_n527), .A2(G49), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n512), .A2(G74), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n566), .A2(G651), .B1(new_n534), .B2(G87), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(G288));
  INV_X1    g143(.A(G61), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(new_n510), .B2(new_n511), .ZN(new_n570));
  AND2_X1   g145(.A1(G73), .A2(G543), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(G86), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n573), .B1(new_n510), .B2(new_n511), .ZN(new_n574));
  NAND2_X1  g149(.A1(G48), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n525), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n572), .A2(new_n577), .ZN(G305));
  NAND2_X1  g153(.A1(new_n527), .A2(G47), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n534), .A2(G85), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n579), .B(new_n580), .C1(new_n516), .C2(new_n581), .ZN(G290));
  INV_X1    g157(.A(G868), .ZN(new_n583));
  NOR2_X1   g158(.A1(G301), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n534), .A2(G92), .ZN(new_n585));
  XOR2_X1   g160(.A(new_n585), .B(KEYINPUT10), .Z(new_n586));
  AOI22_X1  g161(.A1(new_n512), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(new_n516), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT79), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n524), .A2(G54), .A3(G543), .A4(new_n526), .ZN(new_n590));
  AND3_X1   g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n589), .B1(new_n588), .B2(new_n590), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n586), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT80), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n584), .B1(new_n594), .B2(new_n583), .ZN(G284));
  AOI21_X1  g170(.A(new_n584), .B1(new_n594), .B2(new_n583), .ZN(G321));
  NAND2_X1  g171(.A1(G299), .A2(new_n583), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(new_n583), .B2(G168), .ZN(G297));
  OAI21_X1  g173(.A(new_n597), .B1(new_n583), .B2(G168), .ZN(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n594), .B1(new_n600), .B2(G860), .ZN(G148));
  NAND2_X1  g176(.A1(new_n594), .A2(new_n600), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  OR3_X1    g178(.A1(new_n603), .A2(KEYINPUT81), .A3(new_n583), .ZN(new_n604));
  OAI21_X1  g179(.A(KEYINPUT81), .B1(new_n603), .B2(new_n583), .ZN(new_n605));
  OAI211_X1 g180(.A(new_n604), .B(new_n605), .C1(G868), .C2(new_n551), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g182(.A1(new_n479), .A2(G123), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n459), .A2(G111), .ZN(new_n609));
  OAI21_X1  g184(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n463), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n611), .B1(G135), .B2(new_n612), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT82), .Z(new_n614));
  XNOR2_X1  g189(.A(KEYINPUT83), .B(G2096), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n462), .A2(new_n460), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT12), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT13), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2100), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n616), .A2(new_n620), .ZN(G156));
  XNOR2_X1  g196(.A(G2427), .B(G2438), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2430), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2435), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n625), .A2(KEYINPUT14), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(G1341), .B(G1348), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2443), .B(G2446), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n627), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G2451), .B(G2454), .Z(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n631), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(G14), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT85), .ZN(G401));
  INV_X1    g213(.A(KEYINPUT18), .ZN(new_n639));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  XNOR2_X1  g215(.A(G2067), .B(G2678), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(KEYINPUT17), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n640), .A2(new_n641), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n639), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(G2100), .Z(new_n646));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  AOI21_X1  g222(.A(new_n647), .B1(new_n642), .B2(KEYINPUT18), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(G2096), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(new_n649), .ZN(G227));
  XNOR2_X1  g225(.A(G1956), .B(G2474), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1961), .B(G1966), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1971), .B(G1976), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT19), .Z(new_n655));
  NOR2_X1   g230(.A1(new_n651), .A2(new_n652), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n653), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT86), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n658), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n655), .A2(new_n656), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT20), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1991), .B(G1996), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1981), .B(G1986), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G229));
  MUX2_X1   g245(.A(G24), .B(G290), .S(G16), .Z(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(G1986), .Z(new_n672));
  INV_X1    g247(.A(G29), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(G25), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT87), .Z(new_n675));
  NAND2_X1  g250(.A1(new_n479), .A2(G119), .ZN(new_n676));
  OR2_X1    g251(.A1(G95), .A2(G2105), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n677), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n678));
  INV_X1    g253(.A(G131), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n676), .B(new_n678), .C1(new_n679), .C2(new_n463), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n675), .B1(new_n681), .B2(new_n673), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT35), .B(G1991), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(G16), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G22), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT88), .Z(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(G303), .B2(G16), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1971), .ZN(new_n689));
  NOR2_X1   g264(.A1(G6), .A2(G16), .ZN(new_n690));
  INV_X1    g265(.A(G305), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(G16), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT32), .B(G1981), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n685), .A2(G23), .ZN(new_n695));
  INV_X1    g270(.A(G288), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n685), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT33), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n698), .A2(G1976), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n698), .A2(G1976), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n689), .B(new_n694), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n672), .B(new_n684), .C1(new_n701), .C2(KEYINPUT34), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT89), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n701), .A2(KEYINPUT34), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(KEYINPUT36), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT36), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n704), .A2(new_n708), .A3(new_n705), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT25), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G139), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(new_n463), .ZN(new_n714));
  NAND2_X1  g289(.A1(G115), .A2(G2104), .ZN(new_n715));
  INV_X1    g290(.A(G127), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n472), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n714), .B1(G2105), .B2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT90), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT91), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n722), .A2(new_n673), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n673), .A2(G33), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G2072), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n685), .A2(G4), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n594), .B2(new_n685), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G1348), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(G1348), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n685), .A2(G20), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT23), .Z(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G299), .B2(G16), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G1956), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n727), .A2(new_n730), .A3(new_n731), .A4(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT97), .ZN(new_n737));
  OAI21_X1  g312(.A(KEYINPUT95), .B1(G29), .B2(G32), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n460), .A2(G105), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(KEYINPUT94), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(KEYINPUT94), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n740), .A2(new_n741), .B1(new_n612), .B2(G141), .ZN(new_n742));
  NAND3_X1  g317(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT26), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G129), .B2(new_n479), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n746), .A2(new_n673), .ZN(new_n747));
  MUX2_X1   g322(.A(new_n738), .B(KEYINPUT95), .S(new_n747), .Z(new_n748));
  XOR2_X1   g323(.A(KEYINPUT27), .B(G1996), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n614), .A2(G29), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n479), .A2(G128), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n459), .A2(G116), .ZN(new_n753));
  OAI21_X1  g328(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n754));
  INV_X1    g329(.A(G140), .ZN(new_n755));
  OAI221_X1 g330(.A(new_n752), .B1(new_n753), .B2(new_n754), .C1(new_n755), .C2(new_n463), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G29), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n673), .A2(G26), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT28), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G2067), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT31), .B(G11), .Z(new_n763));
  INV_X1    g338(.A(G28), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n764), .A2(KEYINPUT30), .ZN(new_n765));
  AOI21_X1  g340(.A(G29), .B1(new_n764), .B2(KEYINPUT30), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n763), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n751), .A2(new_n762), .A3(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G1966), .ZN(new_n769));
  NOR2_X1   g344(.A1(G168), .A2(new_n685), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n685), .B2(G21), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n768), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(G5), .A2(G16), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G171), .B2(G16), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G1961), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n673), .A2(G35), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G162), .B2(new_n673), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT29), .B(G2090), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n673), .A2(G27), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G164), .B2(new_n673), .ZN(new_n782));
  INV_X1    g357(.A(G2078), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n750), .A2(new_n772), .A3(new_n780), .A4(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT24), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n673), .B1(new_n786), .B2(G34), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(KEYINPUT92), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(KEYINPUT92), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n786), .B2(G34), .ZN(new_n790));
  AOI22_X1  g365(.A1(G160), .A2(G29), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT93), .ZN(new_n792));
  INV_X1    g367(.A(G2084), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n785), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n685), .A2(G19), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n551), .B2(new_n685), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n797), .A2(G1341), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n771), .A2(new_n769), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT96), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n797), .A2(G1341), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n795), .A2(new_n798), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  OR3_X1    g377(.A1(new_n736), .A2(new_n737), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n737), .B1(new_n736), .B2(new_n802), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n707), .A2(new_n709), .B1(new_n803), .B2(new_n804), .ZN(G311));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  INV_X1    g381(.A(new_n709), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n708), .B1(new_n704), .B2(new_n705), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(G150));
  NAND2_X1  g384(.A1(new_n527), .A2(G55), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n811), .A2(new_n516), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT98), .B(G93), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n534), .A2(new_n813), .ZN(new_n814));
  AND3_X1   g389(.A1(new_n810), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(G860), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT101), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT37), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT100), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n594), .A2(G559), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n815), .A2(KEYINPUT99), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n815), .A2(KEYINPUT99), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n822), .B(new_n823), .C1(new_n550), .C2(new_n549), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n551), .A2(KEYINPUT99), .A3(new_n815), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(KEYINPUT38), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n826), .A2(KEYINPUT38), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n821), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n824), .A2(new_n825), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT38), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n833), .A2(G559), .A3(new_n594), .A4(new_n827), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n830), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT39), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n830), .A2(new_n834), .A3(KEYINPUT39), .ZN(new_n838));
  AND4_X1   g413(.A1(new_n820), .A2(new_n837), .A3(new_n816), .A4(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(G860), .B1(new_n835), .B2(new_n836), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n820), .B1(new_n840), .B2(new_n838), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n819), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(KEYINPUT102), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT102), .ZN(new_n844));
  OAI211_X1 g419(.A(new_n844), .B(new_n819), .C1(new_n839), .C2(new_n841), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(G145));
  XOR2_X1   g421(.A(new_n614), .B(G160), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(G162), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n849));
  NOR3_X1   g424(.A1(new_n472), .A2(KEYINPUT73), .A3(new_n489), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n491), .B1(new_n462), .B2(new_n493), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(KEYINPUT103), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n490), .A2(new_n494), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT103), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n854), .A2(new_n855), .A3(new_n849), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT104), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n505), .A2(new_n506), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n858), .B1(new_n505), .B2(new_n506), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n862), .A2(new_n756), .ZN(new_n863));
  INV_X1    g438(.A(new_n746), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n756), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n864), .B1(new_n863), .B2(new_n865), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n722), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT105), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g446(.A(KEYINPUT105), .B(new_n722), .C1(new_n867), .C2(new_n868), .ZN(new_n872));
  INV_X1    g447(.A(new_n868), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n873), .A2(new_n720), .A3(new_n866), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT106), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n873), .A2(KEYINPUT106), .A3(new_n720), .A4(new_n866), .ZN(new_n877));
  AOI22_X1  g452(.A1(new_n871), .A2(new_n872), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n479), .A2(G130), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n459), .A2(G118), .ZN(new_n880));
  OAI21_X1  g455(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n882), .B1(G142), .B2(new_n612), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n618), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n681), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n848), .B1(new_n878), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n871), .A2(new_n872), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n876), .A2(new_n877), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(new_n885), .ZN(new_n891));
  AOI21_X1  g466(.A(G37), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n878), .A2(new_n886), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT107), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n890), .A2(KEYINPUT107), .A3(new_n885), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(new_n848), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n892), .B(KEYINPUT40), .C1(new_n895), .C2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n900), .A2(new_n848), .A3(new_n896), .ZN(new_n901));
  AOI21_X1  g476(.A(KEYINPUT40), .B1(new_n901), .B2(new_n892), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n899), .A2(new_n902), .ZN(G395));
  XNOR2_X1  g478(.A(new_n831), .B(new_n602), .ZN(new_n904));
  INV_X1    g479(.A(G299), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n593), .B(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT41), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n602), .B(new_n826), .ZN(new_n909));
  INV_X1    g484(.A(new_n906), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT42), .ZN(new_n913));
  XOR2_X1   g488(.A(G303), .B(G288), .Z(new_n914));
  XNOR2_X1  g489(.A(G290), .B(new_n691), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n914), .B(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT42), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n908), .A2(new_n911), .A3(new_n918), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n913), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n917), .B1(new_n913), .B2(new_n919), .ZN(new_n921));
  OAI21_X1  g496(.A(G868), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n922), .B1(G868), .B2(new_n815), .ZN(G295));
  OAI21_X1  g498(.A(new_n922), .B1(G868), .B2(new_n815), .ZN(G331));
  XNOR2_X1  g499(.A(G301), .B(KEYINPUT108), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(G168), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n831), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n925), .B(G286), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n826), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n927), .A2(new_n906), .A3(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n926), .B(new_n826), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n930), .B1(new_n931), .B2(new_n907), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n917), .ZN(new_n933));
  INV_X1    g508(.A(G37), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n916), .B(new_n930), .C1(new_n931), .C2(new_n907), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n933), .A2(new_n938), .A3(new_n934), .A4(new_n935), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT109), .B1(new_n936), .B2(KEYINPUT43), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n937), .A2(KEYINPUT109), .A3(KEYINPUT44), .A4(new_n939), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(G397));
  OAI211_X1 g520(.A(new_n853), .B(new_n856), .C1(new_n860), .C2(new_n859), .ZN(new_n946));
  INV_X1    g521(.A(G1384), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT45), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G40), .ZN(new_n949));
  AOI211_X1 g524(.A(new_n949), .B(new_n465), .C1(new_n468), .C2(new_n475), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(KEYINPUT110), .ZN(new_n952));
  INV_X1    g527(.A(G1996), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n746), .B(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n756), .B(new_n761), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n681), .A2(new_n683), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n681), .A2(new_n683), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n954), .A2(new_n955), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(G290), .B(G1986), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n952), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  XOR2_X1   g535(.A(new_n960), .B(KEYINPUT111), .Z(new_n961));
  NAND3_X1  g536(.A1(new_n946), .A2(KEYINPUT45), .A3(new_n947), .ZN(new_n962));
  INV_X1    g537(.A(new_n465), .ZN(new_n963));
  INV_X1    g538(.A(new_n475), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT70), .B1(new_n474), .B2(G2105), .ZN(new_n965));
  OAI211_X1 g540(.A(G40), .B(new_n963), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n947), .B1(new_n496), .B2(new_n507), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n962), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n946), .A2(new_n947), .A3(new_n950), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(KEYINPUT58), .B(G1341), .ZN(new_n973));
  OAI22_X1  g548(.A1(new_n970), .A2(G1996), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n551), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT59), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n974), .A2(KEYINPUT59), .A3(new_n551), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G1956), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT50), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n981), .B1(new_n946), .B2(new_n947), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n950), .B1(KEYINPUT50), .B2(new_n968), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(KEYINPUT56), .B(G2072), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n962), .A2(new_n969), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  OR2_X1    g562(.A1(G299), .A2(KEYINPUT57), .ZN(new_n988));
  NAND2_X1  g563(.A1(G299), .A2(KEYINPUT57), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n984), .A2(new_n989), .A3(new_n988), .A4(new_n986), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT61), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n979), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT113), .ZN(new_n995));
  AOI22_X1  g570(.A1(new_n499), .A2(new_n504), .B1(new_n479), .B2(G126), .ZN(new_n996));
  AOI21_X1  g571(.A(G1384), .B1(new_n852), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n995), .B1(new_n997), .B2(new_n981), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n968), .A2(KEYINPUT113), .A3(KEYINPUT50), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n981), .B(new_n947), .C1(new_n857), .C2(new_n861), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1000), .A2(new_n950), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1348), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n1002), .A2(new_n1003), .B1(new_n972), .B2(new_n761), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT60), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT80), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n593), .B(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1004), .A2(new_n594), .A3(KEYINPUT60), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1008), .B(new_n1009), .C1(KEYINPUT60), .C2(new_n1004), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n991), .A2(KEYINPUT61), .A3(new_n992), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT124), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT124), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n991), .A2(new_n1013), .A3(KEYINPUT61), .A4(new_n992), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n994), .A2(new_n1010), .A3(new_n1012), .A4(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1016));
  AOI22_X1  g591(.A1(new_n984), .A2(new_n986), .B1(new_n989), .B2(new_n988), .ZN(new_n1017));
  OAI211_X1 g592(.A(KEYINPUT123), .B(new_n992), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n991), .B1(new_n1007), .B2(new_n1004), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT123), .B1(new_n1020), .B2(new_n992), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1015), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G8), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n968), .A2(new_n967), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n947), .B1(new_n857), .B2(new_n861), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n966), .B1(new_n1026), .B2(new_n967), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1025), .B1(new_n1027), .B2(KEYINPUT119), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT119), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1029), .B1(new_n948), .B2(new_n966), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1966), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  AOI221_X4 g606(.A(KEYINPUT103), .B1(new_n495), .B2(KEYINPUT4), .C1(new_n490), .C2(new_n494), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n855), .B1(new_n854), .B2(new_n849), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OR2_X1    g609(.A1(new_n859), .A2(new_n860), .ZN(new_n1035));
  AOI21_X1  g610(.A(G1384), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n966), .B1(new_n1036), .B2(new_n981), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1037), .A2(KEYINPUT120), .A3(new_n793), .A4(new_n1000), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1000), .A2(new_n1001), .A3(new_n793), .A4(new_n950), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT120), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1031), .A2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1024), .B1(new_n1043), .B2(G168), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n1039), .B(KEYINPUT120), .ZN(new_n1045));
  OAI211_X1 g620(.A(KEYINPUT119), .B(new_n950), .C1(new_n1036), .C2(KEYINPUT45), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1025), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1030), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n769), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1045), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT125), .B1(new_n1050), .B2(G8), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1044), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(G8), .B1(new_n1031), .B2(new_n1042), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT125), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1052), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(G286), .B1(new_n1031), .B2(new_n1042), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1045), .A2(new_n1049), .A3(G168), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n1058), .A3(G8), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1053), .A2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1028), .A2(KEYINPUT53), .A3(new_n783), .A4(new_n1030), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n962), .A2(new_n969), .A3(new_n783), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT126), .B(KEYINPUT53), .ZN(new_n1064));
  INV_X1    g639(.A(G1961), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n1063), .A2(new_n1064), .B1(new_n1002), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1062), .A2(G301), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1002), .A2(new_n1065), .ZN(new_n1069));
  INV_X1    g644(.A(new_n948), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n783), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1071));
  AOI211_X1 g646(.A(new_n1071), .B(new_n465), .C1(G2105), .C2(new_n474), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1070), .A2(new_n962), .A3(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1068), .A2(new_n1069), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(G171), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1067), .A2(new_n1075), .A3(KEYINPUT54), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n696), .A2(G1976), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n971), .A2(new_n1077), .A3(G8), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT52), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT114), .B(G1976), .Z(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT52), .B1(G288), .B2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n971), .A2(new_n1077), .A3(G8), .A4(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(G305), .A2(G1981), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G1981), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n572), .A2(new_n577), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT49), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1088), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1084), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT49), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1094), .A2(new_n1083), .A3(new_n1089), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1092), .A2(new_n1095), .A3(G8), .A4(new_n971), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1079), .A2(new_n1082), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(G303), .A2(G8), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n1098), .B(KEYINPUT55), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT112), .B(G1971), .Z(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n970), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(G2090), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1000), .A2(new_n1001), .A3(new_n1104), .A4(new_n950), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1024), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1097), .B1(new_n1100), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n966), .B1(new_n981), .B2(new_n997), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1108), .B(new_n1104), .C1(new_n1036), .C2(new_n981), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1024), .B1(new_n1103), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT118), .B1(new_n1110), .B2(new_n1100), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n982), .A2(G2090), .A3(new_n983), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1101), .B1(new_n962), .B2(new_n969), .ZN(new_n1113));
  OAI21_X1  g688(.A(G8), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT118), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1114), .A2(new_n1115), .A3(new_n1099), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1111), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1076), .A2(new_n1107), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1062), .A2(new_n1066), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(G171), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1066), .A2(G301), .A3(new_n1073), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT54), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1023), .A2(new_n1061), .A3(new_n1123), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1110), .A2(KEYINPUT118), .A3(new_n1100), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1115), .B1(new_n1114), .B2(new_n1099), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1107), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  OAI211_X1 g702(.A(G8), .B(G168), .C1(new_n1031), .C2(new_n1042), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT121), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1128), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1130), .A2(new_n1131), .A3(new_n1107), .A4(new_n1117), .ZN(new_n1132));
  XOR2_X1   g707(.A(KEYINPUT122), .B(KEYINPUT63), .Z(new_n1133));
  NAND3_X1  g708(.A1(new_n1129), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1106), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n1099), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1130), .A2(KEYINPUT63), .A3(new_n1107), .A4(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1135), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1096), .ZN(new_n1140));
  NOR2_X1   g715(.A1(G288), .A2(G1976), .ZN(new_n1141));
  XOR2_X1   g716(.A(new_n1141), .B(KEYINPUT117), .Z(new_n1142));
  OAI21_X1  g717(.A(new_n1086), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n971), .A2(G8), .ZN(new_n1144));
  XOR2_X1   g719(.A(new_n1144), .B(KEYINPUT116), .Z(new_n1145));
  AOI21_X1  g720(.A(new_n1139), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1124), .A2(new_n1138), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1053), .A2(new_n1060), .A3(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1127), .A2(new_n1120), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1148), .B1(new_n1053), .B2(new_n1060), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n961), .B1(new_n1147), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n952), .A2(new_n953), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT46), .ZN(new_n1156));
  INV_X1    g731(.A(new_n955), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n952), .B1(new_n746), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n1159), .B(KEYINPUT47), .Z(new_n1160));
  NOR2_X1   g735(.A1(G290), .A2(G1986), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n952), .A2(new_n1161), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n1162), .A2(KEYINPUT48), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1162), .A2(KEYINPUT48), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n952), .A2(new_n958), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n954), .A2(new_n955), .ZN(new_n1167));
  OAI22_X1  g742(.A1(new_n1167), .A2(new_n956), .B1(G2067), .B2(new_n756), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n952), .A2(new_n1168), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n1160), .A2(new_n1166), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1154), .A2(new_n1170), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g746(.A1(new_n901), .A2(new_n892), .ZN(new_n1173));
  INV_X1    g747(.A(G227), .ZN(new_n1174));
  NAND2_X1  g748(.A1(new_n1174), .A2(G319), .ZN(new_n1175));
  XOR2_X1   g749(.A(new_n1175), .B(KEYINPUT127), .Z(new_n1176));
  NOR3_X1   g750(.A1(G229), .A2(G401), .A3(new_n1176), .ZN(new_n1177));
  NAND3_X1  g751(.A1(new_n1173), .A2(new_n940), .A3(new_n1177), .ZN(G225));
  INV_X1    g752(.A(G225), .ZN(G308));
endmodule


