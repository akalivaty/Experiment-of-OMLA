//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1335, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1409, new_n1410, new_n1411, new_n1412, new_n1413;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n205), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n212), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OR2_X1    g0024(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(KEYINPUT64), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g0028(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n231), .A2(new_n210), .ZN(new_n232));
  INV_X1    g0032(.A(new_n201), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G50), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g0036(.A1(new_n215), .A2(new_n225), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g0037(.A(new_n237), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(G226), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT67), .ZN(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G50), .B(G58), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(KEYINPUT66), .ZN(new_n253));
  XOR2_X1   g0053(.A(G68), .B(G77), .Z(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n251), .B(new_n255), .ZN(G351));
  XNOR2_X1  g0056(.A(KEYINPUT3), .B(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(G222), .A3(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G77), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(G1698), .ZN(new_n261));
  INV_X1    g0061(.A(G223), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n259), .B1(new_n260), .B2(new_n257), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n230), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n268));
  INV_X1    g0068(.A(G274), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n264), .A2(G1), .A3(G13), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n268), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n270), .B1(new_n273), .B2(G226), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n267), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G179), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n278), .B(KEYINPUT68), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  AND3_X1   g0080(.A1(new_n228), .A2(new_n229), .A3(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G58), .ZN(new_n282));
  OR2_X1    g0082(.A1(new_n282), .A2(KEYINPUT8), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(KEYINPUT8), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(new_n210), .A3(G33), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n281), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n202), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n281), .B1(G1), .B2(new_n210), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n292), .B1(new_n293), .B2(new_n202), .ZN(new_n294));
  OAI22_X1  g0094(.A1(new_n276), .A2(G169), .B1(new_n289), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n279), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n294), .A2(new_n289), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT69), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n297), .B(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT9), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n297), .B(KEYINPUT69), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT9), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G190), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n275), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n305), .B1(G200), .B2(new_n275), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n300), .A2(new_n303), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT10), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT10), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n300), .A2(new_n303), .A3(new_n309), .A4(new_n306), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n296), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G68), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G20), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n210), .A2(G33), .ZN(new_n314));
  INV_X1    g0114(.A(new_n287), .ZN(new_n315));
  OAI221_X1 g0115(.A(new_n313), .B1(new_n314), .B2(new_n260), .C1(new_n315), .C2(new_n202), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n228), .A2(new_n229), .A3(new_n280), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT11), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G13), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n321), .A2(G1), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n323), .A2(new_n313), .ZN(new_n324));
  XOR2_X1   g0124(.A(new_n324), .B(KEYINPUT12), .Z(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(new_n312), .B2(new_n293), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n320), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n257), .A2(G226), .A3(new_n258), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT70), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT70), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n257), .A2(new_n331), .A3(G226), .A4(new_n258), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(G33), .A2(G97), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n257), .A2(G232), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n334), .B1(new_n335), .B2(new_n258), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n265), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n270), .B1(new_n273), .B2(G238), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(KEYINPUT13), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT13), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n336), .B1(new_n332), .B2(new_n330), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n342), .B(new_n339), .C1(new_n343), .C2(new_n265), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT71), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT14), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n345), .A2(new_n346), .A3(new_n347), .A4(G169), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n341), .A2(G179), .A3(new_n344), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G169), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n351), .B1(KEYINPUT71), .B2(KEYINPUT14), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n345), .A2(new_n352), .B1(new_n346), .B2(new_n347), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n328), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G200), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n345), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n341), .A2(new_n304), .A3(new_n344), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n328), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  MUX2_X1   g0159(.A(new_n290), .B(new_n293), .S(G77), .Z(new_n360));
  INV_X1    g0160(.A(new_n285), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n361), .A2(new_n315), .ZN(new_n362));
  XNOR2_X1  g0162(.A(KEYINPUT15), .B(G87), .ZN(new_n363));
  OAI22_X1  g0163(.A1(new_n363), .A2(new_n314), .B1(new_n210), .B2(new_n260), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n317), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n257), .A2(G232), .A3(new_n258), .ZN(new_n367));
  INV_X1    g0167(.A(G238), .ZN(new_n368));
  OAI221_X1 g0168(.A(new_n367), .B1(new_n206), .B2(new_n257), .C1(new_n261), .C2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n266), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n270), .B1(new_n273), .B2(G244), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n372), .A2(new_n277), .ZN(new_n373));
  INV_X1    g0173(.A(new_n371), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n374), .B1(new_n369), .B2(new_n266), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n375), .A2(new_n351), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n366), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n372), .A2(new_n355), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n375), .A2(new_n304), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n366), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n311), .A2(new_n354), .A3(new_n359), .A4(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n285), .A2(new_n291), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n293), .B2(new_n285), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  OR2_X1    g0186(.A1(KEYINPUT72), .A2(KEYINPUT3), .ZN(new_n387));
  NAND2_X1  g0187(.A1(KEYINPUT72), .A2(KEYINPUT3), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n387), .A2(G33), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G33), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT3), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G226), .A2(G1698), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n262), .B2(G1698), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n389), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(G33), .A2(G87), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n265), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n270), .ZN(new_n397));
  INV_X1    g0197(.A(G232), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n397), .B1(new_n272), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n304), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n355), .B1(new_n396), .B2(new_n399), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT16), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n282), .A2(new_n312), .ZN(new_n405));
  OAI21_X1  g0205(.A(G20), .B1(new_n405), .B2(new_n201), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n287), .A2(G159), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(G20), .B1(new_n389), .B2(new_n391), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT73), .B1(new_n409), .B2(KEYINPUT7), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT73), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT7), .ZN(new_n412));
  INV_X1    g0212(.A(new_n391), .ZN(new_n413));
  AND2_X1   g0213(.A1(KEYINPUT72), .A2(KEYINPUT3), .ZN(new_n414));
  NOR2_X1   g0214(.A1(KEYINPUT72), .A2(KEYINPUT3), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n413), .B1(new_n416), .B2(G33), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n411), .B(new_n412), .C1(new_n417), .C2(G20), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n409), .A2(KEYINPUT7), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n410), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  AOI211_X1 g0220(.A(new_n404), .B(new_n408), .C1(new_n420), .C2(G68), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n412), .B1(new_n257), .B2(G20), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT3), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(G33), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n387), .A2(new_n388), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n425), .B1(new_n426), .B2(new_n390), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n210), .A2(KEYINPUT7), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n422), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n408), .B1(new_n429), .B2(G68), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n317), .B1(new_n430), .B2(KEYINPUT16), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n386), .B(new_n403), .C1(new_n421), .C2(new_n431), .ZN(new_n432));
  XNOR2_X1  g0232(.A(new_n432), .B(KEYINPUT17), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT18), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n420), .A2(G68), .ZN(new_n435));
  INV_X1    g0235(.A(new_n408), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(KEYINPUT16), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n431), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n385), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n400), .A2(G169), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n440), .B1(new_n277), .B2(new_n400), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n434), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n386), .B1(new_n421), .B2(new_n431), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n444), .A2(KEYINPUT18), .A3(new_n441), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n433), .A2(new_n446), .ZN(new_n447));
  OR3_X1    g0247(.A1(new_n383), .A2(KEYINPUT74), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT74), .B1(new_n383), .B2(new_n447), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n363), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(new_n290), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n290), .B1(G1), .B2(new_n390), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n317), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n451), .ZN(new_n456));
  NOR2_X1   g0256(.A1(G87), .A2(G97), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n457), .A2(new_n206), .B1(new_n334), .B2(new_n210), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT19), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n210), .ZN(new_n460));
  OAI22_X1  g0260(.A1(new_n458), .A2(new_n459), .B1(new_n334), .B2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n389), .A2(new_n210), .A3(G68), .A4(new_n391), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n453), .B(new_n456), .C1(new_n463), .C2(new_n281), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT78), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n389), .A2(G244), .A3(G1698), .A4(new_n391), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G116), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n368), .A2(G1698), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n389), .A2(new_n391), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n466), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n266), .ZN(new_n471));
  INV_X1    g0271(.A(G45), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n472), .A2(new_n269), .A3(G1), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n218), .B1(new_n209), .B2(G45), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n271), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n351), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n281), .B1(new_n461), .B2(new_n462), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(new_n452), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT78), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(new_n480), .A3(new_n456), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n471), .A2(new_n277), .A3(new_n475), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n465), .A2(new_n477), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n471), .A2(G190), .A3(new_n475), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n317), .A2(new_n454), .A3(new_n217), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n478), .A2(new_n452), .A3(new_n485), .ZN(new_n486));
  OR2_X1    g0286(.A1(new_n473), .A2(new_n474), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n470), .A2(new_n266), .B1(new_n271), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n484), .B(new_n486), .C1(new_n355), .C2(new_n488), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n483), .A2(KEYINPUT79), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(KEYINPUT79), .B1(new_n483), .B2(new_n489), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n290), .A2(G97), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n493), .B1(new_n455), .B2(G97), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G97), .A2(G107), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n207), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT75), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT6), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n207), .A2(new_n498), .A3(new_n499), .A4(new_n496), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n205), .A2(KEYINPUT6), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n501), .A2(G20), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n287), .A2(G77), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n390), .B1(new_n414), .B2(new_n415), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n428), .B1(new_n506), .B2(new_n424), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n391), .A2(new_n424), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT7), .B1(new_n508), .B2(new_n210), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n504), .B(new_n505), .C1(new_n510), .C2(new_n206), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n495), .B1(new_n511), .B2(new_n317), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n472), .A2(G1), .ZN(new_n513));
  AND2_X1   g0313(.A1(KEYINPUT5), .A2(G41), .ZN(new_n514));
  NOR2_X1   g0314(.A1(KEYINPUT5), .A2(G41), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(new_n271), .A3(G257), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n513), .B(G274), .C1(new_n515), .C2(new_n514), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n517), .A2(KEYINPUT77), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT77), .B1(new_n517), .B2(new_n518), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g0321(.A1(KEYINPUT4), .A2(G244), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n257), .A2(new_n258), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G283), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT76), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT76), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n526), .A2(G33), .A3(G283), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n391), .A2(new_n424), .A3(G250), .A4(G1698), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n523), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n389), .A2(G244), .A3(new_n258), .A4(new_n391), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT4), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n265), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(G200), .B1(new_n521), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n530), .A2(new_n533), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n266), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n517), .A2(new_n518), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(G190), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n512), .A2(new_n535), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(G33), .B1(new_n387), .B2(new_n388), .ZN(new_n542));
  OAI211_X1 g0342(.A(KEYINPUT7), .B(new_n210), .C1(new_n542), .C2(new_n425), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n206), .B1(new_n543), .B2(new_n422), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n504), .A2(new_n505), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n317), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n494), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT77), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n538), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n517), .A2(KEYINPUT77), .A3(new_n518), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n537), .A2(new_n551), .A3(new_n277), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n351), .B1(new_n534), .B2(new_n538), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n547), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n541), .A2(new_n554), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n516), .A2(new_n271), .A3(G264), .ZN(new_n556));
  NAND2_X1  g0356(.A1(G257), .A2(G1698), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n218), .B2(G1698), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n389), .A2(new_n391), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(G33), .A2(G294), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n556), .B1(new_n561), .B2(new_n266), .ZN(new_n562));
  AOI21_X1  g0362(.A(G169), .B1(new_n562), .B2(new_n518), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n265), .B1(new_n559), .B2(new_n560), .ZN(new_n564));
  INV_X1    g0364(.A(new_n518), .ZN(new_n565));
  NOR4_X1   g0365(.A1(new_n564), .A2(new_n556), .A3(G179), .A4(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT86), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n562), .A2(new_n277), .A3(new_n518), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT86), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n564), .A2(new_n565), .A3(new_n556), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n568), .B(new_n569), .C1(G169), .C2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT22), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n573), .A2(new_n217), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n389), .A2(new_n210), .A3(new_n391), .A4(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n210), .A2(G87), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n573), .B1(new_n508), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n467), .A2(G20), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT23), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n210), .B2(G107), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n578), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n575), .A2(new_n577), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n583), .A2(KEYINPUT85), .A3(KEYINPUT24), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT24), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n575), .A2(new_n577), .A3(new_n585), .A4(new_n582), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(KEYINPUT85), .B1(new_n583), .B2(KEYINPUT24), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n317), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n322), .A2(G20), .A3(new_n206), .ZN(new_n590));
  XNOR2_X1  g0390(.A(new_n590), .B(KEYINPUT25), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(G107), .B2(new_n455), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n572), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n562), .A2(new_n304), .A3(new_n518), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n570), .B2(G200), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n589), .A2(new_n596), .A3(new_n592), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n555), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n516), .A2(new_n271), .A3(G270), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n518), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT80), .ZN(new_n601));
  NAND2_X1  g0401(.A1(G264), .A2(G1698), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n219), .B2(G1698), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n389), .A2(new_n391), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n508), .A2(G303), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n266), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT80), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n599), .A2(new_n608), .A3(new_n518), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n601), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  OR2_X1    g0410(.A1(new_n610), .A2(G190), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n355), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT81), .B1(new_n455), .B2(G116), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT81), .ZN(new_n615));
  INV_X1    g0415(.A(G116), .ZN(new_n616));
  NOR4_X1   g0416(.A1(new_n317), .A2(new_n454), .A3(new_n615), .A4(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n210), .A2(G116), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  OAI22_X1  g0419(.A1(new_n614), .A2(new_n617), .B1(new_n323), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT20), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n317), .A2(new_n619), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n210), .B1(new_n205), .B2(G33), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n623), .B1(new_n525), .B2(new_n527), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n621), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT83), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI211_X1 g0427(.A(KEYINPUT83), .B(new_n621), .C1(new_n622), .C2(new_n624), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n622), .ZN(new_n630));
  INV_X1    g0430(.A(new_n623), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n528), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n630), .A2(KEYINPUT82), .A3(KEYINPUT20), .A4(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n632), .A2(KEYINPUT20), .A3(new_n317), .A4(new_n619), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT82), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n620), .B1(new_n629), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n613), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(KEYINPUT84), .A2(KEYINPUT21), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n610), .A2(G169), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n640), .B1(new_n638), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n620), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n627), .A2(new_n633), .A3(new_n636), .A4(new_n628), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n610), .A2(G169), .ZN(new_n646));
  INV_X1    g0446(.A(new_n640), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n601), .A2(new_n607), .A3(G179), .A4(new_n609), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n639), .A2(new_n642), .A3(new_n648), .A4(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n598), .A2(new_n652), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n450), .A2(new_n492), .A3(new_n653), .ZN(G372));
  INV_X1    g0454(.A(KEYINPUT87), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n487), .A2(new_n655), .A3(new_n271), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n475), .A2(KEYINPUT87), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n470), .A2(new_n266), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n482), .B(new_n464), .C1(G169), .C2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n547), .A2(new_n552), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n484), .B(new_n486), .C1(new_n355), .C2(new_n658), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n660), .A2(new_n553), .A3(new_n661), .A4(new_n659), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n659), .B1(new_n662), .B2(KEYINPUT26), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n568), .B1(G169), .B2(new_n570), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n664), .B1(new_n589), .B2(new_n592), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n666), .A2(new_n642), .A3(new_n648), .A4(new_n651), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n541), .A2(new_n554), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n589), .A2(new_n596), .A3(new_n592), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n661), .A2(new_n659), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n663), .B1(new_n667), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n483), .A2(new_n489), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT79), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n483), .A2(KEYINPUT79), .A3(new_n489), .ZN(new_n676));
  INV_X1    g0476(.A(new_n554), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(KEYINPUT26), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n672), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n450), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n345), .A2(new_n352), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n346), .A2(new_n347), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n684), .A2(new_n348), .A3(new_n349), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n685), .A2(new_n328), .B1(new_n359), .B2(new_n378), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT17), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n432), .B(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT88), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n439), .B2(new_n442), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n444), .A2(KEYINPUT88), .A3(new_n441), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n690), .A2(new_n691), .A3(KEYINPUT18), .ZN(new_n692));
  AOI21_X1  g0492(.A(KEYINPUT18), .B1(new_n690), .B2(new_n691), .ZN(new_n693));
  OAI22_X1  g0493(.A1(new_n686), .A2(new_n688), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n308), .A2(new_n310), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n296), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n681), .A2(new_n696), .ZN(G369));
  NAND3_X1  g0497(.A1(new_n642), .A2(new_n648), .A3(new_n651), .ZN(new_n698));
  OR3_X1    g0498(.A1(new_n323), .A2(KEYINPUT27), .A3(G20), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT27), .B1(new_n323), .B2(G20), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(G213), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G343), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n645), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n698), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n652), .B2(new_n704), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G330), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n593), .A2(new_n703), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n594), .A2(new_n597), .A3(new_n708), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n567), .A2(new_n571), .B1(new_n589), .B2(new_n592), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n703), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n707), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n703), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n698), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n709), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n666), .A2(new_n703), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n713), .A2(new_n718), .ZN(G399));
  INV_X1    g0519(.A(new_n213), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(G41), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n457), .A2(new_n206), .A3(new_n616), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n721), .A2(new_n722), .A3(new_n209), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n723), .B1(new_n235), .B2(new_n721), .ZN(new_n724));
  XOR2_X1   g0524(.A(new_n724), .B(KEYINPUT89), .Z(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT28), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT93), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n710), .A2(new_n668), .A3(new_n669), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n648), .A2(new_n651), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n645), .B1(new_n611), .B2(new_n612), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n647), .B1(new_n645), .B2(new_n646), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n728), .A2(new_n492), .A3(new_n732), .A4(new_n714), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(KEYINPUT92), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT92), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n653), .A2(new_n735), .A3(new_n492), .A4(new_n714), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n488), .A2(new_n562), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(new_n649), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n534), .A2(new_n538), .ZN(new_n740));
  AOI21_X1  g0540(.A(KEYINPUT30), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n739), .A2(KEYINPUT30), .A3(new_n740), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n537), .A2(new_n551), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n570), .A2(G179), .ZN(new_n745));
  INV_X1    g0545(.A(new_n658), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n744), .A2(new_n745), .A3(new_n610), .A4(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n742), .A2(new_n743), .A3(new_n747), .ZN(new_n748));
  XOR2_X1   g0548(.A(KEYINPUT90), .B(KEYINPUT31), .Z(new_n749));
  NOR2_X1   g0549(.A1(new_n714), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n743), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n741), .ZN(new_n753));
  AND2_X1   g0553(.A1(new_n746), .A2(new_n610), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n754), .A2(KEYINPUT91), .A3(new_n744), .A4(new_n745), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT91), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n747), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n714), .B1(new_n753), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n751), .B1(new_n759), .B2(KEYINPUT31), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n737), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n727), .B1(new_n762), .B2(G330), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n760), .B1(new_n734), .B2(new_n736), .ZN(new_n764));
  INV_X1    g0564(.A(G330), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n764), .A2(KEYINPUT93), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(KEYINPUT26), .B1(new_n670), .B2(new_n554), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n659), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n594), .A2(new_n642), .A3(new_n648), .A4(new_n651), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n769), .B1(new_n671), .B2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT26), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n675), .A2(new_n677), .A3(new_n772), .A4(new_n676), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n703), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(KEYINPUT29), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n703), .B1(new_n672), .B2(new_n679), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n775), .B1(KEYINPUT29), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n767), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n726), .B1(new_n779), .B2(G1), .ZN(G364));
  XNOR2_X1  g0580(.A(new_n707), .B(KEYINPUT94), .ZN(new_n781));
  INV_X1    g0581(.A(new_n721), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n321), .A2(G20), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G45), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n782), .A2(G1), .A3(new_n784), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n785), .A2(KEYINPUT95), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(KEYINPUT95), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n781), .B(new_n788), .C1(G330), .C2(new_n706), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n231), .B1(G20), .B2(new_n351), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n255), .A2(new_n472), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n720), .A2(new_n417), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n798), .B1(new_n472), .B2(new_n235), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n796), .B1(new_n800), .B2(KEYINPUT97), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n801), .B1(KEYINPUT97), .B2(new_n800), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n720), .A2(new_n508), .ZN(new_n803));
  XNOR2_X1  g0603(.A(G355), .B(KEYINPUT96), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n803), .A2(new_n804), .B1(new_n616), .B2(new_n720), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n795), .B1(new_n802), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n790), .ZN(new_n807));
  NAND2_X1  g0607(.A1(G20), .A2(G190), .ZN(new_n808));
  NOR3_X1   g0608(.A1(new_n808), .A2(new_n355), .A3(G179), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n210), .A2(G190), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NOR3_X1   g0612(.A1(new_n812), .A2(G179), .A3(new_n355), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n257), .B1(new_n217), .B2(new_n810), .C1(new_n814), .C2(new_n206), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT99), .Z(new_n816));
  NOR2_X1   g0616(.A1(new_n277), .A2(new_n355), .ZN(new_n817));
  INV_X1    g0617(.A(new_n808), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n817), .A2(new_n811), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n819), .A2(new_n202), .B1(new_n820), .B2(new_n312), .ZN(new_n821));
  NOR2_X1   g0621(.A1(G179), .A2(G200), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(G190), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(G20), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(new_n205), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n811), .A2(G179), .A3(new_n355), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NOR3_X1   g0628(.A1(new_n808), .A2(new_n277), .A3(G200), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n828), .A2(G77), .B1(new_n829), .B2(G58), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n821), .B(new_n826), .C1(KEYINPUT98), .C2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n830), .A2(KEYINPUT98), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT32), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n811), .A2(new_n822), .ZN(new_n834));
  INV_X1    g0634(.A(G159), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n834), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n837), .A2(KEYINPUT32), .A3(G159), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n832), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n816), .A2(new_n831), .A3(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(G283), .ZN(new_n841));
  INV_X1    g0641(.A(G303), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n814), .A2(new_n841), .B1(new_n842), .B2(new_n810), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n257), .B(new_n843), .C1(G322), .C2(new_n829), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n824), .A2(G294), .ZN(new_n845));
  OR2_X1    g0645(.A1(new_n834), .A2(KEYINPUT100), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n834), .A2(KEYINPUT100), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(G329), .ZN(new_n850));
  INV_X1    g0650(.A(new_n820), .ZN(new_n851));
  NOR2_X1   g0651(.A1(KEYINPUT33), .A2(G317), .ZN(new_n852));
  AND2_X1   g0652(.A1(KEYINPUT33), .A2(G317), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(G311), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n854), .B1(new_n855), .B2(new_n827), .ZN(new_n856));
  INV_X1    g0656(.A(new_n819), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n856), .B1(G326), .B2(new_n857), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n844), .A2(new_n845), .A3(new_n850), .A4(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n807), .B1(new_n840), .B2(new_n859), .ZN(new_n860));
  NOR3_X1   g0660(.A1(new_n806), .A2(new_n860), .A3(new_n788), .ZN(new_n861));
  INV_X1    g0661(.A(new_n793), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n861), .B1(new_n706), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n789), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT101), .ZN(G396));
  AOI21_X1  g0665(.A(new_n714), .B1(new_n360), .B2(new_n365), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n377), .B1(new_n381), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT104), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n366), .B(new_n714), .C1(new_n373), .C2(new_n376), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n868), .B1(new_n867), .B2(new_n869), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n776), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n659), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n670), .A2(new_n554), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n874), .B1(new_n875), .B2(new_n772), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n729), .A2(new_n731), .A3(new_n665), .ZN(new_n877));
  INV_X1    g0677(.A(new_n670), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n555), .A2(new_n597), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n876), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n772), .B1(new_n492), .B2(new_n677), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n872), .B(new_n714), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n873), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n767), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n762), .A2(new_n727), .A3(G330), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT93), .B1(new_n764), .B2(new_n765), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n887), .A2(new_n873), .A3(new_n882), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n884), .A2(new_n888), .A3(new_n788), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n790), .A2(new_n791), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n788), .B1(new_n260), .B2(new_n890), .ZN(new_n891));
  XOR2_X1   g0691(.A(KEYINPUT102), .B(G283), .Z(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n893), .A2(new_n851), .B1(G107), .B2(new_n809), .ZN(new_n894));
  OAI221_X1 g0694(.A(new_n894), .B1(new_n842), .B2(new_n819), .C1(new_n848), .C2(new_n855), .ZN(new_n895));
  INV_X1    g0695(.A(new_n829), .ZN(new_n896));
  INV_X1    g0696(.A(G294), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n508), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n813), .A2(G87), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n616), .B2(new_n827), .ZN(new_n900));
  NOR4_X1   g0700(.A1(new_n895), .A2(new_n826), .A3(new_n898), .A4(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n814), .A2(new_n312), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(G50), .B2(new_n809), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n903), .B(new_n417), .C1(new_n282), .C2(new_n825), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(G132), .B2(new_n849), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT103), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n851), .A2(G150), .B1(G143), .B2(new_n829), .ZN(new_n907));
  INV_X1    g0707(.A(G137), .ZN(new_n908));
  OAI221_X1 g0708(.A(new_n907), .B1(new_n908), .B2(new_n819), .C1(new_n835), .C2(new_n827), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(KEYINPUT34), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n901), .B1(new_n906), .B2(new_n910), .ZN(new_n911));
  OAI221_X1 g0711(.A(new_n891), .B1(new_n872), .B2(new_n792), .C1(new_n807), .C2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n889), .A2(new_n912), .ZN(G384));
  NOR2_X1   g0713(.A1(new_n783), .A2(new_n209), .ZN(new_n914));
  INV_X1    g0714(.A(new_n749), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n759), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(KEYINPUT31), .B2(new_n759), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n737), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n328), .A2(new_n703), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n354), .A2(new_n359), .A3(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n328), .B(new_n703), .C1(new_n685), .C2(new_n358), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n872), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n918), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n408), .B1(new_n420), .B2(G68), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n281), .B1(new_n926), .B2(KEYINPUT16), .ZN(new_n927));
  AOI211_X1 g0727(.A(new_n412), .B(G20), .C1(new_n389), .C2(new_n391), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n412), .B1(new_n417), .B2(G20), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n928), .B1(new_n929), .B2(KEYINPUT73), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n312), .B1(new_n930), .B2(new_n418), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n404), .B1(new_n931), .B2(new_n408), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n385), .B1(new_n927), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n933), .A2(new_n701), .ZN(new_n934));
  INV_X1    g0734(.A(new_n446), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n934), .B1(new_n935), .B2(new_n688), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n432), .B1(new_n439), .B2(new_n701), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT37), .B1(new_n444), .B2(new_n441), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n701), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n441), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n432), .B1(new_n933), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(KEYINPUT37), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n936), .A2(new_n945), .A3(KEYINPUT38), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT38), .ZN(new_n947));
  INV_X1    g0747(.A(new_n934), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(new_n433), .B2(new_n446), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n938), .A2(new_n939), .B1(new_n943), .B2(KEYINPUT37), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n946), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n925), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT40), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n433), .B1(new_n692), .B2(new_n693), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n439), .A2(new_n701), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n439), .A2(new_n442), .A3(new_n689), .ZN(new_n958));
  AOI21_X1  g0758(.A(KEYINPUT88), .B1(new_n444), .B2(new_n441), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(KEYINPUT37), .B1(new_n960), .B2(new_n937), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n956), .A2(new_n957), .B1(new_n961), .B2(new_n940), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n946), .B1(new_n962), .B2(KEYINPUT38), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n925), .A2(KEYINPUT40), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n955), .A2(new_n964), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n450), .A2(new_n918), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n965), .B(new_n966), .Z(new_n967));
  NOR2_X1   g0767(.A1(new_n967), .A2(new_n765), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n922), .B1(new_n882), .B2(new_n869), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n952), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n434), .B1(new_n958), .B2(new_n959), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n690), .A2(new_n691), .A3(KEYINPUT18), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n972), .A2(new_n973), .A3(new_n701), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT106), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT39), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n978), .B(new_n946), .C1(new_n962), .C2(KEYINPUT38), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n952), .A2(KEYINPUT39), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n685), .A2(new_n328), .A3(new_n714), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n971), .A2(KEYINPUT106), .A3(new_n974), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n977), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n450), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n696), .B1(new_n987), .B2(new_n777), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n986), .B(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n914), .B1(new_n969), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n989), .B2(new_n969), .ZN(new_n991));
  NOR3_X1   g0791(.A1(new_n234), .A2(new_n260), .A3(new_n405), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n312), .A2(G50), .ZN(new_n993));
  OAI211_X1 g0793(.A(G1), .B(new_n321), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT105), .Z(new_n996));
  OR2_X1    g0796(.A1(new_n996), .A2(KEYINPUT35), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(KEYINPUT35), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n997), .A2(G116), .A3(new_n232), .A4(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT36), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n991), .A2(new_n994), .A3(new_n1000), .ZN(G367));
  NOR2_X1   g0801(.A1(new_n714), .A2(new_n486), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n659), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n878), .B2(new_n1002), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT43), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n512), .A2(new_n714), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n668), .A2(new_n1007), .B1(new_n554), .B2(new_n714), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT107), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n554), .B1(new_n1009), .B2(new_n594), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT108), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1012), .A2(new_n714), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n716), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1009), .A2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT42), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1006), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1018), .B(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n713), .A2(new_n1009), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1020), .B(new_n1021), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n721), .B(KEYINPUT41), .Z(new_n1023));
  INV_X1    g0823(.A(KEYINPUT44), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1009), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1024), .B1(new_n1025), .B2(new_n718), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(KEYINPUT110), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n716), .A2(new_n717), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1028), .A2(KEYINPUT44), .A3(new_n1009), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(KEYINPUT109), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT110), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1031), .B(new_n1024), .C1(new_n1025), .C2(new_n718), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT109), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1028), .A2(new_n1033), .A3(KEYINPUT44), .A4(new_n1009), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1027), .A2(new_n1030), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1028), .A2(new_n1009), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT45), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n713), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1035), .A2(new_n1037), .A3(new_n713), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n712), .A2(new_n715), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n1015), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n707), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n781), .B2(new_n1045), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n767), .A2(new_n777), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(KEYINPUT111), .B1(new_n1042), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1048), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT111), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1050), .A2(new_n1051), .A3(new_n1041), .A4(new_n1040), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1023), .B1(new_n1053), .B2(new_n779), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n784), .A2(G1), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1022), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n814), .A2(new_n260), .B1(new_n834), .B2(new_n908), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n508), .B(new_n1057), .C1(G58), .C2(new_n809), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n828), .A2(G50), .B1(new_n851), .B2(G159), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n857), .A2(G143), .B1(G150), .B2(new_n829), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n824), .A2(G68), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n810), .A2(new_n616), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1063), .A2(KEYINPUT46), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT112), .Z(new_n1065));
  NOR2_X1   g0865(.A1(new_n819), .A2(new_n855), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n417), .B(new_n1066), .C1(G97), .C2(new_n813), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n851), .A2(G294), .B1(new_n837), .B2(G317), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n893), .A2(new_n828), .B1(G303), .B2(new_n829), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1063), .A2(KEYINPUT46), .B1(G107), .B2(new_n824), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1062), .B1(new_n1065), .B2(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n807), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n788), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1004), .A2(new_n793), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n797), .A2(new_n246), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1078), .B(new_n794), .C1(new_n213), .C2(new_n363), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1056), .A2(new_n1080), .ZN(G387));
  INV_X1    g0881(.A(KEYINPUT116), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1047), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n778), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1084), .A2(new_n1048), .A3(new_n721), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n803), .A2(new_n722), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(G107), .B2(new_n213), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n243), .A2(G45), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n285), .A2(new_n202), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT50), .Z(new_n1090));
  AOI211_X1 g0890(.A(G45), .B(new_n722), .C1(G68), .C2(G77), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n798), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1087), .B1(new_n1088), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1076), .B1(new_n1093), .B2(new_n795), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n893), .A2(new_n824), .B1(G294), .B2(new_n809), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(G303), .A2(new_n828), .B1(new_n857), .B2(G322), .ZN(new_n1096));
  INV_X1    g0896(.A(G317), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n1096), .B1(new_n855), .B2(new_n820), .C1(new_n1097), .C2(new_n896), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT48), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1095), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(new_n1099), .B2(new_n1098), .ZN(new_n1101));
  OR2_X1    g0901(.A1(new_n1101), .A2(KEYINPUT49), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n417), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(KEYINPUT49), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n813), .A2(G116), .B1(G326), .B2(new_n837), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n814), .A2(new_n205), .B1(new_n835), .B2(new_n819), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n809), .A2(G77), .ZN(new_n1108));
  INV_X1    g0908(.A(G150), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n1108), .B1(new_n834), .B2(new_n1109), .C1(new_n896), .C2(new_n202), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n361), .A2(new_n820), .B1(new_n827), .B2(new_n312), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n451), .A2(new_n824), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n417), .ZN(new_n1113));
  NOR4_X1   g0913(.A1(new_n1107), .A2(new_n1110), .A3(new_n1111), .A4(new_n1113), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT114), .Z(new_n1115));
  AOI21_X1  g0915(.A(new_n807), .B1(new_n1106), .B2(new_n1115), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1094), .B(new_n1116), .C1(new_n712), .C2(new_n793), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT115), .Z(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n1047), .B2(new_n1055), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1082), .B1(new_n1085), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1085), .A2(new_n1082), .A3(new_n1119), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(G393));
  AOI21_X1  g0923(.A(new_n782), .B1(new_n1042), .B2(new_n1048), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n1053), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n508), .B1(new_n814), .B2(new_n206), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(G116), .B2(new_n824), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n896), .A2(new_n855), .B1(new_n819), .B2(new_n1097), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT52), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n851), .A2(G303), .B1(new_n837), .B2(G322), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n809), .A2(new_n893), .B1(new_n828), .B2(G294), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1127), .A2(new_n1129), .A3(new_n1130), .A4(new_n1131), .ZN(new_n1132));
  XOR2_X1   g0932(.A(new_n1132), .B(KEYINPUT118), .Z(new_n1133));
  OAI221_X1 g0933(.A(new_n899), .B1(new_n202), .B2(new_n820), .C1(new_n361), .C2(new_n827), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n825), .A2(new_n260), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n1134), .A2(new_n1103), .A3(new_n1135), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n896), .A2(new_n835), .B1(new_n819), .B2(new_n1109), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT51), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n837), .A2(G143), .B1(G68), .B2(new_n809), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT117), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1136), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n790), .B1(new_n1133), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n251), .A2(new_n798), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n795), .B1(G97), .B2(new_n720), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n788), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1142), .B(new_n1146), .C1(new_n1025), .C2(new_n862), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1055), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1147), .B1(new_n1042), .B2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1125), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(G390));
  NAND2_X1  g0951(.A1(new_n887), .A2(new_n924), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n869), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n776), .B2(new_n872), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n982), .B1(new_n1154), .B2(new_n922), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1155), .A2(new_n979), .A3(new_n980), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n669), .A2(new_n670), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n555), .B(new_n1157), .C1(new_n698), .C2(new_n710), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n769), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(new_n773), .A3(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1160), .A2(new_n872), .A3(new_n714), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n869), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n922), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n983), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT119), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1164), .A2(new_n963), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1165), .B1(new_n1164), .B2(new_n963), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1152), .B(new_n1156), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g0968(.A(KEYINPUT120), .B(new_n1156), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n918), .A2(G330), .A3(new_n872), .A4(new_n1163), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1153), .B1(new_n774), .B2(new_n872), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n982), .B1(new_n1173), .B2(new_n922), .ZN(new_n1174));
  NOR3_X1   g0974(.A1(new_n949), .A2(new_n950), .A3(new_n947), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n937), .B1(new_n690), .B2(new_n691), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT37), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n940), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n688), .B1(new_n972), .B2(new_n973), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n957), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1178), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1175), .B1(new_n947), .B2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(KEYINPUT119), .B1(new_n1174), .B2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1164), .A2(new_n963), .A3(new_n1165), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(KEYINPUT120), .B1(new_n1185), .B2(new_n1156), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1168), .B1(new_n1172), .B2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n918), .A2(G330), .A3(new_n872), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1162), .B1(new_n1188), .B2(new_n922), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1152), .A2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n872), .B1(new_n763), .B2(new_n766), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1171), .B1(new_n1191), .B2(new_n922), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1190), .B1(new_n1192), .B2(new_n1154), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n450), .A2(G330), .A3(new_n918), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1194), .B(new_n696), .C1(new_n987), .C2(new_n777), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1193), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n782), .B1(new_n1187), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1168), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n978), .B1(new_n946), .B2(new_n951), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n1182), .B2(new_n978), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1183), .A2(new_n1184), .B1(new_n1201), .B2(new_n1155), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1170), .B1(new_n1202), .B2(KEYINPUT120), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1156), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT120), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1199), .B1(new_n1203), .B2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n923), .B1(new_n885), .B2(new_n886), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1170), .B1(new_n1208), .B2(new_n1163), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1154), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1209), .A2(new_n1210), .B1(new_n1152), .B2(new_n1189), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1211), .A2(new_n1195), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1207), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1198), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1207), .A2(new_n1055), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n788), .B1(new_n361), .B2(new_n890), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n902), .B1(G107), .B2(new_n851), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1217), .B(new_n508), .C1(new_n217), .C2(new_n810), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n828), .A2(G97), .B1(new_n829), .B2(G116), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1219), .B1(new_n841), .B2(new_n819), .C1(new_n848), .C2(new_n897), .ZN(new_n1220));
  NOR3_X1   g1020(.A1(new_n1218), .A2(new_n1220), .A3(new_n1135), .ZN(new_n1221));
  INV_X1    g1021(.A(G128), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n257), .B1(new_n819), .B2(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n810), .A2(new_n1109), .ZN(new_n1224));
  XOR2_X1   g1024(.A(KEYINPUT121), .B(KEYINPUT53), .Z(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n1224), .A2(new_n1226), .B1(new_n835), .B2(new_n825), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n1223), .B(new_n1227), .C1(new_n1224), .C2(new_n1226), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n813), .A2(G50), .B1(new_n829), .B2(G132), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(KEYINPUT54), .B(G143), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n828), .A2(new_n1231), .B1(new_n851), .B2(G137), .ZN(new_n1232));
  INV_X1    g1032(.A(G125), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1229), .B(new_n1232), .C1(new_n848), .C2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1221), .B1(new_n1228), .B2(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1236), .A2(KEYINPUT122), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(KEYINPUT122), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n790), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1216), .B1(new_n1237), .B2(new_n1239), .C1(new_n981), .C2(new_n792), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1214), .A2(new_n1215), .A3(new_n1240), .ZN(G378));
  OAI21_X1  g1041(.A(new_n1196), .B1(new_n1187), .B2(new_n1211), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT57), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n955), .A2(G330), .A3(new_n964), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n299), .A2(new_n701), .ZN(new_n1246));
  XOR2_X1   g1046(.A(new_n311), .B(new_n1246), .Z(new_n1247));
  XOR2_X1   g1047(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1248));
  AND2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n971), .A2(KEYINPUT106), .A3(new_n974), .ZN(new_n1252));
  AOI21_X1  g1052(.A(KEYINPUT106), .B1(new_n971), .B2(new_n974), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1251), .B1(new_n1254), .B2(new_n984), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n977), .A2(new_n984), .A3(new_n1251), .A4(new_n985), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1245), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1251), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n986), .A2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1260), .A2(new_n1244), .A3(new_n1256), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1242), .A2(new_n1243), .A3(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1243), .B1(new_n1242), .B2(new_n1262), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n721), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1251), .A2(new_n791), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n890), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1076), .B1(G50), .B2(new_n1267), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n857), .A2(G116), .B1(G107), .B2(new_n829), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n205), .B2(new_n820), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n813), .A2(G58), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1271), .B1(new_n363), .B2(new_n827), .ZN(new_n1272));
  AOI211_X1 g1072(.A(G41), .B(new_n1272), .C1(G77), .C2(new_n809), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1273), .A2(new_n1103), .A3(new_n1061), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n1270), .B(new_n1274), .C1(G283), .C2(new_n849), .ZN(new_n1275));
  OR2_X1    g1075(.A1(new_n1275), .A2(KEYINPUT58), .ZN(new_n1276));
  INV_X1    g1076(.A(G132), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n819), .A2(new_n1233), .B1(new_n820), .B2(new_n1277), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n1231), .A2(new_n809), .B1(new_n829), .B2(G128), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n908), .B2(new_n827), .ZN(new_n1280));
  AOI211_X1 g1080(.A(new_n1278), .B(new_n1280), .C1(G150), .C2(new_n824), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  OR2_X1    g1082(.A1(new_n1282), .A2(KEYINPUT59), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(KEYINPUT59), .ZN(new_n1284));
  INV_X1    g1084(.A(G41), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n390), .B(new_n1285), .C1(new_n814), .C2(new_n835), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1286), .B1(G124), .B2(new_n837), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1283), .A2(new_n1284), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1275), .A2(KEYINPUT58), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1285), .B1(new_n1103), .B2(new_n390), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n202), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1276), .A2(new_n1288), .A3(new_n1289), .A4(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1268), .B1(new_n1292), .B2(new_n790), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n1262), .A2(new_n1055), .B1(new_n1266), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1265), .A2(new_n1294), .ZN(G375));
  INV_X1    g1095(.A(new_n1023), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1195), .B(new_n1190), .C1(new_n1192), .C2(new_n1154), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1197), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n922), .A2(new_n791), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1076), .B1(G68), .B2(new_n1267), .ZN(new_n1300));
  OAI22_X1  g1100(.A1(new_n896), .A2(new_n841), .B1(new_n820), .B2(new_n616), .ZN(new_n1301));
  AOI211_X1 g1101(.A(new_n257), .B(new_n1301), .C1(G77), .C2(new_n813), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n849), .A2(G303), .ZN(new_n1303));
  OAI22_X1  g1103(.A1(new_n810), .A2(new_n205), .B1(new_n827), .B2(new_n206), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1304), .B1(G294), .B2(new_n857), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1302), .A2(new_n1112), .A3(new_n1303), .A4(new_n1305), .ZN(new_n1306));
  OAI221_X1 g1106(.A(new_n1271), .B1(new_n1109), .B2(new_n827), .C1(new_n835), .C2(new_n810), .ZN(new_n1307));
  AOI211_X1 g1107(.A(new_n1103), .B(new_n1307), .C1(G50), .C2(new_n824), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1308), .B1(new_n1222), .B2(new_n848), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(new_n1309), .B(KEYINPUT123), .ZN(new_n1310));
  AOI22_X1  g1110(.A1(G132), .A2(new_n857), .B1(new_n851), .B2(new_n1231), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1311), .B1(new_n908), .B2(new_n896), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1306), .B1(new_n1310), .B2(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1300), .B1(new_n1313), .B2(new_n790), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1299), .A2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(new_n1211), .B2(new_n1148), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1298), .A2(new_n1317), .ZN(G381));
  INV_X1    g1118(.A(new_n1294), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1195), .B1(new_n1207), .B2(new_n1212), .ZN(new_n1320));
  AND3_X1   g1120(.A1(new_n1260), .A2(new_n1244), .A3(new_n1256), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1244), .B1(new_n1260), .B2(new_n1256), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(KEYINPUT57), .B1(new_n1320), .B2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1242), .A2(new_n1262), .A3(new_n1243), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1319), .B1(new_n1326), .B2(new_n721), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1056), .A2(new_n1150), .A3(new_n1080), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  AND3_X1   g1129(.A1(new_n1214), .A2(new_n1215), .A3(new_n1240), .ZN(new_n1330));
  INV_X1    g1130(.A(G396), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1121), .A2(new_n1331), .A3(new_n1122), .ZN(new_n1332));
  NOR3_X1   g1132(.A1(new_n1332), .A2(G381), .A3(G384), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1327), .A2(new_n1329), .A3(new_n1330), .A4(new_n1333), .ZN(G407));
  NAND2_X1  g1134(.A1(new_n1327), .A2(new_n1330), .ZN(new_n1335));
  OAI211_X1 g1135(.A(G407), .B(G213), .C1(G343), .C2(new_n1335), .ZN(G409));
  INV_X1    g1136(.A(KEYINPUT125), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n782), .B1(new_n1193), .B2(new_n1196), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1297), .A2(KEYINPUT60), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT60), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1340), .B1(new_n1211), .B2(new_n1195), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1338), .B1(new_n1339), .B2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT124), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1342), .A2(new_n1343), .A3(G384), .A4(new_n1317), .ZN(new_n1344));
  INV_X1    g1144(.A(G384), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n721), .B1(new_n1211), .B2(new_n1195), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1297), .A2(KEYINPUT60), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1211), .A2(new_n1340), .A3(new_n1195), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1346), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1345), .B1(new_n1349), .B2(new_n1316), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1344), .A2(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1316), .B1(new_n1352), .B2(new_n1338), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1343), .B1(new_n1353), .B2(G384), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1337), .B1(new_n1351), .B2(new_n1354), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1342), .A2(G384), .A3(new_n1317), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1356), .A2(KEYINPUT124), .ZN(new_n1357));
  NAND4_X1  g1157(.A1(new_n1357), .A2(KEYINPUT125), .A3(new_n1344), .A4(new_n1350), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1355), .A2(new_n1358), .ZN(new_n1359));
  INV_X1    g1159(.A(new_n1359), .ZN(new_n1360));
  INV_X1    g1160(.A(G213), .ZN(new_n1361));
  NOR2_X1   g1161(.A1(new_n1361), .A2(G343), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1265), .A2(G378), .A3(new_n1294), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1242), .A2(new_n1262), .A3(new_n1296), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1294), .A2(new_n1364), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1330), .A2(new_n1365), .ZN(new_n1366));
  AOI21_X1  g1166(.A(new_n1362), .B1(new_n1363), .B2(new_n1366), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1360), .A2(new_n1367), .A3(KEYINPUT63), .ZN(new_n1368));
  AOI21_X1  g1168(.A(new_n1150), .B1(new_n1056), .B2(new_n1080), .ZN(new_n1369));
  INV_X1    g1169(.A(KEYINPUT127), .ZN(new_n1370));
  INV_X1    g1170(.A(new_n1122), .ZN(new_n1371));
  OAI21_X1  g1171(.A(G396), .B1(new_n1371), .B2(new_n1120), .ZN(new_n1372));
  AOI21_X1  g1172(.A(new_n1370), .B1(new_n1372), .B2(new_n1332), .ZN(new_n1373));
  AND3_X1   g1173(.A1(new_n1372), .A2(new_n1332), .A3(new_n1370), .ZN(new_n1374));
  OAI22_X1  g1174(.A1(new_n1329), .A2(new_n1369), .B1(new_n1373), .B2(new_n1374), .ZN(new_n1375));
  INV_X1    g1175(.A(new_n1369), .ZN(new_n1376));
  NOR2_X1   g1176(.A1(new_n1374), .A2(new_n1373), .ZN(new_n1377));
  NAND3_X1  g1177(.A1(new_n1376), .A2(new_n1377), .A3(new_n1328), .ZN(new_n1378));
  INV_X1    g1178(.A(KEYINPUT61), .ZN(new_n1379));
  NAND3_X1  g1179(.A1(new_n1375), .A2(new_n1378), .A3(new_n1379), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1360), .A2(new_n1367), .ZN(new_n1381));
  INV_X1    g1181(.A(KEYINPUT63), .ZN(new_n1382));
  AOI21_X1  g1182(.A(new_n1380), .B1(new_n1381), .B2(new_n1382), .ZN(new_n1383));
  NAND2_X1  g1183(.A1(new_n1362), .A2(G2897), .ZN(new_n1384));
  AND2_X1   g1184(.A1(new_n1344), .A2(new_n1350), .ZN(new_n1385));
  AOI21_X1  g1185(.A(new_n1384), .B1(new_n1385), .B2(new_n1357), .ZN(new_n1386));
  INV_X1    g1186(.A(new_n1386), .ZN(new_n1387));
  NAND3_X1  g1187(.A1(new_n1355), .A2(new_n1358), .A3(new_n1384), .ZN(new_n1388));
  AOI21_X1  g1188(.A(G378), .B1(new_n1294), .B2(new_n1364), .ZN(new_n1389));
  AOI21_X1  g1189(.A(new_n1389), .B1(new_n1327), .B2(G378), .ZN(new_n1390));
  OAI211_X1 g1190(.A(new_n1387), .B(new_n1388), .C1(new_n1390), .C2(new_n1362), .ZN(new_n1391));
  INV_X1    g1191(.A(KEYINPUT126), .ZN(new_n1392));
  NOR2_X1   g1192(.A1(new_n1391), .A2(new_n1392), .ZN(new_n1393));
  NAND2_X1  g1193(.A1(new_n1363), .A2(new_n1366), .ZN(new_n1394));
  INV_X1    g1194(.A(new_n1362), .ZN(new_n1395));
  AOI21_X1  g1195(.A(new_n1386), .B1(new_n1394), .B2(new_n1395), .ZN(new_n1396));
  AOI21_X1  g1196(.A(KEYINPUT126), .B1(new_n1396), .B2(new_n1388), .ZN(new_n1397));
  OAI211_X1 g1197(.A(new_n1368), .B(new_n1383), .C1(new_n1393), .C2(new_n1397), .ZN(new_n1398));
  AOI21_X1  g1198(.A(new_n782), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1399));
  NOR3_X1   g1199(.A1(new_n1399), .A2(new_n1330), .A3(new_n1319), .ZN(new_n1400));
  OAI21_X1  g1200(.A(new_n1395), .B1(new_n1400), .B2(new_n1389), .ZN(new_n1401));
  OAI21_X1  g1201(.A(KEYINPUT62), .B1(new_n1401), .B2(new_n1359), .ZN(new_n1402));
  INV_X1    g1202(.A(KEYINPUT62), .ZN(new_n1403));
  NAND3_X1  g1203(.A1(new_n1360), .A2(new_n1367), .A3(new_n1403), .ZN(new_n1404));
  NAND4_X1  g1204(.A1(new_n1402), .A2(new_n1379), .A3(new_n1404), .A4(new_n1391), .ZN(new_n1405));
  NAND2_X1  g1205(.A1(new_n1375), .A2(new_n1378), .ZN(new_n1406));
  NAND2_X1  g1206(.A1(new_n1405), .A2(new_n1406), .ZN(new_n1407));
  NAND2_X1  g1207(.A1(new_n1398), .A2(new_n1407), .ZN(G405));
  NAND2_X1  g1208(.A1(G375), .A2(G378), .ZN(new_n1409));
  NAND2_X1  g1209(.A1(new_n1409), .A2(new_n1335), .ZN(new_n1410));
  OAI21_X1  g1210(.A(new_n1410), .B1(new_n1354), .B2(new_n1351), .ZN(new_n1411));
  NAND3_X1  g1211(.A1(new_n1360), .A2(new_n1335), .A3(new_n1409), .ZN(new_n1412));
  NAND2_X1  g1212(.A1(new_n1411), .A2(new_n1412), .ZN(new_n1413));
  XNOR2_X1  g1213(.A(new_n1413), .B(new_n1406), .ZN(G402));
endmodule


