//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n550,
    new_n552, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n613, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1200, new_n1201, new_n1202,
    new_n1203;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT67), .Z(G319));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n458), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(KEYINPUT68), .B1(new_n460), .B2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n462), .A2(new_n458), .A3(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n459), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G137), .ZN(new_n465));
  NAND2_X1  g040(.A1(G101), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n458), .A2(G2104), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n468), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n464), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n461), .A2(new_n463), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(new_n469), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(new_n478), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n478), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n481), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND3_X1  g064(.A1(new_n478), .A2(G102), .A3(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(G114), .A2(G2104), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n492), .B1(new_n464), .B2(G126), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n490), .B1(new_n493), .B2(new_n478), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n482), .A2(G138), .A3(new_n478), .A4(new_n469), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n496), .A2(new_n497), .A3(new_n478), .A4(G138), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n498), .B1(new_n496), .B2(new_n497), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n495), .A2(KEYINPUT4), .B1(new_n471), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n494), .A2(new_n500), .ZN(G164));
  AND2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  OR2_X1    g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  NAND3_X1  g080(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g082(.A(G543), .B1(KEYINPUT70), .B2(KEYINPUT5), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n507), .A2(new_n508), .B1(new_n503), .B2(new_n502), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n505), .A2(G50), .B1(new_n510), .B2(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(new_n506), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n515), .A2(G62), .ZN(new_n516));
  AND2_X1   g091(.A1(G75), .A2(G543), .ZN(new_n517));
  OAI211_X1 g092(.A(KEYINPUT71), .B(G651), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n511), .A2(new_n518), .A3(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  AND2_X1   g099(.A1(new_n510), .A2(G89), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n504), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G51), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n527), .B(new_n528), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n525), .A2(new_n531), .ZN(G168));
  INV_X1    g107(.A(G52), .ZN(new_n533));
  XNOR2_X1  g108(.A(KEYINPUT72), .B(G90), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n529), .A2(new_n533), .B1(new_n509), .B2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n521), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n535), .A2(new_n537), .ZN(G171));
  XNOR2_X1  g113(.A(KEYINPUT73), .B(G43), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n505), .A2(new_n539), .B1(new_n510), .B2(G81), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(KEYINPUT74), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(KEYINPUT74), .ZN(new_n543));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(new_n515), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n542), .A2(new_n543), .B1(G651), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT75), .ZN(G188));
  NAND3_X1  g130(.A1(new_n505), .A2(KEYINPUT9), .A3(G53), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n529), .B2(new_n558), .ZN(new_n559));
  AND2_X1   g134(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n545), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n563), .A2(G651), .B1(G91), .B2(new_n510), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n560), .A2(new_n564), .ZN(G299));
  INV_X1    g140(.A(G171), .ZN(G301));
  AND2_X1   g141(.A1(G168), .A2(KEYINPUT76), .ZN(new_n567));
  NOR2_X1   g142(.A1(G168), .A2(KEYINPUT76), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n567), .A2(new_n568), .ZN(G286));
  OR3_X1    g144(.A1(new_n507), .A2(G74), .A3(new_n508), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n505), .A2(G49), .B1(new_n570), .B2(G651), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n572));
  INV_X1    g147(.A(G87), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n509), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n510), .A2(KEYINPUT77), .A3(G87), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n571), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT78), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n571), .A2(new_n578), .A3(new_n575), .A4(new_n574), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(new_n579), .ZN(G288));
  OAI211_X1 g155(.A(G48), .B(G543), .C1(new_n502), .C2(new_n503), .ZN(new_n581));
  INV_X1    g156(.A(G86), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n509), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g158(.A(G61), .B1(new_n507), .B2(new_n508), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(KEYINPUT79), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT79), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n515), .A2(new_n587), .A3(G61), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n583), .B1(new_n589), .B2(G651), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G305));
  INV_X1    g166(.A(G47), .ZN(new_n592));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  OAI22_X1  g168(.A1(new_n529), .A2(new_n592), .B1(new_n509), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n595), .A2(new_n521), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n545), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(new_n505), .B2(G54), .ZN(new_n603));
  INV_X1    g178(.A(G92), .ZN(new_n604));
  OAI21_X1  g179(.A(KEYINPUT10), .B1(new_n509), .B2(new_n604), .ZN(new_n605));
  OR3_X1    g180(.A1(new_n509), .A2(KEYINPUT10), .A3(new_n604), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n603), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n599), .B1(new_n608), .B2(G868), .ZN(G321));
  XOR2_X1   g184(.A(G321), .B(KEYINPUT80), .Z(G284));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(G299), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(G286), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(new_n611), .ZN(G297));
  OAI21_X1  g189(.A(new_n612), .B1(new_n613), .B2(new_n611), .ZN(G280));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n608), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n547), .A2(G651), .ZN(new_n618));
  INV_X1    g193(.A(new_n543), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n541), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(new_n611), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n607), .A2(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n611), .B2(new_n622), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g199(.A1(new_n478), .A2(G111), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT82), .Z(new_n626));
  OAI211_X1 g201(.A(new_n626), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n484), .A2(G123), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n480), .A2(G135), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(G2096), .Z(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n632));
  NOR3_X1   g207(.A1(new_n458), .A2(new_n460), .A3(G2105), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(KEYINPUT13), .B(G2100), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n631), .A2(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2435), .ZN(new_n639));
  XOR2_X1   g214(.A(G2427), .B(G2438), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(KEYINPUT14), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT16), .Z(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n642), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n642), .B(new_n644), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(new_n647), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n649), .A2(new_n651), .A3(new_n653), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(G14), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT83), .ZN(G401));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n659), .B1(new_n662), .B2(KEYINPUT18), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2096), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2100), .ZN(new_n665));
  AND2_X1   g240(.A1(new_n662), .A2(KEYINPUT17), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n660), .A2(new_n661), .ZN(new_n667));
  AOI21_X1  g242(.A(KEYINPUT18), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n665), .B(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(G227));
  XOR2_X1   g245(.A(G1956), .B(G2474), .Z(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n671), .A2(new_n672), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n677), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n674), .A2(new_n676), .A3(new_n678), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n681), .B(new_n682), .C1(new_n680), .C2(new_n679), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT21), .B(G1986), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1991), .B(G1996), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT84), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT22), .B(G1981), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n688), .B(new_n689), .Z(G229));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G25), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n480), .A2(G131), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n484), .A2(G119), .ZN(new_n694));
  NOR2_X1   g269(.A1(G95), .A2(G2105), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT85), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n696), .B(G2104), .C1(G107), .C2(new_n478), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n693), .A2(new_n694), .A3(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n692), .B1(new_n699), .B2(new_n691), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT35), .B(G1991), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G24), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(new_n597), .B2(new_n703), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G1986), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n700), .A2(new_n701), .ZN(new_n707));
  NOR3_X1   g282(.A1(new_n702), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n703), .A2(G22), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G166), .B2(new_n703), .ZN(new_n711));
  INV_X1    g286(.A(G1971), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  MUX2_X1   g288(.A(G23), .B(new_n576), .S(G16), .Z(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT33), .B(G1976), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n703), .A2(G6), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(new_n590), .B2(new_n703), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT32), .B(G1981), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n718), .B(new_n719), .Z(new_n720));
  AND3_X1   g295(.A1(new_n713), .A2(new_n716), .A3(new_n720), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n721), .A2(KEYINPUT34), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(KEYINPUT34), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n709), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT86), .B(KEYINPUT36), .Z(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT91), .B(KEYINPUT23), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n703), .A2(G20), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G299), .B2(G16), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1956), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n691), .A2(G27), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G164), .B2(new_n691), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G2078), .ZN(new_n735));
  NAND2_X1  g310(.A1(G115), .A2(G2104), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n469), .A2(new_n470), .ZN(new_n737));
  INV_X1    g312(.A(G127), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G2105), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n478), .A2(G103), .A3(G2104), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT25), .Z(new_n742));
  INV_X1    g317(.A(G139), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n740), .B(new_n742), .C1(new_n743), .C2(new_n479), .ZN(new_n744));
  MUX2_X1   g319(.A(G33), .B(new_n744), .S(G29), .Z(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G2072), .ZN(new_n746));
  NOR2_X1   g321(.A1(G16), .A2(G21), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G168), .B2(G16), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G1966), .ZN(new_n750));
  NOR2_X1   g325(.A1(G5), .A2(G16), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G171), .B2(G16), .ZN(new_n752));
  OAI22_X1  g327(.A1(new_n749), .A2(new_n750), .B1(G1961), .B2(new_n752), .ZN(new_n753));
  NOR3_X1   g328(.A1(new_n735), .A2(new_n746), .A3(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n691), .A2(G26), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n480), .A2(G140), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n484), .A2(G128), .ZN(new_n759));
  NOR2_X1   g334(.A1(G104), .A2(G2105), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT88), .Z(new_n761));
  OAI211_X1 g336(.A(new_n761), .B(G2104), .C1(G116), .C2(new_n478), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n758), .A2(new_n759), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n757), .B1(new_n763), .B2(G29), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G2067), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n480), .A2(G141), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n484), .A2(G129), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n478), .A2(G105), .A3(G2104), .ZN(new_n768));
  NAND3_X1  g343(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT26), .Z(new_n770));
  NAND4_X1  g345(.A1(new_n766), .A2(new_n767), .A3(new_n768), .A4(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G29), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G29), .B2(G32), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT27), .B(G1996), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT90), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  AND4_X1   g352(.A1(new_n732), .A2(new_n754), .A3(new_n765), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n691), .A2(G35), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G162), .B2(new_n691), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT29), .B(G2090), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  AND2_X1   g357(.A1(KEYINPUT24), .A2(G34), .ZN(new_n783));
  NOR2_X1   g358(.A1(KEYINPUT24), .A2(G34), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n783), .A2(new_n784), .A3(G29), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n476), .B2(G29), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G2084), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT30), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(G28), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(G28), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n789), .A2(new_n790), .A3(new_n691), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n787), .B(new_n791), .C1(new_n691), .C2(new_n630), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n750), .B2(new_n749), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n774), .A2(new_n776), .B1(G1961), .B2(new_n752), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n778), .A2(new_n782), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n724), .B2(new_n726), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n703), .A2(G4), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n608), .B2(new_n703), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(G1348), .Z(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT31), .B(G11), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n727), .A2(new_n796), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n703), .A2(G19), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n548), .B2(new_n703), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT87), .B(G1341), .Z(new_n804));
  XOR2_X1   g379(.A(new_n803), .B(new_n804), .Z(new_n805));
  NOR2_X1   g380(.A1(new_n801), .A2(new_n805), .ZN(G311));
  INV_X1    g381(.A(G311), .ZN(G150));
  AOI22_X1  g382(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n808));
  OR3_X1    g383(.A1(new_n808), .A2(KEYINPUT92), .A3(new_n521), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n505), .A2(G55), .B1(new_n510), .B2(G93), .ZN(new_n810));
  OAI21_X1  g385(.A(KEYINPUT92), .B1(new_n808), .B2(new_n521), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n812), .A2(KEYINPUT93), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(KEYINPUT93), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(G860), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT94), .B(KEYINPUT37), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n608), .A2(G559), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT38), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT39), .Z(new_n821));
  NAND3_X1  g396(.A1(new_n813), .A2(new_n620), .A3(new_n814), .ZN(new_n822));
  INV_X1    g397(.A(new_n812), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n548), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n821), .B(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n818), .B1(new_n826), .B2(G860), .ZN(G145));
  XNOR2_X1  g402(.A(new_n630), .B(new_n476), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(new_n488), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT97), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n744), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(KEYINPUT96), .B2(new_n744), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(new_n763), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n698), .B(KEYINPUT99), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n484), .A2(G130), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT98), .ZN(new_n837));
  OR2_X1    g412(.A1(G106), .A2(G2105), .ZN(new_n838));
  INV_X1    g413(.A(G118), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n460), .B1(new_n839), .B2(G2105), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n480), .A2(G142), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n835), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(KEYINPUT95), .B1(new_n494), .B2(new_n500), .ZN(new_n844));
  INV_X1    g419(.A(new_n490), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n462), .B1(new_n458), .B2(G2104), .ZN(new_n846));
  NOR3_X1   g421(.A1(new_n460), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n847));
  OAI211_X1 g422(.A(G126), .B(new_n469), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(new_n491), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n845), .B1(new_n849), .B2(G2105), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n499), .A2(new_n471), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT95), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n850), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n844), .A2(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n698), .A2(KEYINPUT99), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n698), .A2(KEYINPUT99), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n857), .A2(new_n841), .A3(new_n837), .A4(new_n858), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n843), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n856), .B1(new_n843), .B2(new_n859), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n834), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n843), .A2(new_n859), .ZN(new_n863));
  INV_X1    g438(.A(new_n856), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n834), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n843), .A2(new_n856), .A3(new_n859), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n771), .B(new_n634), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n862), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n869), .B1(new_n862), .B2(new_n868), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n830), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(KEYINPUT101), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT101), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n874), .B(new_n830), .C1(new_n870), .C2(new_n871), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n862), .A2(new_n868), .ZN(new_n877));
  INV_X1    g452(.A(new_n869), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n862), .A2(new_n868), .A3(new_n869), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(new_n829), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(KEYINPUT100), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n879), .A2(new_n883), .A3(new_n829), .A4(new_n880), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G37), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n876), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT40), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT40), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n876), .A2(new_n885), .A3(new_n889), .A4(new_n886), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(G395));
  NAND2_X1  g466(.A1(new_n825), .A2(new_n622), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n822), .B(new_n824), .C1(G559), .C2(new_n607), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n608), .A2(new_n564), .A3(new_n560), .ZN(new_n896));
  NAND2_X1  g471(.A1(G299), .A2(new_n607), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT41), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n894), .A2(new_n895), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n895), .B1(new_n894), .B2(new_n899), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n898), .B(KEYINPUT102), .Z(new_n904));
  OR2_X1    g479(.A1(new_n904), .A2(new_n894), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT108), .ZN(new_n906));
  XNOR2_X1  g481(.A(G305), .B(new_n576), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(G290), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n576), .B(new_n590), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n597), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n912));
  XNOR2_X1  g487(.A(G303), .B(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(KEYINPUT104), .ZN(new_n914));
  XNOR2_X1  g489(.A(G303), .B(KEYINPUT105), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n911), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n908), .A2(new_n914), .A3(new_n917), .A4(new_n910), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n906), .B1(new_n922), .B2(KEYINPUT42), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n906), .A3(KEYINPUT42), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n903), .B(new_n905), .C1(new_n923), .C2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n902), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n927), .A2(new_n905), .A3(new_n900), .ZN(new_n928));
  INV_X1    g503(.A(new_n923), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(new_n929), .A3(new_n924), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n919), .A2(new_n921), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n920), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n926), .A2(new_n930), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n934), .B1(new_n926), .B2(new_n930), .ZN(new_n936));
  OAI21_X1  g511(.A(G868), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n815), .A2(new_n611), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(G295));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n938), .ZN(G331));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n941));
  OAI21_X1  g516(.A(G171), .B1(new_n567), .B2(new_n568), .ZN(new_n942));
  NAND2_X1  g517(.A1(G301), .A2(G168), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n825), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n944), .A2(new_n822), .A3(new_n824), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n948), .A2(new_n904), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT41), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n898), .B(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n951), .B1(new_n947), .B2(new_n946), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n932), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n948), .A2(new_n899), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n954), .B(new_n931), .C1(new_n898), .C2(new_n948), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(new_n955), .A3(new_n886), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n953), .A2(new_n955), .A3(KEYINPUT109), .A4(new_n886), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n941), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n948), .A2(new_n898), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n932), .B1(new_n961), .B2(new_n952), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n962), .A2(new_n955), .A3(new_n886), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n963), .A2(new_n941), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT44), .B1(new_n960), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n953), .A2(new_n955), .A3(new_n941), .A4(new_n886), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n965), .A2(new_n970), .ZN(G397));
  INV_X1    g546(.A(KEYINPUT119), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n850), .A2(new_n853), .ZN(new_n973));
  INV_X1    g548(.A(G1384), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT45), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n465), .A2(new_n466), .ZN(new_n976));
  OAI211_X1 g551(.A(G40), .B(new_n475), .C1(new_n976), .C2(G2105), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n972), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  OAI211_X1 g553(.A(KEYINPUT45), .B(new_n974), .C1(new_n494), .C2(new_n500), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT120), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n973), .A2(KEYINPUT120), .A3(KEYINPUT45), .A4(new_n974), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n478), .B1(new_n472), .B2(new_n473), .ZN(new_n984));
  INV_X1    g559(.A(G40), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n467), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(G1384), .B1(new_n850), .B2(new_n853), .ZN(new_n987));
  OAI211_X1 g562(.A(KEYINPUT119), .B(new_n986), .C1(new_n987), .C2(KEYINPUT45), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n989), .A2(G2078), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n978), .A2(new_n983), .A3(new_n988), .A4(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT50), .B1(new_n973), .B2(new_n974), .ZN(new_n992));
  OAI211_X1 g567(.A(KEYINPUT50), .B(new_n974), .C1(new_n494), .C2(new_n500), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n986), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G1961), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n991), .A2(G301), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT125), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n494), .A2(new_n500), .A3(KEYINPUT95), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n854), .B1(new_n850), .B2(new_n853), .ZN(new_n1001));
  OAI211_X1 g576(.A(KEYINPUT45), .B(new_n974), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G2078), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n974), .B1(new_n494), .B2(new_n500), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n977), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1002), .A2(new_n1003), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n999), .B1(new_n1007), .B2(new_n989), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n1007), .A2(new_n999), .A3(new_n989), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n998), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(G1384), .B1(new_n844), .B2(new_n855), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n977), .B1(new_n1011), .B2(KEYINPUT45), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n856), .A2(new_n974), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n1005), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1012), .A2(new_n1014), .A3(new_n990), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n997), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1007), .A2(new_n989), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT125), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1007), .A2(new_n999), .A3(new_n989), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1016), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1010), .B(KEYINPUT54), .C1(new_n1020), .C2(G301), .ZN(new_n1021));
  INV_X1    g596(.A(G8), .ZN(new_n1022));
  NOR2_X1   g597(.A1(G168), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT51), .B1(new_n1023), .B2(KEYINPUT124), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n978), .A2(new_n983), .A3(new_n988), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n750), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1004), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n977), .B1(new_n1028), .B2(new_n993), .ZN(new_n1029));
  INV_X1    g604(.A(G2084), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1026), .A2(new_n1031), .ZN(new_n1032));
  OR2_X1    g607(.A1(new_n525), .A2(new_n531), .ZN(new_n1033));
  OAI211_X1 g608(.A(G8), .B(new_n1024), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1032), .A2(G8), .A3(new_n1033), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1023), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1024), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n1025), .A2(new_n750), .B1(new_n1030), .B2(new_n1029), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1036), .B(new_n1037), .C1(new_n1038), .C2(new_n1022), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1034), .A2(new_n1035), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT114), .ZN(new_n1041));
  OAI211_X1 g616(.A(G303), .B(G8), .C1(new_n1041), .C2(KEYINPUT55), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(KEYINPUT55), .ZN(new_n1043));
  XOR2_X1   g618(.A(new_n1043), .B(KEYINPUT115), .Z(new_n1044));
  XNOR2_X1  g619(.A(new_n1042), .B(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G2090), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1029), .A2(KEYINPUT113), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n986), .B1(new_n987), .B2(KEYINPUT45), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1049), .B1(KEYINPUT45), .B2(new_n1011), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1048), .B1(new_n1050), .B2(G1971), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT113), .B1(new_n1029), .B2(new_n1047), .ZN(new_n1052));
  OAI211_X1 g627(.A(G8), .B(new_n1046), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT49), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT117), .ZN(new_n1055));
  INV_X1    g630(.A(G1981), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n590), .A2(new_n1056), .ZN(new_n1057));
  AOI211_X1 g632(.A(G1981), .B(new_n583), .C1(new_n589), .C2(G651), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n1057), .A2(new_n1058), .A3(KEYINPUT116), .ZN(new_n1059));
  NAND3_X1  g634(.A1(G305), .A2(KEYINPUT116), .A3(G1981), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1055), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT116), .B1(new_n590), .B2(new_n1056), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(new_n1056), .B2(new_n590), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1064), .A2(KEYINPUT117), .A3(new_n1054), .A4(new_n1060), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1004), .A2(new_n977), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1066), .A2(new_n1022), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1062), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1976), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1067), .B1(new_n1069), .B2(new_n576), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT52), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT52), .B1(G288), .B2(new_n1069), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1072), .B(new_n1067), .C1(new_n1069), .C2(new_n576), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1068), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n995), .A2(G2090), .ZN(new_n1075));
  AOI21_X1  g650(.A(G1971), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1076));
  OAI21_X1  g651(.A(G8), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(new_n1045), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1053), .A2(new_n1074), .A3(new_n1078), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1021), .A2(new_n1040), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n991), .A2(new_n997), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1081), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT126), .B1(new_n1082), .B2(G301), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT126), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1009), .A2(new_n1008), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1084), .B(G171), .C1(new_n1085), .C2(new_n1081), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1020), .A2(G301), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1083), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(G1956), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n995), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(KEYINPUT121), .A2(KEYINPUT57), .ZN(new_n1096));
  NAND3_X1  g671(.A1(G299), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n560), .A2(new_n1093), .A3(new_n1094), .A4(new_n564), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g675(.A(KEYINPUT56), .B(G2072), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1002), .A2(new_n1006), .A3(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1092), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(G2067), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1066), .A2(KEYINPUT122), .A3(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n987), .A2(new_n1104), .A3(new_n986), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1105), .B(new_n1108), .C1(new_n1029), .C2(G1348), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1103), .A2(new_n608), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1100), .B1(new_n1092), .B2(new_n1102), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1092), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1114), .B1(new_n1115), .B2(new_n1111), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  OAI211_X1 g693(.A(KEYINPUT123), .B(new_n1114), .C1(new_n1115), .C2(new_n1111), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(G1996), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1066), .ZN(new_n1122));
  XOR2_X1   g697(.A(KEYINPUT58), .B(G1341), .Z(new_n1123));
  AOI22_X1  g698(.A1(new_n1050), .A2(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(KEYINPUT59), .B1(new_n1124), .B2(new_n620), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1126), .B1(new_n1127), .B2(G1996), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(new_n1129), .A3(new_n548), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1125), .A2(new_n1130), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n608), .A2(KEYINPUT60), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1109), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1109), .A2(new_n1132), .ZN(new_n1134));
  OAI22_X1  g709(.A1(new_n1133), .A2(new_n1134), .B1(KEYINPUT60), .B2(new_n608), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1112), .A2(KEYINPUT61), .A3(new_n1103), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1131), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1113), .B1(new_n1120), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1080), .A2(new_n1090), .A3(new_n1138), .ZN(new_n1139));
  XOR2_X1   g714(.A(new_n1058), .B(KEYINPUT118), .Z(new_n1140));
  NAND2_X1  g715(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1140), .B1(new_n1141), .B2(G288), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n1067), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1074), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1143), .B1(new_n1053), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT63), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1053), .A2(new_n1074), .A3(new_n1078), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1038), .A2(new_n1022), .A3(G286), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1146), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(G8), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1146), .B1(new_n1151), .B2(new_n1045), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1152), .A2(new_n1053), .A3(new_n1074), .A4(new_n1148), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1145), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1040), .A2(KEYINPUT62), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT62), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1034), .A2(new_n1157), .A3(new_n1035), .A4(new_n1039), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1155), .A2(new_n1156), .A3(new_n1079), .A4(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1139), .A2(new_n1154), .A3(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1013), .A2(new_n1005), .A3(new_n986), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT110), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1013), .A2(KEYINPUT110), .A3(new_n1005), .A4(new_n986), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n772), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1161), .A2(G1996), .ZN(new_n1166));
  OAI22_X1  g741(.A1(new_n1165), .A2(new_n1166), .B1(G1996), .B2(new_n772), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n763), .B(G2067), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT111), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1168), .A2(KEYINPUT111), .A3(new_n1169), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1167), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(KEYINPUT112), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT112), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1167), .A2(new_n1172), .A3(new_n1176), .A4(new_n1173), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n698), .A2(new_n701), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n698), .A2(new_n701), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1168), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1175), .A2(new_n1177), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1161), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n597), .B(G1986), .Z(new_n1183));
  AOI21_X1  g758(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1160), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1168), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1175), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1187));
  OR2_X1    g762(.A1(new_n763), .A2(G2067), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1186), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  XOR2_X1   g764(.A(new_n1166), .B(KEYINPUT46), .Z(new_n1190));
  OAI211_X1 g765(.A(new_n1190), .B(new_n1170), .C1(new_n772), .C2(new_n1186), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT47), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1191), .B(new_n1192), .ZN(new_n1193));
  NOR3_X1   g768(.A1(new_n1161), .A2(G1986), .A3(G290), .ZN(new_n1194));
  XOR2_X1   g769(.A(new_n1194), .B(KEYINPUT48), .Z(new_n1195));
  AND4_X1   g770(.A1(new_n1175), .A2(new_n1177), .A3(new_n1180), .A4(new_n1195), .ZN(new_n1196));
  NOR3_X1   g771(.A1(new_n1189), .A2(new_n1193), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1185), .A2(new_n1197), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g773(.A1(new_n657), .A2(new_n456), .A3(new_n669), .ZN(new_n1200));
  XNOR2_X1  g774(.A(new_n1200), .B(KEYINPUT127), .ZN(new_n1201));
  AOI21_X1  g775(.A(new_n1201), .B1(new_n966), .B2(new_n967), .ZN(new_n1202));
  INV_X1    g776(.A(G229), .ZN(new_n1203));
  AND3_X1   g777(.A1(new_n887), .A2(new_n1202), .A3(new_n1203), .ZN(G308));
  NAND3_X1  g778(.A1(new_n887), .A2(new_n1202), .A3(new_n1203), .ZN(G225));
endmodule


