//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 0 0 0 1 1 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT28), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT64), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT64), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n190), .B1(new_n195), .B2(new_n189), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT0), .A2(G128), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT0), .A2(G128), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT65), .B1(new_n196), .B2(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT66), .B1(new_n191), .B2(G143), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT64), .B(G146), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G143), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT66), .ZN(new_n206));
  AND4_X1   g020(.A1(new_n206), .A2(new_n192), .A3(new_n194), .A4(G143), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n198), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT11), .ZN(new_n209));
  INV_X1    g023(.A(G134), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(G137), .ZN(new_n211));
  INV_X1    g025(.A(G137), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(KEYINPUT11), .A3(G134), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n210), .A2(G137), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n211), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G131), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(KEYINPUT67), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n217), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n219), .A2(new_n211), .A3(new_n213), .A4(new_n214), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n222));
  AOI21_X1  g036(.A(G143), .B1(new_n192), .B2(new_n194), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n222), .B(new_n200), .C1(new_n223), .C2(new_n190), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n202), .A2(new_n208), .A3(new_n221), .A4(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n215), .A2(new_n216), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n212), .A2(G134), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(new_n214), .A3(G131), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G128), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n192), .A2(new_n194), .A3(G143), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT1), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT68), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT1), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n230), .B1(new_n231), .B2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(new_n196), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G128), .ZN(new_n240));
  INV_X1    g054(.A(new_n203), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n231), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n192), .A2(new_n194), .A3(new_n206), .A4(G143), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n240), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n229), .B1(new_n238), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n225), .A2(new_n245), .ZN(new_n246));
  OR2_X1    g060(.A1(KEYINPUT71), .A2(G116), .ZN(new_n247));
  NAND2_X1  g061(.A1(KEYINPUT71), .A2(G116), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(G119), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n250));
  INV_X1    g064(.A(G119), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(KEYINPUT70), .A2(G119), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(G116), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT2), .B(G113), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT72), .ZN(new_n258));
  INV_X1    g072(.A(new_n256), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(new_n249), .A3(new_n254), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n255), .A2(KEYINPUT72), .A3(new_n256), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n246), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n263), .A2(new_n225), .A3(new_n245), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n188), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n188), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(G237), .A2(G953), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G210), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n271), .B(KEYINPUT27), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT26), .B(G101), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n272), .B(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NOR3_X1   g089(.A1(new_n267), .A2(new_n269), .A3(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT74), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n187), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n266), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n263), .B1(new_n225), .B2(new_n245), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT28), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(new_n268), .A3(new_n274), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT30), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n246), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT69), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n246), .A2(KEYINPUT69), .A3(new_n283), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n225), .A2(new_n245), .A3(KEYINPUT30), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n289), .A2(new_n264), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n279), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n282), .B1(new_n291), .B2(new_n274), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n278), .B1(new_n292), .B2(new_n277), .ZN(new_n293));
  INV_X1    g107(.A(G902), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT75), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n295), .B1(new_n276), .B2(KEYINPUT29), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n281), .A2(KEYINPUT29), .A3(new_n268), .A4(new_n274), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n297), .A2(KEYINPUT75), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n294), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G472), .B1(new_n293), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(G472), .A2(G902), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n301), .B(KEYINPUT73), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT69), .B1(new_n246), .B2(new_n283), .ZN(new_n303));
  AOI211_X1 g117(.A(new_n285), .B(KEYINPUT30), .C1(new_n225), .C2(new_n245), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n290), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT31), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n279), .A2(new_n275), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n275), .B1(new_n267), .B2(new_n269), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n306), .B1(new_n305), .B2(new_n307), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n302), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT32), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT32), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n314), .B(new_n302), .C1(new_n310), .C2(new_n311), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n300), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G217), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n318), .B1(G234), .B2(new_n294), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT16), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(G125), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT76), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(G125), .ZN(new_n324));
  INV_X1    g138(.A(G125), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G140), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT16), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n328), .A2(new_n320), .A3(new_n321), .A4(G125), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n323), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n191), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n323), .A2(new_n327), .A3(G146), .A4(new_n329), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT23), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n252), .A2(G128), .A3(new_n253), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n230), .A2(G119), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT70), .B(G119), .ZN(new_n338));
  AOI21_X1  g152(.A(KEYINPUT23), .B1(new_n338), .B2(new_n230), .ZN(new_n339));
  OAI21_X1  g153(.A(G110), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n335), .A2(new_n336), .ZN(new_n341));
  XOR2_X1   g155(.A(KEYINPUT24), .B(G110), .Z(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n333), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(G125), .B(G140), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n204), .A2(new_n345), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n332), .A2(new_n346), .ZN(new_n347));
  NOR3_X1   g161(.A1(new_n337), .A2(new_n339), .A3(G110), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n341), .A2(new_n342), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(KEYINPUT22), .B(G137), .ZN(new_n351));
  INV_X1    g165(.A(G953), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(G221), .A3(G234), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n351), .B(new_n353), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n344), .A2(new_n350), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n354), .B1(new_n344), .B2(new_n350), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT25), .B1(new_n357), .B2(new_n294), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n344), .A2(new_n350), .ZN(new_n359));
  INV_X1    g173(.A(new_n354), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n344), .A2(new_n350), .A3(new_n354), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n361), .A2(KEYINPUT25), .A3(new_n294), .A4(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n319), .B1(new_n358), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT77), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n361), .A2(new_n294), .A3(new_n362), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT25), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n363), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT77), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n371), .A3(new_n319), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n319), .A2(G902), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(KEYINPUT78), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n357), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n366), .A2(new_n372), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(G214), .B1(G237), .B2(G902), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n249), .A2(new_n254), .A3(KEYINPUT5), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n381), .B(G113), .C1(KEYINPUT5), .C2(new_n254), .ZN(new_n382));
  INV_X1    g196(.A(G104), .ZN(new_n383));
  OAI21_X1  g197(.A(KEYINPUT3), .B1(new_n383), .B2(G107), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT3), .ZN(new_n385));
  INV_X1    g199(.A(G107), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(G104), .ZN(new_n387));
  INV_X1    g201(.A(G101), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n383), .A2(G107), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n384), .A2(new_n387), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n383), .A2(G107), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n386), .A2(G104), .ZN(new_n392));
  OAI21_X1  g206(.A(G101), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n382), .A2(new_n260), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n384), .A2(new_n387), .A3(new_n389), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G101), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(KEYINPUT4), .A3(new_n390), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n397), .A2(new_n400), .A3(G101), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n396), .B1(new_n263), .B2(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(G110), .B(G122), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n404), .B(new_n396), .C1(new_n263), .C2(new_n402), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(KEYINPUT6), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n352), .A2(G224), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(KEYINPUT79), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n224), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n197), .B1(new_n242), .B2(new_n243), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n325), .B1(new_n414), .B2(new_n202), .ZN(new_n415));
  INV_X1    g229(.A(new_n190), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n416), .B1(new_n204), .B2(G143), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n239), .B1(G143), .B2(new_n204), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n417), .B1(new_n418), .B2(new_n230), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n236), .A2(new_n230), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n420), .B1(new_n205), .B2(new_n207), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n419), .A2(new_n325), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n411), .B1(new_n415), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n202), .A2(new_n208), .A3(new_n224), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(G125), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n426), .A2(new_n422), .A3(new_n410), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT6), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n403), .A2(new_n429), .A3(new_n405), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n408), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT80), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT80), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n408), .A2(new_n428), .A3(new_n433), .A4(new_n430), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  XOR2_X1   g249(.A(KEYINPUT81), .B(KEYINPUT8), .Z(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(new_n404), .ZN(new_n437));
  INV_X1    g251(.A(new_n396), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n395), .B1(new_n382), .B2(new_n260), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT7), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n440), .B(new_n407), .C1(new_n427), .C2(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT83), .B(KEYINPUT7), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n411), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT82), .ZN(new_n445));
  AOI22_X1  g259(.A1(new_n445), .A2(new_n422), .B1(new_n425), .B2(G125), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n423), .A2(KEYINPUT82), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n444), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n294), .B1(new_n442), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n435), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(G210), .B1(G237), .B2(G902), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n435), .A2(new_n452), .A3(new_n450), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n380), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(G110), .B(G140), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n352), .A2(G227), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n457), .B(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n221), .ZN(new_n460));
  OAI21_X1  g274(.A(G128), .B1(new_n190), .B2(new_n232), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n242), .A2(new_n243), .A3(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n395), .B1(new_n462), .B2(new_n244), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT10), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n419), .A2(new_n421), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n394), .A2(new_n464), .ZN(new_n466));
  AOI22_X1  g280(.A1(new_n463), .A2(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OR2_X1    g281(.A1(new_n425), .A2(new_n402), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n460), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n466), .B1(new_n238), .B2(new_n244), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n242), .A2(new_n243), .A3(new_n461), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n394), .B1(new_n421), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n470), .B1(new_n472), .B2(KEYINPUT10), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n425), .A2(new_n402), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n473), .A2(new_n474), .A3(new_n221), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n459), .B1(new_n469), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n467), .A2(new_n468), .A3(new_n460), .ZN(new_n477));
  INV_X1    g291(.A(new_n459), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n419), .A2(new_n421), .A3(new_n394), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n463), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT12), .B1(new_n480), .B2(new_n221), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT12), .ZN(new_n482));
  AOI211_X1 g296(.A(new_n482), .B(new_n460), .C1(new_n463), .C2(new_n479), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n477), .B(new_n478), .C1(new_n481), .C2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(G902), .B1(new_n476), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(G469), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n477), .B1(new_n481), .B2(new_n483), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n459), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n221), .B1(new_n473), .B2(new_n474), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n477), .A2(new_n490), .A3(new_n478), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n489), .A2(G469), .A3(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n486), .A2(new_n294), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n487), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT9), .B(G234), .ZN(new_n496));
  OAI21_X1  g310(.A(G221), .B1(new_n496), .B2(G902), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n230), .A2(G143), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT13), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n210), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n189), .A2(G128), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n230), .A2(G143), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT13), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n503), .A3(new_n210), .ZN(new_n505));
  AOI22_X1  g319(.A1(new_n501), .A2(new_n504), .B1(new_n505), .B2(KEYINPUT88), .ZN(new_n506));
  OR2_X1    g320(.A1(new_n505), .A2(KEYINPUT88), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n247), .A2(G122), .A3(new_n248), .ZN(new_n508));
  INV_X1    g322(.A(G122), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(G116), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(new_n386), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n386), .B1(new_n508), .B2(new_n510), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n506), .B(new_n507), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n502), .A2(new_n503), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(G134), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n505), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT14), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n508), .A2(new_n518), .A3(new_n510), .ZN(new_n519));
  OAI21_X1  g333(.A(G107), .B1(new_n508), .B2(new_n518), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n511), .B(new_n517), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  NOR3_X1   g335(.A1(new_n496), .A2(new_n318), .A3(G953), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n514), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT89), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT89), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n514), .A2(new_n521), .A3(new_n525), .A4(new_n522), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n514), .A2(new_n521), .ZN(new_n527));
  INV_X1    g341(.A(new_n522), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n524), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n294), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT91), .ZN(new_n532));
  INV_X1    g346(.A(G478), .ZN(new_n533));
  OAI22_X1  g347(.A1(new_n531), .A2(new_n532), .B1(KEYINPUT15), .B2(new_n533), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n530), .A2(KEYINPUT90), .A3(new_n294), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT90), .B1(new_n530), .B2(new_n294), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n533), .A2(KEYINPUT15), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n538), .B1(new_n531), .B2(KEYINPUT91), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n534), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT87), .ZN(new_n541));
  XOR2_X1   g355(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(G113), .B(G122), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n544), .B(new_n383), .ZN(new_n545));
  INV_X1    g359(.A(G237), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(new_n352), .A3(G214), .ZN(new_n547));
  NOR2_X1   g361(.A1(KEYINPUT85), .A2(G143), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n270), .B(G214), .C1(KEYINPUT85), .C2(G143), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AND2_X1   g365(.A1(KEYINPUT18), .A2(G131), .ZN(new_n552));
  OR2_X1    g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n552), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n346), .B1(new_n191), .B2(new_n345), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n551), .A2(KEYINPUT17), .A3(G131), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n331), .A2(new_n557), .A3(new_n332), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT86), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n331), .A2(new_n557), .A3(KEYINPUT86), .A4(new_n332), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n551), .A2(G131), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT17), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n549), .A2(new_n550), .A3(new_n216), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n545), .B(new_n556), .C1(new_n560), .C2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n545), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n345), .B(KEYINPUT19), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n204), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n562), .A2(new_n564), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n571), .A3(new_n332), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n556), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n568), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n567), .A2(new_n575), .ZN(new_n576));
  OR2_X1    g390(.A1(G475), .A2(G902), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n541), .B(new_n543), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n577), .B1(new_n567), .B2(new_n575), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT87), .B1(new_n579), .B2(new_n542), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT20), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n578), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n556), .B1(new_n560), .B2(new_n566), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n584), .A2(new_n568), .ZN(new_n585));
  INV_X1    g399(.A(new_n567), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n294), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(G475), .ZN(new_n588));
  INV_X1    g402(.A(G234), .ZN(new_n589));
  OAI211_X1 g403(.A(G952), .B(new_n352), .C1(new_n589), .C2(new_n546), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(KEYINPUT92), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  OAI211_X1 g406(.A(G902), .B(G953), .C1(new_n589), .C2(new_n546), .ZN(new_n593));
  XOR2_X1   g407(.A(new_n593), .B(KEYINPUT93), .Z(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT21), .B(G898), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n592), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n540), .A2(new_n583), .A3(new_n588), .A4(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n498), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n317), .A2(new_n378), .A3(new_n456), .A4(new_n600), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT94), .B(G101), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G3));
  AOI21_X1  g417(.A(new_n452), .B1(new_n435), .B2(new_n450), .ZN(new_n604));
  AOI211_X1 g418(.A(new_n453), .B(new_n449), .C1(new_n432), .C2(new_n434), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n379), .B(new_n598), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n535), .ZN(new_n607));
  INV_X1    g421(.A(new_n536), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(new_n533), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n610), .B1(new_n527), .B2(new_n528), .ZN(new_n611));
  AOI22_X1  g425(.A1(new_n530), .A2(new_n610), .B1(new_n523), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(G478), .A3(new_n294), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n583), .A2(new_n588), .B1(new_n609), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n606), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n312), .ZN(new_n617));
  OAI211_X1 g431(.A(KEYINPUT95), .B(new_n294), .C1(new_n310), .C2(new_n311), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n618), .A2(G472), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT95), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n289), .A2(new_n264), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n286), .B2(new_n287), .ZN(new_n622));
  INV_X1    g436(.A(new_n307), .ZN(new_n623));
  OAI21_X1  g437(.A(KEYINPUT31), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n624), .A2(new_n309), .A3(new_n308), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n620), .B1(new_n626), .B2(G902), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n617), .B1(new_n619), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n498), .A2(new_n377), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n616), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(new_n630), .B(KEYINPUT96), .Z(new_n631));
  XOR2_X1   g445(.A(KEYINPUT34), .B(G104), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  NAND2_X1  g447(.A1(new_n579), .A2(new_n542), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n578), .A2(new_n580), .A3(new_n634), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n635), .A2(new_n588), .ZN(new_n636));
  INV_X1    g450(.A(new_n540), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n606), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n639), .A2(new_n628), .A3(new_n629), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT35), .B(G107), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  OAI21_X1  g456(.A(new_n379), .B1(new_n604), .B2(new_n605), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n360), .A2(KEYINPUT36), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT97), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(new_n359), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n375), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n366), .A2(new_n372), .A3(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(new_n497), .A3(new_n495), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n643), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n599), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n650), .A2(new_n628), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT37), .B(G110), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G12));
  AND2_X1   g468(.A1(new_n650), .A2(new_n317), .ZN(new_n655));
  INV_X1    g469(.A(G900), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n592), .B1(new_n595), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n638), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT98), .B(G128), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G30));
  NOR2_X1   g475(.A1(new_n604), .A2(new_n605), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT38), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n663), .A2(new_n380), .A3(new_n648), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n657), .B(KEYINPUT39), .Z(new_n665));
  NAND3_X1  g479(.A1(new_n495), .A2(new_n497), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT100), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n667), .A2(KEYINPUT40), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(KEYINPUT40), .ZN(new_n669));
  INV_X1    g483(.A(G472), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n275), .B1(new_n279), .B2(new_n280), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT99), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n671), .A2(KEYINPUT99), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n672), .B(new_n673), .C1(new_n622), .C2(new_n623), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n670), .B1(new_n674), .B2(new_n294), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(new_n313), .B2(new_n315), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n583), .A2(new_n588), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n637), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n664), .A2(new_n668), .A3(new_n669), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G143), .ZN(G45));
  INV_X1    g495(.A(new_n657), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n614), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n655), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G146), .ZN(G48));
  AOI21_X1  g500(.A(new_n377), .B1(new_n300), .B2(new_n316), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n485), .A2(new_n486), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(new_n497), .A3(new_n487), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n616), .A2(new_n687), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT41), .B(G113), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G15));
  NAND3_X1  g507(.A1(new_n639), .A2(new_n687), .A3(new_n690), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G116), .ZN(G18));
  AOI21_X1  g509(.A(new_n371), .B1(new_n370), .B2(new_n319), .ZN(new_n696));
  INV_X1    g510(.A(new_n319), .ZN(new_n697));
  AOI211_X1 g511(.A(KEYINPUT77), .B(new_n697), .C1(new_n369), .C2(new_n363), .ZN(new_n698));
  INV_X1    g512(.A(new_n647), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n696), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n700), .A2(new_n599), .ZN(new_n701));
  INV_X1    g515(.A(new_n315), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n314), .B1(new_n625), .B2(new_n302), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n278), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n274), .B1(new_n305), .B2(new_n266), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n277), .B1(new_n706), .B2(new_n276), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n276), .A2(new_n295), .A3(KEYINPUT29), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n297), .A2(KEYINPUT75), .ZN(new_n710));
  AOI21_X1  g524(.A(G902), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n670), .B1(new_n708), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n701), .B1(new_n704), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n456), .A2(new_n690), .ZN(new_n714));
  OAI21_X1  g528(.A(KEYINPUT101), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n643), .A2(new_n689), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT101), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n716), .A2(new_n317), .A3(new_n717), .A4(new_n701), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G119), .ZN(G21));
  AOI21_X1  g534(.A(new_n670), .B1(new_n625), .B2(new_n294), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n617), .A2(new_n721), .A3(new_n377), .ZN(new_n722));
  INV_X1    g536(.A(new_n678), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n689), .A2(new_n597), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n722), .A2(new_n456), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  INV_X1    g540(.A(KEYINPUT102), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n727), .B1(new_n614), .B2(new_n682), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n614), .A2(new_n727), .A3(new_n682), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n700), .A2(new_n721), .A3(new_n617), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n716), .A2(new_n729), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G125), .ZN(G27));
  NAND2_X1  g547(.A1(new_n609), .A2(new_n613), .ZN(new_n734));
  AND4_X1   g548(.A1(new_n727), .A2(new_n677), .A3(new_n734), .A4(new_n682), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n728), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n454), .A2(new_n379), .A3(new_n455), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n493), .B1(new_n485), .B2(new_n486), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT103), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n492), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n489), .A2(KEYINPUT103), .A3(G469), .A4(new_n491), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n738), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n497), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n737), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n736), .A2(new_n687), .A3(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT42), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n736), .A2(new_n687), .A3(new_n744), .A4(KEYINPUT42), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G131), .ZN(G33));
  NAND3_X1  g564(.A1(new_n687), .A2(new_n744), .A3(new_n658), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G134), .ZN(G36));
  AND2_X1   g566(.A1(new_n489), .A2(new_n491), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n753), .A2(KEYINPUT45), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(KEYINPUT45), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(G469), .A3(new_n755), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n756), .A2(new_n494), .ZN(new_n757));
  OR2_X1    g571(.A1(new_n757), .A2(KEYINPUT46), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n756), .A2(KEYINPUT46), .A3(new_n494), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(new_n487), .A3(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n497), .A3(new_n665), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n734), .A2(new_n583), .A3(new_n588), .ZN(new_n762));
  XOR2_X1   g576(.A(new_n762), .B(KEYINPUT43), .Z(new_n763));
  INV_X1    g577(.A(new_n628), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n764), .A3(new_n648), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n761), .A2(new_n737), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n768), .B1(new_n766), .B2(new_n765), .ZN(new_n769));
  XOR2_X1   g583(.A(KEYINPUT104), .B(G137), .Z(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(G39));
  NAND2_X1  g585(.A1(new_n760), .A2(new_n497), .ZN(new_n772));
  XNOR2_X1  g586(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT47), .ZN(new_n775));
  AOI22_X1  g589(.A1(new_n760), .A2(new_n497), .B1(KEYINPUT105), .B2(new_n775), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n317), .A2(new_n737), .A3(new_n378), .A4(new_n683), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT106), .ZN(new_n778));
  OR3_X1    g592(.A1(new_n774), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G140), .ZN(G42));
  NAND2_X1  g594(.A1(new_n688), .A2(new_n487), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT107), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT49), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n676), .A2(new_n378), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n497), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n762), .A2(new_n380), .A3(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n783), .A2(new_n663), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  XOR2_X1   g602(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n789));
  NOR2_X1   g603(.A1(new_n737), .A2(new_n689), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n785), .A2(new_n592), .A3(new_n790), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n791), .A2(new_n677), .A3(new_n734), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n763), .A2(new_n592), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n793), .A2(KEYINPUT114), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(KEYINPUT114), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n796), .A2(new_n790), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n792), .B1(new_n797), .B2(new_n731), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n796), .A2(new_n722), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n782), .A2(KEYINPUT115), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n782), .A2(KEYINPUT115), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n800), .A2(new_n786), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n802), .B1(new_n774), .B2(new_n776), .ZN(new_n803));
  INV_X1    g617(.A(new_n737), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n799), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n798), .A2(new_n805), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n663), .A2(new_n380), .A3(new_n690), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n799), .A2(KEYINPUT50), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n796), .A2(new_n722), .A3(new_n807), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT50), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n806), .B1(KEYINPUT116), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n808), .A2(new_n814), .A3(new_n811), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n789), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  OAI211_X1 g630(.A(G952), .B(new_n352), .C1(new_n791), .C2(new_n615), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n817), .B1(new_n799), .B2(new_n716), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT48), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n797), .A2(new_n819), .A3(new_n687), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n819), .B1(new_n797), .B2(new_n687), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n818), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT117), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n818), .B(KEYINPUT117), .C1(new_n820), .C2(new_n821), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n812), .A2(KEYINPUT51), .A3(new_n805), .A4(new_n798), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n676), .A2(new_n643), .A3(new_n678), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT109), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n738), .A2(new_n740), .A3(new_n741), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n497), .B1(new_n657), .B2(KEYINPUT108), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n832), .B1(KEYINPUT108), .B2(new_n657), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n366), .A2(new_n372), .A3(new_n647), .A4(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n830), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n700), .A2(new_n742), .A3(KEYINPUT109), .A4(new_n833), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n829), .A2(new_n837), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n650), .B(new_n317), .C1(new_n658), .C2(new_n684), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(new_n839), .A3(new_n732), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT52), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n838), .A2(new_n839), .A3(new_n842), .A4(new_n732), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n736), .A2(new_n731), .A3(new_n744), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n636), .A2(new_n540), .A3(new_n682), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n846), .A2(new_n649), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n317), .A3(new_n804), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n845), .A2(new_n751), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n749), .A2(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n652), .A2(new_n601), .A3(new_n725), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n628), .A2(new_n629), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n615), .B1(new_n677), .B2(new_n540), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(new_n456), .A3(new_n598), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n687), .B(new_n690), .C1(new_n616), .C2(new_n639), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n851), .A2(new_n719), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n844), .A2(new_n850), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT53), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT111), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n841), .A2(new_n860), .A3(new_n843), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n652), .A2(new_n601), .A3(new_n725), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n863), .B1(new_n718), .B2(new_n715), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n691), .A2(new_n694), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n852), .A2(new_n854), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n864), .A2(new_n749), .A3(new_n867), .A4(new_n849), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n860), .B1(new_n841), .B2(new_n843), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n862), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n828), .B(new_n859), .C1(new_n870), .C2(KEYINPUT53), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT112), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT110), .B1(new_n858), .B2(KEYINPUT53), .ZN(new_n874));
  INV_X1    g688(.A(new_n869), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n850), .A2(new_n857), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n875), .A2(new_n876), .A3(KEYINPUT53), .A4(new_n861), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT110), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT53), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n878), .B(new_n879), .C1(new_n868), .C2(new_n844), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n874), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT54), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n875), .A2(new_n876), .A3(new_n861), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n879), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n884), .A2(KEYINPUT112), .A3(new_n828), .A4(new_n859), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n873), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n816), .A2(new_n827), .A3(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(G952), .A2(G953), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n788), .B1(new_n887), .B2(new_n888), .ZN(G75));
  INV_X1    g703(.A(KEYINPUT56), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n408), .A2(new_n430), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(new_n428), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT55), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n884), .A2(new_n859), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n894), .A2(G210), .A3(G902), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT118), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n890), .B(new_n893), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n897), .B1(new_n896), .B2(new_n895), .ZN(new_n898));
  OR2_X1    g712(.A1(new_n352), .A2(G952), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(KEYINPUT119), .Z(new_n900));
  AND2_X1   g714(.A1(new_n895), .A2(new_n890), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n900), .B1(new_n901), .B2(new_n893), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n898), .A2(new_n902), .ZN(G51));
  INV_X1    g717(.A(new_n900), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n894), .A2(KEYINPUT54), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n871), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n493), .B(KEYINPUT57), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n476), .A2(new_n484), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT120), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n894), .A2(G902), .ZN(new_n912));
  OR2_X1    g726(.A1(new_n912), .A2(new_n756), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n904), .B1(new_n911), .B2(new_n913), .ZN(G54));
  NAND4_X1  g728(.A1(new_n894), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n915));
  INV_X1    g729(.A(new_n576), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n915), .A2(new_n916), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n904), .B1(new_n917), .B2(new_n918), .ZN(G60));
  NAND2_X1  g733(.A1(G478), .A2(G902), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT59), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n612), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n904), .B1(new_n906), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n612), .B1(new_n886), .B2(new_n921), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n923), .B1(new_n924), .B2(KEYINPUT121), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT121), .ZN(new_n926));
  AOI211_X1 g740(.A(new_n926), .B(new_n612), .C1(new_n886), .C2(new_n921), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n925), .A2(new_n927), .ZN(G63));
  INV_X1    g742(.A(KEYINPUT61), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n929), .A2(KEYINPUT124), .ZN(new_n930));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT122), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT60), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n894), .A2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n357), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n904), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n646), .B(KEYINPUT123), .Z(new_n937));
  NAND3_X1  g751(.A1(new_n894), .A2(new_n933), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n930), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n929), .A2(KEYINPUT124), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(G66));
  XOR2_X1   g755(.A(new_n857), .B(KEYINPUT125), .Z(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n352), .ZN(new_n943));
  INV_X1    g757(.A(G224), .ZN(new_n944));
  OAI21_X1  g758(.A(G953), .B1(new_n596), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n891), .B1(G898), .B2(new_n352), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(G69));
  NAND2_X1  g762(.A1(new_n288), .A2(new_n289), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(new_n569), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n950), .B1(G900), .B2(G953), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n687), .A2(new_n456), .A3(new_n723), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n751), .B1(new_n761), .B2(new_n952), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n839), .A2(new_n732), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n779), .A2(new_n769), .A3(new_n749), .A4(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n951), .B1(new_n957), .B2(G953), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n352), .B1(G227), .B2(G900), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n958), .B1(KEYINPUT126), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n680), .A2(new_n954), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT62), .Z(new_n963));
  NAND3_X1  g777(.A1(new_n687), .A2(new_n804), .A3(new_n853), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n964), .A2(new_n667), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n963), .A2(new_n769), .A3(new_n779), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n352), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n961), .B1(new_n967), .B2(new_n950), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n960), .A2(KEYINPUT126), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n968), .B(new_n969), .ZN(G72));
  NAND2_X1  g784(.A1(G472), .A2(G902), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT63), .Z(new_n972));
  OAI21_X1  g786(.A(new_n972), .B1(new_n957), .B2(new_n942), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n973), .A2(KEYINPUT127), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n622), .A2(new_n279), .A3(new_n274), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n973), .A2(KEYINPUT127), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n291), .A2(new_n275), .ZN(new_n978));
  INV_X1    g792(.A(new_n972), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n978), .A2(new_n975), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n881), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n972), .B1(new_n966), .B2(new_n942), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n904), .B1(new_n982), .B2(new_n978), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n977), .A2(new_n981), .A3(new_n983), .ZN(G57));
endmodule


