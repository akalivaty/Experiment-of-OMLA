//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 0 1 1 0 0 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n437, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n582, new_n583, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1194, new_n1195, new_n1196, new_n1197;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT66), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT67), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT68), .Z(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT70), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT70), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G101), .ZN(new_n468));
  NOR3_X1   g043(.A1(new_n467), .A2(new_n468), .A3(G2105), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n473), .A2(G137), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n470), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT71), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n470), .A2(KEYINPUT71), .A3(new_n472), .A4(new_n474), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n469), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G125), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n471), .A2(G2104), .ZN(new_n482));
  OAI21_X1  g057(.A(KEYINPUT69), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n472), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n480), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(G113), .A2(G2104), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g064(.A(G2105), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n479), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT72), .ZN(G160));
  NAND2_X1  g067(.A1(new_n470), .A2(new_n472), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(new_n473), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G124), .ZN(new_n495));
  XOR2_X1   g070(.A(new_n495), .B(KEYINPUT73), .Z(new_n496));
  NOR2_X1   g071(.A1(new_n493), .A2(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G136), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n473), .A2(G112), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n496), .A2(new_n501), .ZN(G162));
  AND3_X1   g077(.A1(new_n472), .A2(new_n484), .A3(new_n485), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n485), .B1(new_n472), .B2(new_n484), .ZN(new_n504));
  OAI211_X1 g079(.A(G138), .B(new_n473), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT4), .A2(G138), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n470), .A2(new_n473), .A3(new_n472), .A4(new_n508), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n470), .A2(G126), .A3(G2105), .A4(new_n472), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT75), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT74), .A2(G114), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT74), .A2(G114), .ZN(new_n513));
  OAI21_X1  g088(.A(G2105), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(G102), .A2(G2105), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n514), .A2(G2104), .A3(new_n515), .ZN(new_n516));
  AND3_X1   g091(.A1(new_n510), .A2(new_n511), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n511), .B1(new_n510), .B2(new_n516), .ZN(new_n518));
  OAI211_X1 g093(.A(new_n507), .B(new_n509), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(G164));
  AOI21_X1  g095(.A(KEYINPUT78), .B1(KEYINPUT77), .B2(KEYINPUT5), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT78), .A2(KEYINPUT5), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n521), .A2(G543), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT6), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(G651), .ZN(new_n529));
  INV_X1    g104(.A(G651), .ZN(new_n530));
  OAI21_X1  g105(.A(KEYINPUT76), .B1(new_n530), .B2(KEYINPUT6), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT76), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n532), .A2(new_n528), .A3(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n529), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n527), .A2(G88), .A3(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(G543), .ZN(new_n536));
  AOI211_X1 g111(.A(new_n536), .B(new_n529), .C1(new_n531), .C2(new_n533), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G50), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n525), .A2(G62), .A3(new_n526), .ZN(new_n539));
  NAND2_X1  g114(.A1(G75), .A2(G543), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g116(.A(new_n535), .B(new_n538), .C1(new_n541), .C2(new_n530), .ZN(G303));
  INV_X1    g117(.A(G303), .ZN(G166));
  NAND2_X1  g118(.A1(new_n534), .A2(G543), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT79), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n545), .A2(G51), .ZN(new_n546));
  NAND3_X1  g121(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT7), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n534), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n525), .A2(new_n526), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n546), .A2(new_n551), .ZN(G168));
  NAND2_X1  g127(.A1(G77), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G64), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n550), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G651), .ZN(new_n556));
  INV_X1    g131(.A(G90), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n527), .A2(new_n534), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n559), .B1(G52), .B2(new_n545), .ZN(G171));
  INV_X1    g135(.A(new_n558), .ZN(new_n561));
  NAND2_X1  g136(.A1(G68), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G56), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n550), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n561), .A2(G81), .B1(G651), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n545), .A2(G43), .ZN(new_n566));
  AND2_X1   g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n550), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n561), .A2(G91), .B1(G651), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(KEYINPUT80), .A2(G53), .ZN(new_n577));
  OR3_X1    g152(.A1(new_n544), .A2(KEYINPUT9), .A3(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(KEYINPUT9), .B1(new_n544), .B2(new_n577), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n576), .A2(new_n580), .ZN(G299));
  XNOR2_X1  g156(.A(new_n537), .B(KEYINPUT79), .ZN(new_n582));
  INV_X1    g157(.A(G52), .ZN(new_n583));
  OAI221_X1 g158(.A(new_n556), .B1(new_n557), .B2(new_n558), .C1(new_n582), .C2(new_n583), .ZN(G301));
  INV_X1    g159(.A(G168), .ZN(G286));
  NAND2_X1  g160(.A1(new_n561), .A2(G87), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n527), .B2(G74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n537), .A2(G49), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  INV_X1    g164(.A(new_n524), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n526), .B(G61), .C1(new_n590), .C2(new_n521), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n593), .A2(G651), .B1(new_n537), .B2(G48), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n534), .A2(new_n525), .A3(G86), .A4(new_n526), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(KEYINPUT81), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT81), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n527), .A2(new_n597), .A3(G86), .A4(new_n534), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n594), .A2(new_n596), .A3(new_n598), .ZN(G305));
  NAND2_X1  g174(.A1(G72), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G60), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n550), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n561), .A2(G85), .B1(G651), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n545), .A2(G47), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  AND3_X1   g181(.A1(new_n527), .A2(G92), .A3(new_n534), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT10), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n545), .A2(G54), .ZN(new_n609));
  XNOR2_X1  g184(.A(KEYINPUT82), .B(G66), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n527), .A2(new_n610), .B1(G79), .B2(G543), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n611), .A2(new_n530), .ZN(new_n612));
  AND3_X1   g187(.A1(new_n608), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(new_n613), .B2(G868), .ZN(G284));
  OAI21_X1  g189(.A(new_n606), .B1(new_n613), .B2(G868), .ZN(G321));
  XOR2_X1   g190(.A(G299), .B(KEYINPUT83), .Z(new_n616));
  MUX2_X1   g191(.A(new_n616), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g192(.A(new_n616), .B(G286), .S(G868), .Z(G280));
  XOR2_X1   g193(.A(KEYINPUT84), .B(G559), .Z(new_n619));
  OAI21_X1  g194(.A(new_n613), .B1(G860), .B2(new_n619), .ZN(G148));
  NAND2_X1  g195(.A1(new_n613), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n567), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g199(.A1(new_n503), .A2(new_n504), .ZN(new_n625));
  OR3_X1    g200(.A1(new_n625), .A2(G2105), .A3(new_n467), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT12), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n628), .A2(G2100), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(G2100), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n497), .A2(G135), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT85), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n494), .A2(G123), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n473), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND3_X1  g212(.A1(new_n629), .A2(new_n630), .A3(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G1341), .B(G1348), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2451), .B(G2454), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT86), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n648), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(G14), .A3(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(G401));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT87), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT17), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2084), .B(G2090), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n661), .B1(new_n658), .B2(new_n660), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n659), .B2(new_n660), .ZN(new_n664));
  INV_X1    g239(.A(new_n660), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n665), .A2(new_n661), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n658), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT18), .ZN(new_n668));
  NOR3_X1   g243(.A1(new_n662), .A2(new_n664), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2096), .B(G2100), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G227));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT89), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n677), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(new_n675), .B2(new_n678), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n680), .B(KEYINPUT90), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n675), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT91), .B(KEYINPUT20), .Z(new_n686));
  OR2_X1    g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n686), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n683), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n693), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G229));
  MUX2_X1   g272(.A(G6), .B(G305), .S(G16), .Z(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT32), .B(G1981), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n698), .B(new_n699), .Z(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G23), .ZN(new_n702));
  INV_X1    g277(.A(G288), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n701), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT33), .B(G1976), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n701), .A2(G22), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G166), .B2(new_n701), .ZN(new_n708));
  INV_X1    g283(.A(G1971), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n700), .A2(new_n706), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(KEYINPUT34), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT93), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n711), .A2(KEYINPUT34), .ZN(new_n714));
  NOR2_X1   g289(.A1(G25), .A2(G29), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n497), .A2(G131), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n494), .A2(G119), .ZN(new_n717));
  OR2_X1    g292(.A1(G95), .A2(G2105), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n718), .B(G2104), .C1(G107), .C2(new_n473), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n716), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n715), .B1(new_n721), .B2(G29), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT35), .B(G1991), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT92), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n722), .B(new_n724), .ZN(new_n725));
  MUX2_X1   g300(.A(G24), .B(G290), .S(G16), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G1986), .ZN(new_n727));
  NOR4_X1   g302(.A1(new_n714), .A2(KEYINPUT94), .A3(new_n725), .A4(new_n727), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n713), .A2(new_n728), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n729), .A2(KEYINPUT36), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n713), .A2(new_n728), .A3(KEYINPUT36), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n613), .A2(new_n701), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G4), .B2(new_n701), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT95), .B(G1348), .Z(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n701), .A2(G20), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT23), .Z(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G299), .B2(G16), .ZN(new_n738));
  INV_X1    g313(.A(G1956), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n735), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G29), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G33), .ZN(new_n743));
  NAND2_X1  g318(.A1(G115), .A2(G2104), .ZN(new_n744));
  INV_X1    g319(.A(G127), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n625), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n473), .B1(new_n746), .B2(KEYINPUT99), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(KEYINPUT99), .B2(new_n746), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT98), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n750), .A2(KEYINPUT25), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(KEYINPUT25), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n751), .A2(new_n752), .B1(G139), .B2(new_n497), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n748), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(KEYINPUT100), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT100), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n748), .A2(new_n756), .A3(new_n753), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n743), .B1(new_n759), .B2(new_n742), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n760), .A2(G2072), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(G2072), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n701), .A2(G19), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n567), .B2(new_n701), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G1341), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n733), .B2(new_n734), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n741), .A2(new_n761), .A3(new_n762), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n742), .A2(G27), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G164), .B2(new_n742), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G2078), .ZN(new_n770));
  NOR2_X1   g345(.A1(G29), .A2(G35), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G162), .B2(G29), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT101), .B(KEYINPUT29), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n770), .B1(new_n774), .B2(G2090), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT30), .B(G28), .ZN(new_n776));
  OR2_X1    g351(.A1(KEYINPUT31), .A2(G11), .ZN(new_n777));
  NAND2_X1  g352(.A1(KEYINPUT31), .A2(G11), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n776), .A2(new_n742), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n636), .B2(new_n742), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n497), .A2(G141), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n494), .A2(G129), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n467), .A2(G2105), .ZN(new_n783));
  NAND3_X1  g358(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT26), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n783), .A2(G105), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n781), .A2(new_n782), .A3(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n790), .A2(new_n742), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n742), .B2(G32), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT27), .B(G1996), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n780), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(G1966), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n701), .A2(G21), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G168), .B2(new_n701), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n794), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n797), .A2(G1966), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n701), .A2(G5), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G171), .B2(new_n701), .ZN(new_n803));
  INV_X1    g378(.A(G1961), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT96), .B(KEYINPUT28), .Z(new_n806));
  NAND2_X1  g381(.A1(new_n742), .A2(G26), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n497), .A2(G140), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n494), .A2(G128), .ZN(new_n811));
  OR2_X1    g386(.A1(G104), .A2(G2105), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n812), .B(G2104), .C1(G116), .C2(new_n473), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n809), .B1(new_n814), .B2(G29), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT97), .B(G2067), .ZN(new_n817));
  OAI22_X1  g392(.A1(new_n792), .A2(new_n793), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(new_n817), .B2(new_n816), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n775), .A2(new_n801), .A3(new_n805), .A4(new_n819), .ZN(new_n820));
  AND2_X1   g395(.A1(KEYINPUT24), .A2(G34), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n742), .B1(KEYINPUT24), .B2(G34), .ZN(new_n822));
  OAI22_X1  g397(.A1(G160), .A2(new_n742), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n823), .A2(G2084), .ZN(new_n824));
  OAI22_X1  g399(.A1(new_n774), .A2(G2090), .B1(G2084), .B2(new_n823), .ZN(new_n825));
  NOR4_X1   g400(.A1(new_n767), .A2(new_n820), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n730), .A2(new_n731), .A3(new_n826), .ZN(G150));
  INV_X1    g402(.A(G150), .ZN(G311));
  NAND2_X1  g403(.A1(new_n613), .A2(G559), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(G80), .A2(G543), .ZN(new_n832));
  INV_X1    g407(.A(G67), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n550), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(G651), .ZN(new_n835));
  INV_X1    g410(.A(G93), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n836), .B2(new_n558), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(G55), .B2(new_n545), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(new_n567), .ZN(new_n839));
  INV_X1    g414(.A(G55), .ZN(new_n840));
  OAI221_X1 g415(.A(new_n835), .B1(new_n836), .B2(new_n558), .C1(new_n582), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n565), .A2(new_n566), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n831), .B(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT39), .ZN(new_n846));
  AOI21_X1  g421(.A(G860), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n846), .B2(new_n845), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n841), .A2(G860), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT37), .Z(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT103), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n848), .A2(KEYINPUT103), .A3(new_n850), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(G145));
  NAND2_X1  g430(.A1(new_n497), .A2(G142), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n494), .A2(G130), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n473), .A2(G118), .ZN(new_n858));
  OAI21_X1  g433(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n856), .B(new_n857), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n627), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n627), .A2(new_n860), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n720), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n627), .A2(new_n860), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n627), .A2(new_n860), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n864), .A2(new_n721), .A3(new_n865), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n510), .A2(new_n516), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n507), .A2(new_n868), .A3(new_n509), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n789), .B(new_n814), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n758), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n870), .B1(new_n755), .B2(new_n757), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n869), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n759), .A2(new_n870), .ZN(new_n875));
  INV_X1    g450(.A(new_n873), .ZN(new_n876));
  INV_X1    g451(.A(new_n869), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AOI211_X1 g453(.A(KEYINPUT104), .B(new_n867), .C1(new_n874), .C2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n874), .ZN(new_n881));
  INV_X1    g456(.A(new_n867), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI22_X1  g458(.A1(new_n879), .A2(new_n883), .B1(new_n881), .B2(new_n882), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n636), .B(G160), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(G162), .Z(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(G37), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n882), .B1(new_n881), .B2(KEYINPUT105), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n889), .B1(KEYINPUT105), .B2(new_n881), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n890), .B(new_n886), .C1(new_n883), .C2(new_n879), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n888), .A2(KEYINPUT40), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT40), .B1(new_n888), .B2(new_n891), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(G395));
  XOR2_X1   g469(.A(new_n621), .B(new_n844), .Z(new_n895));
  INV_X1    g470(.A(G299), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n613), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n608), .A2(new_n609), .A3(new_n612), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(G299), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT41), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n897), .A2(KEYINPUT41), .A3(new_n899), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n895), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n897), .A2(new_n899), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n903), .B1(new_n905), .B2(new_n895), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(KEYINPUT42), .ZN(new_n907));
  XNOR2_X1  g482(.A(G290), .B(G305), .ZN(new_n908));
  XNOR2_X1  g483(.A(G288), .B(G303), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n908), .B(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT42), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n903), .B(new_n912), .C1(new_n905), .C2(new_n895), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n907), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n911), .B1(new_n907), .B2(new_n913), .ZN(new_n915));
  OAI21_X1  g490(.A(G868), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(G868), .B2(new_n838), .ZN(G295));
  OAI21_X1  g492(.A(new_n916), .B1(G868), .B2(new_n838), .ZN(G331));
  NAND2_X1  g493(.A1(G168), .A2(G171), .ZN(new_n919));
  OAI21_X1  g494(.A(G301), .B1(new_n546), .B2(new_n551), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n921), .A2(new_n844), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n922), .A2(new_n904), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n924), .B1(new_n921), .B2(new_n844), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n921), .A2(new_n844), .A3(new_n924), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n923), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n904), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n921), .A2(new_n844), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n930), .B(new_n901), .C1(new_n932), .C2(new_n922), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n928), .A2(new_n933), .A3(new_n910), .ZN(new_n934));
  INV_X1    g509(.A(G37), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n910), .B1(new_n928), .B2(new_n933), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n939));
  INV_X1    g514(.A(new_n922), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n926), .A2(new_n940), .A3(new_n927), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n902), .A2(new_n900), .ZN(new_n942));
  AOI22_X1  g517(.A1(new_n941), .A2(new_n942), .B1(new_n931), .B2(new_n923), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n934), .B(new_n935), .C1(new_n943), .C2(new_n910), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT44), .B1(new_n939), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(new_n938), .B2(new_n945), .ZN(new_n949));
  OAI211_X1 g524(.A(KEYINPUT107), .B(KEYINPUT43), .C1(new_n936), .C2(new_n937), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(new_n944), .B2(KEYINPUT43), .ZN(new_n952));
  INV_X1    g527(.A(new_n936), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n941), .A2(new_n942), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n923), .A2(new_n931), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n911), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n953), .A2(new_n957), .A3(KEYINPUT108), .A4(new_n945), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n949), .A2(new_n950), .B1(new_n952), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n947), .B1(new_n959), .B2(KEYINPUT44), .ZN(G397));
  NAND3_X1  g535(.A1(new_n479), .A2(new_n490), .A3(G40), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n479), .A2(new_n490), .A3(KEYINPUT109), .A4(G40), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n869), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n965), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT111), .ZN(new_n971));
  INV_X1    g546(.A(G2067), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n814), .B(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G1996), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n973), .B1(new_n974), .B2(new_n790), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n971), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n970), .A2(new_n974), .A3(new_n790), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n720), .B(new_n723), .Z(new_n979));
  AOI21_X1  g554(.A(new_n978), .B1(new_n971), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(G290), .A2(G1986), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(G290), .A2(G1986), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n982), .A2(KEYINPUT110), .A3(new_n983), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n984), .B(new_n970), .C1(KEYINPUT110), .C2(new_n983), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n980), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT63), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n593), .A2(G651), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n537), .A2(G48), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n988), .A2(new_n989), .A3(new_n595), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(G1981), .ZN(new_n991));
  INV_X1    g566(.A(G1981), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n594), .A2(new_n992), .A3(new_n596), .A4(new_n598), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT113), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT49), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n991), .A2(new_n993), .A3(KEYINPUT113), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT114), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n996), .A2(new_n1001), .A3(new_n997), .A4(new_n998), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n994), .A2(new_n997), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n506), .A2(new_n505), .B1(new_n497), .B2(new_n508), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1384), .B1(new_n1005), .B2(new_n868), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n963), .A2(new_n1006), .A3(new_n964), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(G8), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT112), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1007), .A2(KEYINPUT112), .A3(G8), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1004), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n703), .A2(G1976), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n1007), .A2(KEYINPUT112), .A3(G8), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT112), .B1(new_n1007), .B2(G8), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  AOI22_X1  g591(.A1(new_n1003), .A2(new_n1012), .B1(new_n1016), .B2(KEYINPUT52), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(new_n703), .B2(G1976), .ZN(new_n1019));
  OR2_X1    g594(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(G168), .A2(G8), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n969), .A2(KEYINPUT115), .A3(new_n963), .A4(new_n964), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n519), .A2(KEYINPUT45), .A3(new_n966), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G40), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n488), .B1(new_n625), .B2(new_n480), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1025), .B1(new_n1026), .B2(G2105), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT109), .B1(new_n1027), .B2(new_n479), .ZN(new_n1028));
  INV_X1    g603(.A(new_n964), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT115), .B1(new_n1030), .B2(new_n969), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n795), .B1(new_n1024), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT50), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n869), .A2(new_n1033), .A3(new_n966), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n963), .A2(new_n1034), .A3(new_n964), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1033), .B1(new_n519), .B2(new_n966), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G2084), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1021), .B1(new_n1032), .B2(new_n1039), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1017), .A2(new_n1020), .A3(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G2090), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n519), .A2(new_n966), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT50), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1030), .A2(new_n1047), .A3(new_n1049), .A4(new_n1034), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n869), .A2(KEYINPUT45), .A3(new_n966), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n963), .A2(new_n1051), .A3(new_n964), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT45), .B1(new_n519), .B2(new_n966), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n709), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1050), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G8), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1046), .B1(new_n1056), .B2(KEYINPUT116), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(KEYINPUT116), .B2(new_n1056), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n987), .B1(new_n1041), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G8), .ZN(new_n1060));
  AOI211_X1 g635(.A(new_n1060), .B(new_n1045), .C1(new_n1050), .C2(new_n1054), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n519), .A2(new_n1033), .A3(new_n966), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n967), .A2(KEYINPUT50), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1030), .A2(new_n1047), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n1054), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1046), .B1(new_n1065), .B2(G8), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1066), .A2(KEYINPUT63), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1061), .B1(new_n1067), .B2(new_n1040), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1070));
  INV_X1    g645(.A(new_n993), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1003), .A2(new_n1012), .ZN(new_n1072));
  NOR2_X1   g647(.A1(G288), .A2(G1976), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1071), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI22_X1  g649(.A1(new_n1068), .A2(new_n1069), .B1(new_n1070), .B2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1059), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1032), .A2(new_n1039), .A3(G168), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT123), .B1(new_n1077), .B2(G8), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT122), .ZN(new_n1079));
  OAI21_X1  g654(.A(KEYINPUT51), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT115), .ZN(new_n1081));
  INV_X1    g656(.A(new_n969), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1081), .B1(new_n1082), .B2(new_n965), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1083), .A2(new_n1023), .A3(new_n1022), .ZN(new_n1084));
  AOI22_X1  g659(.A1(new_n1084), .A2(new_n795), .B1(new_n1038), .B2(new_n1037), .ZN(new_n1085));
  NOR2_X1   g660(.A1(G286), .A2(KEYINPUT123), .ZN(new_n1086));
  OAI22_X1  g661(.A1(new_n1085), .A2(new_n1086), .B1(new_n1079), .B2(KEYINPUT51), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1087), .A2(G8), .A3(new_n1077), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1080), .A2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1066), .A2(new_n1061), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1090), .A2(new_n1017), .A3(new_n1020), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1030), .A2(KEYINPUT119), .A3(new_n1049), .A4(new_n1034), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT119), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1093), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1092), .A2(new_n1094), .A3(new_n804), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT124), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1092), .A2(new_n1094), .A3(KEYINPUT124), .A4(new_n804), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n1100));
  OR3_X1    g675(.A1(new_n1052), .A2(G2078), .A3(new_n1053), .ZN(new_n1101));
  NOR4_X1   g676(.A1(new_n1082), .A2(new_n1100), .A3(G2078), .A4(new_n961), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1100), .A2(new_n1101), .B1(new_n1102), .B2(new_n1051), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(G171), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1101), .A2(new_n1100), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1100), .A2(G2078), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1083), .A2(new_n1023), .A3(new_n1022), .A4(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1106), .A2(new_n1108), .A3(new_n1095), .A4(G301), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1109), .A2(KEYINPUT54), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1091), .B1(new_n1105), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT54), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1099), .A2(new_n1103), .A3(G301), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1106), .A2(new_n1108), .A3(new_n1095), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1114), .A2(G171), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1112), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1089), .A2(new_n1111), .A3(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1063), .A2(new_n1062), .A3(new_n963), .A4(new_n964), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n739), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1048), .A2(new_n968), .ZN(new_n1120));
  XNOR2_X1  g695(.A(KEYINPUT56), .B(G2072), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1030), .A2(new_n1120), .A3(new_n1051), .A4(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT57), .B1(G299), .B2(KEYINPUT117), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT117), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT57), .ZN(new_n1126));
  AOI211_X1 g701(.A(new_n1125), .B(new_n1126), .C1(new_n576), .C2(new_n580), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1123), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1092), .A2(new_n1094), .A3(new_n734), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n963), .A2(new_n1006), .A3(new_n972), .A4(new_n964), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT118), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1132), .B(new_n1133), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1128), .A2(new_n1119), .A3(new_n1122), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n613), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1130), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1136), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1128), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1139), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1131), .A2(new_n1134), .A3(KEYINPUT60), .A4(new_n898), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1130), .A2(KEYINPUT61), .A3(new_n1136), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1131), .A2(new_n1134), .A3(KEYINPUT60), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n613), .ZN(new_n1147));
  AOI21_X1  g722(.A(KEYINPUT60), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1145), .A2(new_n1149), .ZN(new_n1150));
  OR2_X1    g725(.A1(KEYINPUT58), .A2(G1341), .ZN(new_n1151));
  NAND2_X1  g726(.A1(KEYINPUT58), .A2(G1341), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1007), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(KEYINPUT120), .B(G1996), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1052), .A2(new_n1053), .A3(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n567), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(KEYINPUT59), .B1(new_n1156), .B2(KEYINPUT121), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(KEYINPUT121), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1157), .B(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1138), .B1(new_n1150), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1076), .B1(new_n1117), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT62), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1080), .A2(new_n1162), .A3(new_n1088), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1162), .B1(new_n1080), .B2(new_n1088), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1115), .A2(new_n1020), .A3(new_n1017), .A4(new_n1090), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n986), .B1(new_n1161), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(new_n971), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n976), .A2(new_n721), .A3(new_n723), .A4(new_n977), .ZN(new_n1169));
  OR2_X1    g744(.A1(new_n814), .A2(G2067), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1168), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n1171), .A2(KEYINPUT125), .ZN(new_n1172));
  INV_X1    g747(.A(new_n973), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n971), .B1(new_n789), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n970), .A2(new_n974), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1175), .B(KEYINPUT46), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  XOR2_X1   g752(.A(new_n1177), .B(KEYINPUT47), .Z(new_n1178));
  NAND2_X1  g753(.A1(new_n970), .A2(new_n981), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1179), .B(KEYINPUT48), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n980), .A2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1171), .A2(KEYINPUT125), .ZN(new_n1182));
  NOR4_X1   g757(.A1(new_n1172), .A2(new_n1178), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1167), .A2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g759(.A1(new_n888), .A2(new_n891), .ZN(new_n1186));
  NOR2_X1   g760(.A1(G227), .A2(new_n461), .ZN(new_n1187));
  AND2_X1   g761(.A1(new_n655), .A2(new_n1187), .ZN(new_n1188));
  OR2_X1    g762(.A1(new_n1188), .A2(KEYINPUT126), .ZN(new_n1189));
  NAND2_X1  g763(.A1(new_n1188), .A2(KEYINPUT126), .ZN(new_n1190));
  AND3_X1   g764(.A1(new_n696), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g765(.A1(new_n1186), .A2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g766(.A1(new_n1192), .A2(new_n959), .ZN(G308));
  NAND3_X1  g767(.A1(new_n696), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1194));
  AOI21_X1  g768(.A(new_n1194), .B1(new_n888), .B2(new_n891), .ZN(new_n1195));
  AND2_X1   g769(.A1(new_n949), .A2(new_n950), .ZN(new_n1196));
  AND2_X1   g770(.A1(new_n952), .A2(new_n958), .ZN(new_n1197));
  OAI21_X1  g771(.A(new_n1195), .B1(new_n1196), .B2(new_n1197), .ZN(G225));
endmodule


