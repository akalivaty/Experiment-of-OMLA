//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1295, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(new_n203), .A2(G50), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  NOR3_X1   g0008(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT64), .Z(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(G250), .B1(G257), .B2(G264), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n215), .A2(KEYINPUT0), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(KEYINPUT0), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT1), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  AND2_X1   g0023(.A1(new_n211), .A2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n216), .B(new_n217), .C1(new_n218), .C2(new_n224), .ZN(new_n225));
  AOI211_X1 g0025(.A(new_n209), .B(new_n225), .C1(new_n218), .C2(new_n224), .ZN(G361));
  XOR2_X1   g0026(.A(G238), .B(G244), .Z(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G232), .ZN(new_n228));
  XOR2_X1   g0028(.A(KEYINPUT2), .B(G226), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G264), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XOR2_X1   g0034(.A(G87), .B(G116), .Z(new_n235));
  XOR2_X1   g0035(.A(G97), .B(G107), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  INV_X1    g0037(.A(G50), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n238), .A2(G68), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n202), .A2(G50), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n237), .B(new_n243), .Z(G351));
  INV_X1    g0044(.A(G169), .ZN(new_n245));
  AOI21_X1  g0045(.A(new_n208), .B1(G33), .B2(G41), .ZN(new_n246));
  INV_X1    g0046(.A(G1), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G45), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT5), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n249), .A2(G41), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n248), .B1(new_n250), .B2(KEYINPUT76), .ZN(new_n251));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  OAI21_X1  g0052(.A(KEYINPUT76), .B1(new_n252), .B2(KEYINPUT5), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(KEYINPUT5), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n246), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  AND2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  OAI211_X1 g0058(.A(G257), .B(G1698), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  OAI211_X1 g0060(.A(G250), .B(new_n260), .C1(new_n257), .C2(new_n258), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G294), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n259), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  AOI22_X1  g0063(.A1(G264), .A2(new_n256), .B1(new_n263), .B2(new_n246), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  OAI211_X1 g0065(.A(G1), .B(G13), .C1(new_n265), .C2(new_n252), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n251), .A2(new_n255), .A3(G274), .A4(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n245), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n263), .A2(new_n246), .ZN(new_n269));
  INV_X1    g0069(.A(new_n255), .ZN(new_n270));
  INV_X1    g0070(.A(G45), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(G1), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT76), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n272), .B1(new_n254), .B2(new_n273), .ZN(new_n274));
  OAI211_X1 g0074(.A(G264), .B(new_n266), .C1(new_n270), .C2(new_n274), .ZN(new_n275));
  AND4_X1   g0075(.A1(G179), .A2(new_n269), .A3(new_n275), .A4(new_n267), .ZN(new_n276));
  OAI21_X1  g0076(.A(KEYINPUT85), .B1(new_n268), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n247), .A2(G13), .A3(G20), .ZN(new_n278));
  OR3_X1    g0078(.A1(new_n278), .A2(KEYINPUT25), .A3(G107), .ZN(new_n279));
  OAI21_X1  g0079(.A(KEYINPUT25), .B1(new_n278), .B2(G107), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n208), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n247), .A2(G33), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(new_n278), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G107), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n279), .B(new_n280), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT84), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n278), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(new_n282), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(G107), .A3(new_n284), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n292), .A2(KEYINPUT84), .A3(new_n279), .A4(new_n280), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT23), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n295), .B1(new_n207), .B2(G107), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n286), .A2(KEYINPUT23), .A3(G20), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n207), .B(G87), .C1(new_n257), .C2(new_n258), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT22), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT3), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n265), .ZN(new_n304));
  NAND2_X1  g0104(.A1(KEYINPUT3), .A2(G33), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT22), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n306), .A2(new_n307), .A3(new_n207), .A4(G87), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n300), .B1(new_n302), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT24), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n282), .B1(new_n309), .B2(KEYINPUT24), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n294), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n269), .A2(new_n275), .A3(new_n267), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G169), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n264), .A2(G179), .A3(new_n267), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT85), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n277), .A2(new_n313), .A3(new_n318), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n309), .A2(KEYINPUT24), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n320), .A2(new_n282), .A3(new_n310), .ZN(new_n321));
  INV_X1    g0121(.A(new_n314), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G190), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n314), .A2(G200), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n321), .A2(new_n323), .A3(new_n294), .A4(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n319), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT86), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT86), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n319), .A2(new_n328), .A3(new_n325), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT70), .ZN(new_n331));
  AOI21_X1  g0131(.A(G1698), .B1(new_n304), .B2(new_n305), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G222), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n333), .B(KEYINPUT65), .ZN(new_n334));
  INV_X1    g0134(.A(new_n306), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n335), .A2(new_n260), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n336), .A2(G223), .B1(new_n335), .B2(G77), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n266), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n247), .B1(G41), .B2(G45), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G274), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n246), .A2(new_n340), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n342), .B1(new_n343), .B2(G226), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  OR3_X1    g0145(.A1(new_n338), .A2(KEYINPUT66), .A3(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT66), .B1(new_n338), .B2(new_n345), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n331), .B1(new_n348), .B2(G190), .ZN(new_n349));
  INV_X1    g0149(.A(G190), .ZN(new_n350));
  AOI211_X1 g0150(.A(KEYINPUT70), .B(new_n350), .C1(new_n346), .C2(new_n347), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT10), .ZN(new_n353));
  OAI21_X1  g0153(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n354), .B(KEYINPUT68), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT67), .ZN(new_n356));
  NOR2_X1   g0156(.A1(G20), .A2(G33), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G150), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT8), .B(G58), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n207), .A2(G33), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n355), .B1(new_n356), .B2(new_n361), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n361), .A2(new_n356), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n282), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OR2_X1    g0164(.A1(new_n364), .A2(KEYINPUT69), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(KEYINPUT69), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n278), .A2(G50), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n282), .B1(new_n247), .B2(G20), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n367), .B1(new_n368), .B2(G50), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n365), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT9), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n365), .A2(KEYINPUT9), .A3(new_n366), .A4(new_n369), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n348), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G200), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n352), .A2(new_n353), .A3(new_n374), .A4(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n376), .A2(new_n372), .A3(new_n373), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n349), .A2(new_n351), .ZN(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT10), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n332), .A2(G226), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G33), .A2(G97), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n306), .A2(G232), .A3(G1698), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n246), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n342), .B1(new_n343), .B2(G238), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT13), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT13), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n386), .A2(new_n390), .A3(new_n387), .ZN(new_n391));
  AND3_X1   g0191(.A1(new_n389), .A2(G179), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n389), .A2(KEYINPUT71), .A3(new_n391), .ZN(new_n393));
  OR3_X1    g0193(.A1(new_n388), .A2(KEYINPUT71), .A3(KEYINPUT13), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n395), .A2(KEYINPUT14), .A3(G169), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n393), .A2(new_n394), .A3(G169), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT14), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n392), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n357), .A2(KEYINPUT72), .A3(G50), .ZN(new_n401));
  INV_X1    g0201(.A(G77), .ZN(new_n402));
  OAI221_X1 g0202(.A(new_n401), .B1(new_n207), .B2(G68), .C1(new_n402), .C2(new_n360), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT72), .B1(new_n357), .B2(G50), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n282), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT11), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OR3_X1    g0207(.A1(new_n278), .A2(KEYINPUT12), .A3(G68), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT12), .B1(new_n278), .B2(G68), .ZN(new_n409));
  AOI22_X1  g0209(.A1(G68), .A2(new_n368), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(new_n405), .B2(new_n406), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n400), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n395), .A2(G200), .ZN(new_n414));
  INV_X1    g0214(.A(new_n412), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n350), .B1(new_n388), .B2(KEYINPUT13), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n415), .B1(new_n416), .B2(new_n391), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n413), .B1(new_n414), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n375), .A2(new_n245), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n419), .B(new_n370), .C1(G179), .C2(new_n375), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n368), .A2(G77), .ZN(new_n421));
  XNOR2_X1  g0221(.A(KEYINPUT15), .B(G87), .ZN(new_n422));
  OAI22_X1  g0222(.A1(new_n422), .A2(new_n360), .B1(new_n207), .B2(new_n402), .ZN(new_n423));
  INV_X1    g0223(.A(new_n359), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n423), .B1(new_n357), .B2(new_n424), .ZN(new_n425));
  OAI221_X1 g0225(.A(new_n421), .B1(G77), .B2(new_n278), .C1(new_n425), .C2(new_n283), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n336), .A2(G238), .B1(new_n335), .B2(G107), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n306), .A2(G232), .A3(new_n260), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n246), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n342), .B1(new_n343), .B2(G244), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n426), .B1(new_n433), .B2(G169), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n432), .A2(G179), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n433), .A2(G190), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n426), .B1(new_n432), .B2(G200), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT73), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n304), .A2(new_n207), .A3(new_n305), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT7), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT7), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n304), .A2(new_n443), .A3(new_n207), .A4(new_n305), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n442), .A2(G68), .A3(new_n444), .ZN(new_n445));
  XNOR2_X1  g0245(.A(G58), .B(G68), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n446), .A2(G20), .B1(G159), .B2(new_n357), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n445), .A2(KEYINPUT16), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT16), .B1(new_n445), .B2(new_n447), .ZN(new_n449));
  NOR3_X1   g0249(.A1(new_n448), .A2(new_n449), .A3(new_n283), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n359), .B1(new_n247), .B2(G20), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n451), .A2(new_n291), .B1(new_n290), .B2(new_n359), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n440), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n445), .A2(new_n447), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT16), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n445), .A2(KEYINPUT16), .A3(new_n447), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n457), .A2(new_n282), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n459), .A2(KEYINPUT73), .A3(new_n452), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n266), .A2(G232), .A3(new_n339), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n341), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  OR2_X1    g0263(.A1(G223), .A2(G1698), .ZN(new_n464));
  INV_X1    g0264(.A(G226), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G1698), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n464), .B(new_n466), .C1(new_n257), .C2(new_n258), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G87), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n246), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n245), .B1(new_n463), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n266), .B1(new_n467), .B2(new_n468), .ZN(new_n472));
  INV_X1    g0272(.A(G179), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n472), .A2(new_n462), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n454), .A2(new_n460), .A3(new_n476), .ZN(new_n477));
  OR2_X1    g0277(.A1(new_n477), .A2(KEYINPUT18), .ZN(new_n478));
  INV_X1    g0278(.A(G200), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n479), .B1(new_n463), .B2(new_n470), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n472), .A2(new_n462), .A3(new_n350), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n459), .A2(new_n482), .A3(new_n452), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT17), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n283), .B1(new_n455), .B2(new_n456), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n453), .B1(new_n486), .B2(new_n458), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(KEYINPUT17), .A3(new_n482), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n489), .B1(KEYINPUT18), .B2(new_n477), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n439), .A2(new_n478), .A3(new_n490), .ZN(new_n491));
  AND4_X1   g0291(.A1(new_n381), .A2(new_n418), .A3(new_n420), .A4(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT75), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT74), .ZN(new_n494));
  OAI211_X1 g0294(.A(G244), .B(new_n260), .C1(new_n257), .C2(new_n258), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT4), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n332), .A2(KEYINPUT74), .A3(KEYINPUT4), .A4(G244), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n495), .A2(new_n496), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G33), .A2(G283), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n306), .A2(G250), .A3(G1698), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n493), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n503), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n497), .A2(new_n498), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n505), .A2(KEYINPUT75), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n504), .A2(new_n246), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n256), .A2(G257), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n267), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n508), .A2(new_n473), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n286), .A2(KEYINPUT6), .A3(G97), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n236), .B2(KEYINPUT6), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n514), .A2(G20), .B1(G77), .B2(new_n357), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n442), .A2(G107), .A3(new_n444), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n283), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(G97), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n290), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(new_n285), .B2(new_n518), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n505), .A2(new_n506), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n266), .B1(new_n523), .B2(new_n493), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n510), .B1(new_n524), .B2(new_n507), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n512), .B(new_n522), .C1(new_n525), .C2(G169), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n508), .A2(G190), .A3(new_n511), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n527), .B(new_n521), .C1(new_n525), .C2(new_n479), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(G264), .B(G1698), .C1(new_n257), .C2(new_n258), .ZN(new_n530));
  OAI211_X1 g0330(.A(G257), .B(new_n260), .C1(new_n257), .C2(new_n258), .ZN(new_n531));
  INV_X1    g0331(.A(G303), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n530), .B(new_n531), .C1(new_n532), .C2(new_n306), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n246), .ZN(new_n534));
  OAI211_X1 g0334(.A(G270), .B(new_n266), .C1(new_n270), .C2(new_n274), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n534), .A2(new_n267), .A3(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(G116), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n290), .A2(KEYINPUT82), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT82), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n278), .B2(G116), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n281), .A2(new_n208), .B1(G20), .B2(new_n537), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n501), .B(new_n207), .C1(G33), .C2(new_n518), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n542), .A2(KEYINPUT20), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT20), .B1(new_n542), .B2(new_n543), .ZN(new_n545));
  OAI221_X1 g0345(.A(new_n541), .B1(new_n285), .B2(new_n537), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n536), .A2(new_n546), .A3(G169), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT83), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT21), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT21), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n547), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n546), .B1(new_n536), .B2(G200), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n350), .B2(new_n536), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n536), .A2(new_n473), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n546), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n550), .A2(new_n552), .A3(new_n554), .A4(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n360), .A2(new_n518), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT19), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT78), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT78), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT19), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(KEYINPUT80), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  XNOR2_X1  g0364(.A(KEYINPUT78), .B(KEYINPUT19), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT80), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n565), .B(new_n566), .C1(new_n518), .C2(new_n360), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n306), .A2(new_n207), .A3(G68), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n564), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n383), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n563), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g0371(.A(KEYINPUT79), .B(G87), .Z(new_n572));
  NOR2_X1   g0372(.A1(G97), .A2(G107), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n571), .A2(new_n207), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n282), .B1(new_n569), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n422), .A2(new_n290), .ZN(new_n576));
  INV_X1    g0376(.A(new_n285), .ZN(new_n577));
  INV_X1    g0377(.A(new_n422), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n575), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT81), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT81), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n575), .A2(new_n582), .A3(new_n576), .A4(new_n579), .ZN(new_n583));
  OAI211_X1 g0383(.A(G238), .B(new_n260), .C1(new_n257), .C2(new_n258), .ZN(new_n584));
  OAI211_X1 g0384(.A(G244), .B(G1698), .C1(new_n257), .C2(new_n258), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n584), .B(new_n585), .C1(new_n265), .C2(new_n537), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n246), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n248), .A2(G250), .ZN(new_n588));
  OAI21_X1  g0388(.A(KEYINPUT77), .B1(new_n246), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT77), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n266), .A2(new_n590), .A3(G250), .A4(new_n248), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n589), .A2(new_n591), .B1(G274), .B2(new_n272), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(G169), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n587), .A2(new_n592), .A3(G179), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n581), .A2(new_n583), .A3(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n593), .A2(new_n350), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n479), .B1(new_n587), .B2(new_n592), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n577), .A2(G87), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n575), .A2(new_n576), .A3(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n597), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n557), .A2(new_n605), .ZN(new_n606));
  AND4_X1   g0406(.A1(new_n330), .A2(new_n492), .A3(new_n529), .A4(new_n606), .ZN(G372));
  AND3_X1   g0407(.A1(new_n587), .A2(new_n592), .A3(G179), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n245), .B1(new_n587), .B2(new_n592), .ZN(new_n609));
  OAI21_X1  g0409(.A(KEYINPUT87), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT87), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n594), .A2(new_n611), .A3(new_n595), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n612), .A3(new_n580), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n613), .A2(new_n325), .A3(new_n604), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n315), .A2(new_n316), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n313), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n550), .A2(new_n616), .A3(new_n552), .A4(new_n556), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n614), .A2(new_n526), .A3(new_n528), .A4(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n618), .A2(new_n613), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n580), .A2(KEYINPUT81), .B1(new_n594), .B2(new_n595), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n620), .A2(new_n583), .B1(new_n600), .B2(new_n603), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n508), .A2(new_n511), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n521), .B1(new_n622), .B2(new_n245), .ZN(new_n623));
  XNOR2_X1  g0423(.A(KEYINPUT88), .B(KEYINPUT26), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n621), .A2(new_n623), .A3(new_n512), .A4(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT89), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n508), .A2(new_n473), .A3(new_n511), .ZN(new_n629));
  AOI21_X1  g0429(.A(G169), .B1(new_n508), .B2(new_n511), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n629), .A2(new_n630), .A3(new_n521), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n631), .A2(KEYINPUT89), .A3(new_n621), .A4(new_n625), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT26), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n613), .A2(new_n604), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n633), .B1(new_n526), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n628), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n619), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n492), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n420), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n475), .B1(new_n459), .B2(new_n452), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n640), .B(KEYINPUT18), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n414), .A2(new_n417), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n413), .B1(new_n642), .B2(new_n436), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n641), .B1(new_n643), .B2(new_n489), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n639), .B1(new_n644), .B2(new_n381), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n638), .A2(new_n645), .ZN(G369));
  NAND3_X1  g0446(.A1(new_n247), .A2(new_n207), .A3(G13), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(new_n649), .A3(G213), .ZN(new_n650));
  INV_X1    g0450(.A(G343), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n319), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n313), .A2(new_n652), .ZN(new_n656));
  AOI21_X1  g0456(.A(KEYINPUT91), .B1(new_n330), .B2(new_n656), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n319), .A2(new_n328), .A3(new_n325), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n328), .B1(new_n319), .B2(new_n325), .ZN(new_n659));
  OAI211_X1 g0459(.A(KEYINPUT91), .B(new_n656), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n655), .B1(new_n657), .B2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n552), .A2(new_n556), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n550), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n546), .A2(new_n652), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n557), .B2(new_n665), .ZN(new_n667));
  XOR2_X1   g0467(.A(KEYINPUT90), .B(G330), .Z(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n662), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n313), .A2(new_n615), .A3(new_n653), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n656), .B1(new_n658), .B2(new_n659), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT91), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n652), .B1(new_n663), .B2(new_n550), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(new_n660), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n672), .A2(new_n673), .A3(new_n678), .ZN(G399));
  NOR2_X1   g0479(.A1(new_n213), .A2(G41), .ZN(new_n680));
  INV_X1    g0480(.A(new_n206), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n572), .A2(new_n573), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(G116), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G1), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n682), .B1(new_n680), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT28), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT29), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n637), .A2(new_n688), .A3(new_n653), .ZN(new_n689));
  NOR3_X1   g0489(.A1(new_n602), .A2(new_n598), .A3(new_n599), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n565), .A2(new_n383), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n683), .B1(new_n691), .B2(G20), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n692), .A2(new_n568), .A3(new_n564), .A4(new_n567), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n693), .A2(new_n282), .B1(new_n290), .B2(new_n422), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n596), .A2(KEYINPUT87), .B1(new_n694), .B2(new_n579), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n690), .B1(new_n695), .B2(new_n612), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n696), .A2(KEYINPUT26), .A3(new_n512), .A4(new_n623), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT95), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n624), .B1(new_n526), .B2(new_n605), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT96), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI211_X1 g0502(.A(KEYINPUT96), .B(new_n624), .C1(new_n526), .C2(new_n605), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n631), .A2(KEYINPUT95), .A3(KEYINPUT26), .A4(new_n696), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n699), .A2(new_n702), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n663), .A2(new_n319), .A3(new_n550), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n706), .A2(new_n614), .A3(new_n526), .A4(new_n528), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n707), .A2(new_n613), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n652), .B1(new_n705), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n689), .B1(new_n709), .B2(new_n688), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n330), .A2(new_n529), .A3(new_n606), .A4(new_n653), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT31), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n587), .A2(new_n592), .A3(KEYINPUT92), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(new_n536), .A3(new_n473), .ZN(new_n714));
  AOI21_X1  g0514(.A(KEYINPUT92), .B1(new_n587), .B2(new_n592), .ZN(new_n715));
  OAI21_X1  g0515(.A(KEYINPUT93), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n535), .A2(new_n267), .ZN(new_n717));
  AOI21_X1  g0517(.A(G179), .B1(new_n717), .B2(new_n534), .ZN(new_n718));
  INV_X1    g0518(.A(new_n715), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT93), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n718), .A2(new_n719), .A3(new_n720), .A4(new_n713), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n716), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n322), .B1(new_n508), .B2(new_n511), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT30), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n264), .A2(new_n587), .A3(new_n592), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n555), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n725), .B1(new_n622), .B2(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n525), .A2(KEYINPUT30), .A3(new_n555), .A4(new_n726), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n724), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n653), .B1(new_n730), .B2(KEYINPUT94), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT94), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n724), .A2(new_n732), .A3(new_n728), .A4(new_n729), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n712), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n730), .A2(KEYINPUT31), .A3(new_n652), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n668), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n710), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n687), .B1(new_n738), .B2(G1), .ZN(G364));
  NOR2_X1   g0539(.A1(new_n213), .A2(new_n306), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(new_n271), .B2(new_n681), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(new_n271), .B2(new_n243), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n213), .A2(new_n335), .ZN(new_n744));
  AOI22_X1  g0544(.A1(new_n744), .A2(G355), .B1(new_n537), .B2(new_n213), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(KEYINPUT97), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n745), .A2(KEYINPUT97), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n743), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n208), .B1(G20), .B2(new_n245), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XOR2_X1   g0553(.A(new_n753), .B(KEYINPUT98), .Z(new_n754));
  AND2_X1   g0554(.A1(new_n748), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(G13), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G20), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n247), .B1(new_n757), .B2(G45), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n680), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G179), .A2(G200), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n207), .B1(new_n762), .B2(G190), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G97), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n473), .A2(new_n479), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n207), .A2(G190), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n765), .B1(new_n202), .B2(new_n768), .ZN(new_n769));
  XOR2_X1   g0569(.A(new_n769), .B(KEYINPUT99), .Z(new_n770));
  NAND2_X1  g0570(.A1(new_n767), .A2(new_n762), .ZN(new_n771));
  INV_X1    g0571(.A(G159), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT32), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n207), .A2(new_n350), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n775), .A2(new_n473), .A3(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n473), .A2(G200), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n776), .A2(new_n572), .B1(new_n778), .B2(new_n201), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n767), .A2(new_n777), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n306), .B1(new_n780), .B2(new_n402), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n766), .A2(new_n775), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n238), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n767), .A2(new_n473), .A3(G200), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n286), .ZN(new_n785));
  NOR4_X1   g0585(.A1(new_n779), .A2(new_n781), .A3(new_n783), .A4(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n770), .A2(new_n774), .A3(new_n786), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT100), .Z(new_n788));
  XOR2_X1   g0588(.A(KEYINPUT33), .B(G317), .Z(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n768), .ZN(new_n790));
  INV_X1    g0590(.A(G283), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n335), .B1(new_n784), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n782), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n790), .B(new_n792), .C1(G326), .C2(new_n793), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n776), .B(KEYINPUT101), .Z(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G303), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n764), .A2(G294), .ZN(new_n797));
  INV_X1    g0597(.A(G322), .ZN(new_n798));
  INV_X1    g0598(.A(G311), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n778), .A2(new_n798), .B1(new_n780), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n771), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n800), .B1(G329), .B2(new_n801), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n794), .A2(new_n796), .A3(new_n797), .A4(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(KEYINPUT102), .B1(new_n788), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n752), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n788), .A2(KEYINPUT102), .A3(new_n803), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n755), .B(new_n761), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n751), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n808), .B1(new_n667), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n671), .A2(new_n760), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n669), .B2(new_n667), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n810), .A2(new_n812), .ZN(G396));
  AOI21_X1  g0613(.A(new_n652), .B1(new_n619), .B2(new_n636), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n436), .A2(new_n652), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(KEYINPUT103), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT103), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n436), .A2(new_n817), .A3(new_n652), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n426), .A2(new_n652), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n439), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n814), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n814), .A2(new_n822), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n711), .A2(KEYINPUT31), .B1(new_n731), .B2(new_n733), .ZN(new_n826));
  INV_X1    g0626(.A(new_n736), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n669), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n760), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n828), .B2(new_n825), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n805), .A2(new_n750), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n760), .B1(G77), .B2(new_n831), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n782), .A2(new_n532), .B1(new_n771), .B2(new_n799), .ZN(new_n833));
  INV_X1    g0633(.A(new_n780), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n306), .B(new_n833), .C1(G116), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n795), .A2(G107), .ZN(new_n836));
  INV_X1    g0636(.A(G87), .ZN(new_n837));
  INV_X1    g0637(.A(G294), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n837), .A2(new_n784), .B1(new_n778), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n768), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n839), .B1(G283), .B2(new_n840), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n835), .A2(new_n836), .A3(new_n765), .A4(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n778), .ZN(new_n843));
  AOI22_X1  g0643(.A1(G143), .A2(new_n843), .B1(new_n834), .B2(G159), .ZN(new_n844));
  INV_X1    g0644(.A(G137), .ZN(new_n845));
  INV_X1    g0645(.A(G150), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n844), .B1(new_n845), .B2(new_n782), .C1(new_n846), .C2(new_n768), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT34), .Z(new_n848));
  NOR2_X1   g0648(.A1(new_n784), .A2(new_n202), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n335), .B(new_n849), .C1(G132), .C2(new_n801), .ZN(new_n850));
  INV_X1    g0650(.A(new_n795), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n850), .B1(new_n201), .B2(new_n763), .C1(new_n851), .C2(new_n238), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n842), .B1(new_n848), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n832), .B1(new_n853), .B2(new_n752), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n822), .B2(new_n750), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n830), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(G384));
  NOR2_X1   g0657(.A1(new_n757), .A2(new_n247), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n731), .A2(KEYINPUT31), .A3(new_n733), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n735), .A2(new_n860), .B1(new_n821), .B2(new_n819), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT38), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n440), .B(new_n453), .C1(new_n486), .C2(new_n458), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT73), .B1(new_n459), .B2(new_n452), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n650), .ZN(new_n866));
  INV_X1    g0666(.A(new_n641), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n865), .B(new_n866), .C1(new_n867), .C2(new_n489), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n454), .A2(new_n460), .A3(new_n866), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT37), .B1(new_n487), .B2(new_n482), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n477), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT105), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n477), .A2(new_n870), .A3(KEYINPUT105), .A4(new_n871), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT107), .ZN(new_n876));
  INV_X1    g0676(.A(new_n483), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n876), .B1(new_n877), .B2(new_n640), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n459), .A2(new_n452), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n476), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n880), .A2(KEYINPUT107), .A3(new_n483), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n878), .A2(new_n881), .A3(new_n870), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n874), .A2(new_n875), .B1(KEYINPUT37), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n862), .B1(new_n869), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT104), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n877), .B2(new_n640), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n880), .A2(KEYINPUT104), .A3(new_n483), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n879), .A2(new_n866), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT37), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT37), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n483), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(new_n865), .B2(new_n476), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT105), .B1(new_n893), .B2(new_n870), .ZN(new_n894));
  INV_X1    g0694(.A(new_n875), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n890), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n888), .B1(new_n490), .B2(new_n478), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n896), .A2(new_n898), .A3(KEYINPUT38), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n884), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n415), .A2(new_n652), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n642), .B(new_n901), .C1(new_n400), .C2(new_n412), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n400), .A2(new_n901), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n861), .A2(new_n900), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT40), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT40), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n874), .A2(new_n875), .B1(KEYINPUT37), .B2(new_n889), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n862), .B1(new_n908), .B2(new_n897), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n899), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n861), .A2(new_n907), .A3(new_n910), .A4(new_n904), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n860), .A2(new_n735), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n492), .A2(new_n913), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n912), .B(new_n914), .Z(new_n915));
  NOR2_X1   g0715(.A1(new_n915), .A2(new_n668), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n413), .A2(new_n653), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT106), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT38), .B1(new_n896), .B2(new_n898), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n908), .A2(new_n862), .A3(new_n897), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n920), .B(KEYINPUT39), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT39), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n884), .A2(new_n899), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n924), .B1(new_n899), .B2(new_n909), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n927), .A2(new_n920), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n919), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n436), .A2(new_n653), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(new_n814), .B2(new_n822), .ZN(new_n932));
  INV_X1    g0732(.A(new_n904), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n934), .A2(new_n910), .B1(new_n867), .B2(new_n650), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n929), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n492), .A2(new_n710), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n645), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n936), .B(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n858), .B1(new_n917), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n939), .B2(new_n917), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n514), .A2(KEYINPUT35), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n514), .A2(KEYINPUT35), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n208), .A2(new_n207), .A3(new_n537), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT36), .ZN(new_n946));
  OAI21_X1  g0746(.A(G77), .B1(new_n201), .B2(new_n202), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n239), .B1(new_n206), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n948), .A2(G1), .A3(new_n756), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n941), .A2(new_n946), .A3(new_n949), .ZN(G367));
  NOR2_X1   g0750(.A1(new_n741), .A2(new_n233), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n753), .B1(new_n212), .B2(new_n422), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n760), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n335), .B1(new_n768), .B2(new_n838), .ZN(new_n954));
  INV_X1    g0754(.A(new_n776), .ZN(new_n955));
  AOI21_X1  g0755(.A(KEYINPUT46), .B1(new_n955), .B2(G116), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n954), .B(new_n956), .C1(G107), .C2(new_n764), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n795), .A2(KEYINPUT46), .A3(G116), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n784), .A2(new_n518), .B1(new_n780), .B2(new_n791), .ZN(new_n959));
  XNOR2_X1  g0759(.A(KEYINPUT112), .B(G317), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n959), .B1(new_n801), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n957), .A2(new_n958), .A3(new_n962), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n782), .A2(new_n799), .B1(new_n778), .B2(new_n532), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT111), .Z(new_n965));
  OAI22_X1  g0765(.A1(new_n776), .A2(new_n201), .B1(new_n778), .B2(new_n846), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(G68), .B2(new_n764), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n793), .A2(G143), .B1(new_n801), .B2(G137), .ZN(new_n968));
  AOI22_X1  g0768(.A1(G159), .A2(new_n840), .B1(new_n834), .B2(G50), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n784), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(G77), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n306), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT113), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n963), .A2(new_n965), .B1(new_n970), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT47), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n953), .B1(new_n976), .B2(new_n752), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n603), .A2(new_n653), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n695), .A2(new_n612), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n634), .B2(new_n978), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n977), .B1(new_n980), .B2(new_n809), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n631), .A2(new_n652), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n522), .A2(new_n652), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n526), .A2(new_n528), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n678), .A2(new_n673), .A3(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT45), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n986), .A2(new_n987), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n678), .A2(new_n673), .ZN(new_n990));
  INV_X1    g0790(.A(new_n985), .ZN(new_n991));
  AOI21_X1  g0791(.A(KEYINPUT44), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT44), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n993), .B(new_n985), .C1(new_n678), .C2(new_n673), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n988), .A2(new_n989), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n672), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n995), .A2(KEYINPUT110), .A3(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n677), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n655), .B(new_n998), .C1(new_n657), .C2(new_n661), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n999), .A2(new_n670), .A3(new_n678), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n670), .B1(new_n999), .B2(new_n678), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n828), .B(new_n689), .C1(new_n688), .C2(new_n709), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n996), .A2(KEYINPUT110), .ZN(new_n1005));
  NOR3_X1   g0805(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n672), .B1(new_n992), .B2(new_n994), .C1(new_n989), .C2(new_n988), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n997), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n738), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n680), .B(KEYINPUT41), .Z(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n759), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n672), .A2(new_n991), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n319), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n529), .A2(new_n1017), .A3(new_n983), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n652), .B1(new_n1018), .B2(new_n526), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n676), .A2(new_n660), .A3(new_n677), .A4(new_n985), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1019), .B1(new_n1020), .B2(KEYINPUT42), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n657), .A2(new_n661), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT42), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1022), .A2(new_n1023), .A3(new_n677), .A4(new_n985), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT108), .ZN(new_n1025));
  AND3_X1   g0825(.A1(new_n1021), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1025), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1016), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1020), .A2(KEYINPUT42), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1019), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1020), .A2(KEYINPUT42), .ZN(new_n1032));
  OAI21_X1  g0832(.A(KEYINPUT108), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n980), .B(KEYINPUT43), .Z(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1021), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT109), .ZN(new_n1038));
  AND3_X1   g0838(.A1(new_n1028), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1038), .B1(new_n1028), .B2(new_n1037), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1014), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NOR3_X1   g0841(.A1(new_n1026), .A2(new_n1027), .A3(new_n1034), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1015), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1043));
  OAI21_X1  g0843(.A(KEYINPUT109), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1028), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1044), .A2(new_n1013), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1041), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n981), .B1(new_n1012), .B2(new_n1047), .ZN(G387));
  NAND2_X1  g0848(.A1(new_n999), .A2(new_n678), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n671), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n1000), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n662), .A2(new_n809), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n782), .A2(new_n798), .B1(new_n768), .B2(new_n799), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n778), .A2(new_n960), .B1(new_n780), .B2(new_n532), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1055), .A2(KEYINPUT48), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(KEYINPUT48), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n955), .A2(G294), .B1(new_n764), .B2(G283), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT49), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n784), .A2(new_n537), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n306), .B(new_n1063), .C1(G326), .C2(new_n801), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1061), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n776), .A2(new_n402), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n306), .B1(new_n784), .B2(new_n518), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1066), .B(new_n1067), .C1(G159), .C2(new_n793), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G68), .A2(new_n834), .B1(new_n801), .B2(G150), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G50), .A2(new_n843), .B1(new_n840), .B2(new_n424), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n764), .A2(new_n578), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n805), .B1(new_n1065), .B2(new_n1072), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n230), .A2(new_n271), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n684), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1074), .A2(new_n740), .B1(new_n1075), .B2(new_n744), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n271), .B1(new_n202), .B2(new_n402), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT50), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n424), .B2(new_n238), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n359), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1080));
  NOR4_X1   g0880(.A1(new_n1075), .A2(new_n1077), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n1076), .A2(new_n1081), .B1(G107), .B2(new_n212), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n761), .B(new_n1073), .C1(new_n754), .C2(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n1051), .A2(new_n759), .B1(new_n1052), .B2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n680), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT114), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n1085), .A2(new_n1086), .B1(new_n738), .B2(new_n1051), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n680), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n738), .B2(new_n1051), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1089), .A2(KEYINPUT114), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1084), .B1(new_n1087), .B2(new_n1090), .ZN(G393));
  AND2_X1   g0891(.A1(new_n1008), .A2(new_n680), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT115), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n995), .A2(new_n1093), .A3(new_n996), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n1007), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1093), .B1(new_n995), .B2(new_n996), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n1095), .A2(new_n1096), .B1(new_n1004), .B2(new_n1003), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1092), .A2(new_n1097), .ZN(new_n1098));
  OR3_X1    g0898(.A1(new_n1095), .A2(new_n758), .A3(new_n1096), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT116), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n740), .A2(new_n237), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n753), .B1(new_n212), .B2(new_n518), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n760), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n306), .B(new_n785), .C1(G116), .C2(new_n764), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(G303), .A2(new_n840), .B1(new_n834), .B2(G294), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n955), .A2(G283), .B1(new_n801), .B2(G322), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G317), .A2(new_n793), .B1(new_n843), .B2(G311), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT52), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n782), .A2(new_n846), .B1(new_n778), .B2(new_n772), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT51), .Z(new_n1111));
  OAI21_X1  g0911(.A(new_n306), .B1(new_n784), .B2(new_n837), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G77), .B2(new_n764), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(G50), .A2(new_n840), .B1(new_n801), .B2(G143), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n955), .A2(G68), .B1(new_n834), .B2(new_n424), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n1107), .A2(new_n1109), .B1(new_n1111), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1103), .B1(new_n1117), .B2(new_n752), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n985), .B2(new_n809), .ZN(new_n1119));
  AND3_X1   g0919(.A1(new_n1099), .A2(new_n1100), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1100), .B1(new_n1099), .B2(new_n1119), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1098), .B1(new_n1120), .B2(new_n1121), .ZN(G390));
  OAI21_X1  g0922(.A(new_n918), .B1(new_n932), .B2(new_n933), .ZN(new_n1123));
  OAI21_X1  g0923(.A(KEYINPUT39), .B1(new_n921), .B2(new_n922), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(KEYINPUT106), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1123), .A2(new_n1125), .A3(new_n923), .A4(new_n925), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n737), .A2(new_n822), .A3(new_n904), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n931), .B1(new_n709), .B2(new_n822), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n918), .B(new_n900), .C1(new_n1128), .C2(new_n933), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1126), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n900), .A2(new_n918), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n709), .A2(new_n822), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n930), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1131), .B1(new_n1133), .B2(new_n904), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n926), .A2(new_n928), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1134), .B1(new_n1135), .B2(new_n1123), .ZN(new_n1136));
  OAI211_X1 g0936(.A(G330), .B(new_n822), .C1(new_n826), .C2(new_n859), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1137), .A2(new_n933), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1130), .B1(new_n1136), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1137), .A2(new_n933), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT117), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1137), .A2(KEYINPUT117), .A3(new_n933), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1143), .A2(new_n1127), .A3(new_n1128), .A4(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n932), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n904), .B1(new_n737), .B2(new_n822), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1146), .B1(new_n1147), .B2(new_n1138), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n492), .A2(G330), .A3(new_n913), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1150), .A2(new_n937), .A3(new_n645), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1088), .B1(new_n1140), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1151), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n1138), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1155), .A2(new_n1157), .A3(new_n1130), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1154), .A2(new_n1158), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n759), .B(new_n1130), .C1(new_n1136), .C2(new_n1139), .ZN(new_n1160));
  NOR3_X1   g0960(.A1(new_n926), .A2(new_n928), .A3(new_n750), .ZN(new_n1161));
  INV_X1    g0961(.A(G128), .ZN(new_n1162));
  INV_X1    g0962(.A(G132), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n782), .A2(new_n1162), .B1(new_n778), .B2(new_n1163), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n1164), .B(KEYINPUT118), .Z(new_n1165));
  AOI22_X1  g0965(.A1(new_n971), .A2(G50), .B1(new_n840), .B2(G137), .ZN(new_n1166));
  INV_X1    g0966(.A(G125), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1166), .B1(new_n1167), .B2(new_n771), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT54), .B(G143), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n776), .A2(new_n846), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT53), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n306), .B1(new_n780), .B2(new_n1169), .C1(new_n1170), .C2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n772), .B2(new_n763), .ZN(new_n1174));
  NOR4_X1   g0974(.A1(new_n1165), .A2(new_n1168), .A3(new_n1172), .A4(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n306), .B1(new_n795), .B2(G87), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT119), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n849), .B1(G294), .B2(new_n801), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n402), .B2(new_n763), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n768), .A2(new_n286), .B1(new_n780), .B2(new_n518), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n782), .A2(new_n791), .B1(new_n778), .B2(new_n537), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1175), .B1(new_n1177), .B2(new_n1182), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n760), .B1(new_n424), .B2(new_n831), .C1(new_n1183), .C2(new_n805), .ZN(new_n1184));
  OAI21_X1  g0984(.A(KEYINPUT120), .B1(new_n1161), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n882), .A2(KEYINPUT37), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n894), .B2(new_n895), .ZN(new_n1187));
  AOI21_X1  g0987(.A(KEYINPUT38), .B1(new_n1187), .B2(new_n868), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1188), .A2(new_n922), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n920), .A2(new_n927), .B1(new_n1189), .B2(new_n924), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1190), .A2(new_n749), .A3(new_n1125), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT120), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1184), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1185), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1160), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1159), .A2(new_n1197), .ZN(G378));
  NAND2_X1  g0998(.A1(new_n912), .A2(G330), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n381), .A2(new_n420), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n370), .A2(new_n866), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n381), .A2(new_n420), .A3(new_n1201), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1205), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1201), .B1(new_n381), .B2(new_n420), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1202), .B(new_n639), .C1(new_n377), .C2(new_n380), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1207), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1206), .A2(new_n1210), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n929), .A2(new_n935), .A3(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1211), .B1(new_n929), .B2(new_n935), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1199), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1211), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n918), .B1(new_n1190), .B2(new_n1125), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n934), .A2(new_n910), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n867), .A2(new_n650), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1215), .B1(new_n1216), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(G330), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n906), .B2(new_n911), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n929), .A2(new_n935), .A3(new_n1211), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1220), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1214), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1215), .A2(new_n749), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n760), .B1(G50), .B2(new_n831), .ZN(new_n1227));
  AOI21_X1  g1027(.A(G50), .B1(new_n305), .B2(new_n252), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n784), .A2(new_n201), .B1(new_n771), .B2(new_n791), .ZN(new_n1229));
  NOR4_X1   g1029(.A1(new_n1229), .A2(new_n1066), .A3(G41), .A4(new_n306), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n764), .A2(G68), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n793), .A2(G116), .B1(new_n834), .B2(new_n578), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(G97), .A2(new_n840), .B1(new_n843), .B2(G107), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .A4(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT58), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1228), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  AOI211_X1 g1036(.A(G33), .B(G41), .C1(new_n971), .C2(G159), .ZN(new_n1237));
  XOR2_X1   g1037(.A(KEYINPUT122), .B(G124), .Z(new_n1238));
  OAI22_X1  g1038(.A1(new_n776), .A2(new_n1169), .B1(new_n778), .B2(new_n1162), .ZN(new_n1239));
  XOR2_X1   g1039(.A(new_n1239), .B(KEYINPUT121), .Z(new_n1240));
  NOR2_X1   g1040(.A1(new_n768), .A2(new_n1163), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n782), .A2(new_n1167), .B1(new_n780), .B2(new_n845), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(G150), .C2(new_n764), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1240), .A2(new_n1243), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1237), .B1(new_n771), .B2(new_n1238), .C1(new_n1244), .C2(KEYINPUT59), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1244), .A2(KEYINPUT59), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n1236), .B1(new_n1235), .B2(new_n1234), .C1(new_n1245), .C2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1227), .B1(new_n1247), .B2(new_n752), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n1225), .A2(new_n759), .B1(new_n1226), .B2(new_n1248), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1224), .A2(new_n1214), .B1(new_n1158), .B2(new_n1152), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n680), .B1(new_n1250), .B2(KEYINPUT57), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1149), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1152), .B1(new_n1140), .B2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1225), .A2(new_n1253), .A3(KEYINPUT57), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1249), .B1(new_n1251), .B2(new_n1255), .ZN(G375));
  NAND2_X1  g1056(.A1(new_n933), .A2(new_n749), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n760), .B1(G68), .B2(new_n831), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(G150), .A2(new_n834), .B1(new_n801), .B2(G128), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n335), .B1(new_n971), .B2(G58), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1259), .B(new_n1260), .C1(new_n238), .C2(new_n763), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1169), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n793), .A2(G132), .B1(new_n840), .B2(new_n1262), .ZN(new_n1263));
  OAI221_X1 g1063(.A(new_n1263), .B1(new_n845), .B2(new_n778), .C1(new_n851), .C2(new_n772), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(G116), .A2(new_n840), .B1(new_n834), .B2(G107), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n1265), .B1(new_n791), .B2(new_n778), .C1(new_n851), .C2(new_n518), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n793), .A2(G294), .B1(new_n801), .B2(G303), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1267), .A2(new_n335), .A3(new_n972), .A4(new_n1071), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n1261), .A2(new_n1264), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT123), .ZN(new_n1270));
  OR2_X1    g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n805), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1258), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1149), .A2(new_n759), .B1(new_n1257), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1153), .A2(new_n1011), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1274), .B1(new_n1275), .B2(new_n1276), .ZN(G381));
  NAND2_X1  g1077(.A1(new_n1225), .A2(new_n759), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1226), .A2(new_n1248), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1225), .A2(new_n1253), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT57), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1088), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  AOI211_X1 g1083(.A(G378), .B(new_n1280), .C1(new_n1283), .C2(new_n1254), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1121), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1099), .A2(new_n1100), .A3(new_n1119), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(new_n1285), .A2(new_n1286), .B1(new_n1097), .B2(new_n1092), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1084), .ZN(new_n1288));
  AOI22_X1  g1088(.A1(new_n1089), .A2(KEYINPUT114), .B1(new_n1004), .B2(new_n1003), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1290));
  AOI211_X1 g1090(.A(G396), .B(new_n1288), .C1(new_n1289), .C2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n856), .ZN(new_n1292));
  NOR3_X1   g1092(.A1(G387), .A2(G381), .A3(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1284), .A2(new_n1287), .A3(new_n1293), .ZN(G407));
  NAND2_X1  g1094(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1295), .A2(new_n680), .A3(new_n1254), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1196), .B1(new_n1154), .B2(new_n1158), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1296), .A2(new_n1297), .A3(new_n1249), .ZN(new_n1298));
  OAI211_X1 g1098(.A(G407), .B(G213), .C1(G343), .C2(new_n1298), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1299), .B(KEYINPUT124), .ZN(G409));
  NAND3_X1  g1100(.A1(new_n1225), .A2(new_n1253), .A3(new_n1011), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1249), .A2(new_n1297), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n651), .A2(G213), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1145), .A2(new_n1148), .A3(new_n1151), .A4(KEYINPUT60), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n680), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1153), .A2(KEYINPUT60), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1276), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1306), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1274), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n856), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1276), .B1(KEYINPUT60), .B2(new_n1153), .ZN(new_n1312));
  OAI211_X1 g1112(.A(G384), .B(new_n1274), .C1(new_n1312), .C2(new_n1306), .ZN(new_n1313));
  AND2_X1   g1113(.A1(new_n1311), .A2(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1280), .B1(new_n1283), .B2(new_n1254), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n1304), .B(new_n1314), .C1(new_n1297), .C2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(KEYINPUT62), .ZN(new_n1317));
  OR2_X1    g1117(.A1(new_n1303), .A2(KEYINPUT125), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n651), .A2(G213), .A3(G2897), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1314), .A2(new_n1318), .A3(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1311), .A2(new_n1313), .A3(new_n1318), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1319), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1297), .B1(new_n1296), .B2(new_n1249), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1325));
  OAI211_X1 g1125(.A(new_n1320), .B(new_n1323), .C1(new_n1324), .C2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT61), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(G375), .A2(G378), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT62), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1328), .A2(new_n1329), .A3(new_n1304), .A4(new_n1314), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1317), .A2(new_n1326), .A3(new_n1327), .A4(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(G396), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1332), .B1(new_n1333), .B2(new_n1084), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1334), .A2(new_n1291), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1335), .B1(G387), .B2(KEYINPUT126), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(G393), .A2(G396), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1333), .A2(new_n1332), .A3(new_n1084), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1010), .B1(new_n1008), .B2(new_n738), .ZN(new_n1340));
  OAI211_X1 g1140(.A(new_n1046), .B(new_n1041), .C1(new_n1340), .C2(new_n759), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1339), .B1(new_n1341), .B2(new_n981), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1287), .B1(new_n1336), .B2(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(G387), .A2(new_n1335), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT126), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1345), .B1(new_n1341), .B2(new_n981), .ZN(new_n1346));
  OAI211_X1 g1146(.A(G390), .B(new_n1344), .C1(new_n1335), .C2(new_n1346), .ZN(new_n1347));
  AND2_X1   g1147(.A1(new_n1343), .A2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1331), .A2(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT63), .ZN(new_n1350));
  AOI21_X1  g1150(.A(new_n1348), .B1(new_n1350), .B2(new_n1316), .ZN(new_n1351));
  NAND4_X1  g1151(.A1(new_n1328), .A2(KEYINPUT63), .A3(new_n1304), .A4(new_n1314), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1351), .A2(new_n1327), .A3(new_n1326), .A4(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1349), .A2(new_n1353), .ZN(G405));
  INV_X1    g1154(.A(new_n1314), .ZN(new_n1355));
  OAI21_X1  g1155(.A(new_n1355), .B1(new_n1284), .B2(new_n1324), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1328), .A2(new_n1298), .A3(new_n1314), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1356), .A2(new_n1357), .A3(new_n1348), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1348), .B1(new_n1356), .B2(new_n1357), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1358), .B1(new_n1359), .B2(KEYINPUT127), .ZN(new_n1360));
  INV_X1    g1160(.A(KEYINPUT127), .ZN(new_n1361));
  AOI211_X1 g1161(.A(new_n1361), .B(new_n1348), .C1(new_n1357), .C2(new_n1356), .ZN(new_n1362));
  NOR2_X1   g1162(.A1(new_n1360), .A2(new_n1362), .ZN(G402));
endmodule


