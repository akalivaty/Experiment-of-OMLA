

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581;

  XOR2_X1 U319 ( .A(n305), .B(n304), .Z(n450) );
  AND2_X1 U320 ( .A1(n554), .A2(n549), .ZN(n367) );
  XNOR2_X1 U321 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n413) );
  XNOR2_X1 U322 ( .A(n414), .B(n413), .ZN(n519) );
  XOR2_X1 U323 ( .A(n349), .B(KEYINPUT41), .Z(n554) );
  XOR2_X1 U324 ( .A(n366), .B(n387), .Z(n549) );
  XNOR2_X1 U325 ( .A(n447), .B(G204GAT), .ZN(n448) );
  XNOR2_X1 U326 ( .A(n449), .B(n448), .ZN(G1353GAT) );
  XOR2_X1 U327 ( .A(KEYINPUT72), .B(KEYINPUT75), .Z(n288) );
  XNOR2_X1 U328 ( .A(KEYINPUT33), .B(KEYINPUT77), .ZN(n287) );
  XNOR2_X1 U329 ( .A(n288), .B(n287), .ZN(n305) );
  XOR2_X1 U330 ( .A(G120GAT), .B(G71GAT), .Z(n336) );
  XNOR2_X1 U331 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n289) );
  XNOR2_X1 U332 ( .A(n289), .B(KEYINPUT13), .ZN(n374) );
  XOR2_X1 U333 ( .A(n336), .B(n374), .Z(n291) );
  NAND2_X1 U334 ( .A1(G230GAT), .A2(G233GAT), .ZN(n290) );
  XNOR2_X1 U335 ( .A(n291), .B(n290), .ZN(n298) );
  XOR2_X1 U336 ( .A(KEYINPUT76), .B(KEYINPUT31), .Z(n293) );
  XNOR2_X1 U337 ( .A(KEYINPUT74), .B(KEYINPUT32), .ZN(n292) );
  XNOR2_X1 U338 ( .A(n293), .B(n292), .ZN(n294) );
  XNOR2_X1 U339 ( .A(n294), .B(KEYINPUT71), .ZN(n296) );
  XOR2_X1 U340 ( .A(G176GAT), .B(G64GAT), .Z(n420) );
  XNOR2_X1 U341 ( .A(G204GAT), .B(n420), .ZN(n295) );
  XNOR2_X1 U342 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U343 ( .A(n298), .B(n297), .ZN(n303) );
  XNOR2_X1 U344 ( .A(G106GAT), .B(G78GAT), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n299), .B(G148GAT), .ZN(n311) );
  XOR2_X1 U346 ( .A(G92GAT), .B(KEYINPUT73), .Z(n301) );
  XNOR2_X1 U347 ( .A(G99GAT), .B(G85GAT), .ZN(n300) );
  XNOR2_X1 U348 ( .A(n301), .B(n300), .ZN(n396) );
  XNOR2_X1 U349 ( .A(n311), .B(n396), .ZN(n302) );
  XNOR2_X1 U350 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U351 ( .A(KEYINPUT90), .B(KEYINPUT22), .Z(n307) );
  NAND2_X1 U352 ( .A1(G228GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U353 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U354 ( .A(n308), .B(KEYINPUT23), .Z(n313) );
  XOR2_X1 U355 ( .A(G155GAT), .B(KEYINPUT3), .Z(n310) );
  XNOR2_X1 U356 ( .A(KEYINPUT2), .B(KEYINPUT91), .ZN(n309) );
  XNOR2_X1 U357 ( .A(n310), .B(n309), .ZN(n438) );
  XNOR2_X1 U358 ( .A(n438), .B(n311), .ZN(n312) );
  XNOR2_X1 U359 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U360 ( .A(KEYINPUT94), .B(KEYINPUT24), .Z(n315) );
  XNOR2_X1 U361 ( .A(KEYINPUT92), .B(KEYINPUT93), .ZN(n314) );
  XNOR2_X1 U362 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U363 ( .A(n317), .B(n316), .Z(n319) );
  XOR2_X1 U364 ( .A(G141GAT), .B(G22GAT), .Z(n352) );
  XOR2_X1 U365 ( .A(G50GAT), .B(G162GAT), .Z(n392) );
  XNOR2_X1 U366 ( .A(n352), .B(n392), .ZN(n318) );
  XNOR2_X1 U367 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U368 ( .A(G211GAT), .B(G218GAT), .Z(n321) );
  XNOR2_X1 U369 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n320) );
  XNOR2_X1 U370 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U371 ( .A(G197GAT), .B(n322), .Z(n421) );
  XOR2_X1 U372 ( .A(n323), .B(n421), .Z(n546) );
  XOR2_X1 U373 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n325) );
  XNOR2_X1 U374 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n324) );
  XNOR2_X1 U375 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U376 ( .A(KEYINPUT87), .B(n326), .ZN(n424) );
  XOR2_X1 U377 ( .A(KEYINPUT0), .B(G134GAT), .Z(n328) );
  XNOR2_X1 U378 ( .A(KEYINPUT85), .B(G127GAT), .ZN(n327) );
  XNOR2_X1 U379 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U380 ( .A(G113GAT), .B(n329), .ZN(n444) );
  XNOR2_X1 U381 ( .A(n424), .B(n444), .ZN(n343) );
  XOR2_X1 U382 ( .A(KEYINPUT89), .B(G190GAT), .Z(n331) );
  XNOR2_X1 U383 ( .A(G43GAT), .B(G99GAT), .ZN(n330) );
  XNOR2_X1 U384 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U385 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n333) );
  XNOR2_X1 U386 ( .A(G15GAT), .B(KEYINPUT88), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U388 ( .A(n335), .B(n334), .Z(n341) );
  XOR2_X1 U389 ( .A(n336), .B(G176GAT), .Z(n338) );
  NAND2_X1 U390 ( .A1(G227GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U391 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U392 ( .A(G169GAT), .B(n339), .ZN(n340) );
  XNOR2_X1 U393 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U394 ( .A(n343), .B(n342), .Z(n562) );
  INV_X1 U395 ( .A(n562), .ZN(n548) );
  NAND2_X1 U396 ( .A1(n546), .A2(n548), .ZN(n344) );
  XNOR2_X1 U397 ( .A(n344), .B(KEYINPUT26), .ZN(n536) );
  NAND2_X1 U398 ( .A1(n450), .A2(KEYINPUT65), .ZN(n348) );
  INV_X1 U399 ( .A(n450), .ZN(n346) );
  INV_X1 U400 ( .A(KEYINPUT65), .ZN(n345) );
  NAND2_X1 U401 ( .A1(n346), .A2(n345), .ZN(n347) );
  NAND2_X1 U402 ( .A1(n348), .A2(n347), .ZN(n349) );
  XOR2_X1 U403 ( .A(G15GAT), .B(G1GAT), .Z(n371) );
  XOR2_X1 U404 ( .A(G169GAT), .B(G8GAT), .Z(n415) );
  XOR2_X1 U405 ( .A(n371), .B(n415), .Z(n351) );
  NAND2_X1 U406 ( .A1(G229GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U407 ( .A(n351), .B(n350), .ZN(n353) );
  XOR2_X1 U408 ( .A(n353), .B(n352), .Z(n361) );
  XOR2_X1 U409 ( .A(G197GAT), .B(G113GAT), .Z(n355) );
  XNOR2_X1 U410 ( .A(G50GAT), .B(G36GAT), .ZN(n354) );
  XNOR2_X1 U411 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U412 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n357) );
  XNOR2_X1 U413 ( .A(KEYINPUT66), .B(KEYINPUT69), .ZN(n356) );
  XNOR2_X1 U414 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U415 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U416 ( .A(n361), .B(n360), .ZN(n366) );
  XOR2_X1 U417 ( .A(G29GAT), .B(KEYINPUT68), .Z(n363) );
  XNOR2_X1 U418 ( .A(G43GAT), .B(KEYINPUT67), .ZN(n362) );
  XNOR2_X1 U419 ( .A(n363), .B(n362), .ZN(n365) );
  XOR2_X1 U420 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n364) );
  XOR2_X1 U421 ( .A(n365), .B(n364), .Z(n387) );
  XNOR2_X1 U422 ( .A(n367), .B(KEYINPUT46), .ZN(n405) );
  XOR2_X1 U423 ( .A(G155GAT), .B(G71GAT), .Z(n369) );
  XNOR2_X1 U424 ( .A(G183GAT), .B(G127GAT), .ZN(n368) );
  XNOR2_X1 U425 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U426 ( .A(n370), .B(G78GAT), .Z(n373) );
  XNOR2_X1 U427 ( .A(G22GAT), .B(n371), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n378) );
  XOR2_X1 U429 ( .A(n374), .B(KEYINPUT12), .Z(n376) );
  NAND2_X1 U430 ( .A1(G231GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U431 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U432 ( .A(n378), .B(n377), .Z(n386) );
  XOR2_X1 U433 ( .A(KEYINPUT83), .B(G64GAT), .Z(n380) );
  XNOR2_X1 U434 ( .A(G8GAT), .B(G211GAT), .ZN(n379) );
  XNOR2_X1 U435 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U436 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n382) );
  XNOR2_X1 U437 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n381) );
  XNOR2_X1 U438 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U439 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U440 ( .A(n386), .B(n385), .Z(n574) );
  INV_X1 U441 ( .A(n387), .ZN(n391) );
  XOR2_X1 U442 ( .A(KEYINPUT78), .B(KEYINPUT9), .Z(n389) );
  XNOR2_X1 U443 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U445 ( .A(n391), .B(n390), .Z(n403) );
  XOR2_X1 U446 ( .A(G36GAT), .B(G190GAT), .Z(n418) );
  XOR2_X1 U447 ( .A(n418), .B(n392), .Z(n394) );
  XNOR2_X1 U448 ( .A(G218GAT), .B(G106GAT), .ZN(n393) );
  XNOR2_X1 U449 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U450 ( .A(n395), .B(KEYINPUT79), .Z(n401) );
  XOR2_X1 U451 ( .A(n396), .B(KEYINPUT80), .Z(n398) );
  NAND2_X1 U452 ( .A1(G232GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U453 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U454 ( .A(G134GAT), .B(n399), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U456 ( .A(n403), .B(n402), .Z(n561) );
  INV_X1 U457 ( .A(n561), .ZN(n463) );
  NAND2_X1 U458 ( .A1(n574), .A2(n463), .ZN(n404) );
  OR2_X1 U459 ( .A1(n405), .A2(n404), .ZN(n406) );
  XNOR2_X1 U460 ( .A(n406), .B(KEYINPUT47), .ZN(n412) );
  XNOR2_X1 U461 ( .A(KEYINPUT36), .B(KEYINPUT103), .ZN(n407) );
  XOR2_X1 U462 ( .A(n407), .B(n463), .Z(n578) );
  NOR2_X1 U463 ( .A1(n578), .A2(n574), .ZN(n408) );
  XNOR2_X1 U464 ( .A(KEYINPUT45), .B(n408), .ZN(n409) );
  NAND2_X1 U465 ( .A1(n409), .A2(n450), .ZN(n410) );
  NOR2_X1 U466 ( .A1(n410), .A2(n549), .ZN(n411) );
  NOR2_X1 U467 ( .A1(n412), .A2(n411), .ZN(n414) );
  XOR2_X1 U468 ( .A(G92GAT), .B(n415), .Z(n417) );
  NAND2_X1 U469 ( .A1(G226GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U470 ( .A(n417), .B(n416), .ZN(n419) );
  XOR2_X1 U471 ( .A(n419), .B(n418), .Z(n423) );
  XNOR2_X1 U472 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U473 ( .A(n423), .B(n422), .ZN(n425) );
  XOR2_X1 U474 ( .A(n425), .B(n424), .Z(n511) );
  INV_X1 U475 ( .A(n511), .ZN(n487) );
  NOR2_X1 U476 ( .A1(n519), .A2(n487), .ZN(n426) );
  XNOR2_X1 U477 ( .A(n426), .B(KEYINPUT54), .ZN(n445) );
  XOR2_X1 U478 ( .A(KEYINPUT96), .B(KEYINPUT6), .Z(n428) );
  XNOR2_X1 U479 ( .A(KEYINPUT5), .B(KEYINPUT95), .ZN(n427) );
  XNOR2_X1 U480 ( .A(n428), .B(n427), .ZN(n442) );
  XOR2_X1 U481 ( .A(G148GAT), .B(G120GAT), .Z(n430) );
  XNOR2_X1 U482 ( .A(G29GAT), .B(G141GAT), .ZN(n429) );
  XNOR2_X1 U483 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U484 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n432) );
  XNOR2_X1 U485 ( .A(G1GAT), .B(G57GAT), .ZN(n431) );
  XNOR2_X1 U486 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U487 ( .A(n434), .B(n433), .Z(n440) );
  XOR2_X1 U488 ( .A(G85GAT), .B(G162GAT), .Z(n436) );
  NAND2_X1 U489 ( .A1(G225GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U491 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U493 ( .A(n442), .B(n441), .Z(n443) );
  XOR2_X1 U494 ( .A(n444), .B(n443), .Z(n520) );
  INV_X1 U495 ( .A(n520), .ZN(n483) );
  NAND2_X1 U496 ( .A1(n445), .A2(n483), .ZN(n545) );
  NOR2_X1 U497 ( .A1(n536), .A2(n545), .ZN(n446) );
  XOR2_X1 U498 ( .A(KEYINPUT122), .B(n446), .Z(n579) );
  NOR2_X1 U499 ( .A1(n450), .A2(n579), .ZN(n449) );
  XNOR2_X1 U500 ( .A(KEYINPUT61), .B(KEYINPUT124), .ZN(n447) );
  NAND2_X1 U501 ( .A1(n549), .A2(n450), .ZN(n481) );
  XOR2_X1 U502 ( .A(n511), .B(KEYINPUT27), .Z(n518) );
  XOR2_X1 U503 ( .A(n546), .B(KEYINPUT28), .Z(n494) );
  INV_X1 U504 ( .A(n494), .ZN(n524) );
  NOR2_X1 U505 ( .A1(n518), .A2(n524), .ZN(n451) );
  NAND2_X1 U506 ( .A1(n451), .A2(n548), .ZN(n452) );
  NAND2_X1 U507 ( .A1(n520), .A2(n452), .ZN(n461) );
  NOR2_X1 U508 ( .A1(n548), .A2(n487), .ZN(n453) );
  NOR2_X1 U509 ( .A1(n546), .A2(n453), .ZN(n454) );
  XNOR2_X1 U510 ( .A(n454), .B(KEYINPUT97), .ZN(n455) );
  XNOR2_X1 U511 ( .A(n455), .B(KEYINPUT25), .ZN(n457) );
  NOR2_X1 U512 ( .A1(n536), .A2(n518), .ZN(n456) );
  NOR2_X1 U513 ( .A1(n457), .A2(n456), .ZN(n458) );
  XNOR2_X1 U514 ( .A(KEYINPUT98), .B(n458), .ZN(n459) );
  NAND2_X1 U515 ( .A1(n483), .A2(n459), .ZN(n460) );
  NAND2_X1 U516 ( .A1(n461), .A2(n460), .ZN(n462) );
  XNOR2_X1 U517 ( .A(KEYINPUT99), .B(n462), .ZN(n477) );
  XOR2_X1 U518 ( .A(KEYINPUT84), .B(KEYINPUT16), .Z(n465) );
  INV_X1 U519 ( .A(n574), .ZN(n557) );
  NAND2_X1 U520 ( .A1(n557), .A2(n463), .ZN(n464) );
  XNOR2_X1 U521 ( .A(n465), .B(n464), .ZN(n466) );
  NAND2_X1 U522 ( .A1(n477), .A2(n466), .ZN(n497) );
  NOR2_X1 U523 ( .A1(n481), .A2(n497), .ZN(n475) );
  NAND2_X1 U524 ( .A1(n520), .A2(n475), .ZN(n467) );
  XNOR2_X1 U525 ( .A(n467), .B(KEYINPUT34), .ZN(n468) );
  XOR2_X1 U526 ( .A(n468), .B(KEYINPUT101), .Z(n470) );
  XNOR2_X1 U527 ( .A(G1GAT), .B(KEYINPUT100), .ZN(n469) );
  XNOR2_X1 U528 ( .A(n470), .B(n469), .ZN(G1324GAT) );
  NAND2_X1 U529 ( .A1(n511), .A2(n475), .ZN(n471) );
  XNOR2_X1 U530 ( .A(n471), .B(KEYINPUT102), .ZN(n472) );
  XNOR2_X1 U531 ( .A(G8GAT), .B(n472), .ZN(G1325GAT) );
  XOR2_X1 U532 ( .A(G15GAT), .B(KEYINPUT35), .Z(n474) );
  NAND2_X1 U533 ( .A1(n475), .A2(n562), .ZN(n473) );
  XNOR2_X1 U534 ( .A(n474), .B(n473), .ZN(G1326GAT) );
  NAND2_X1 U535 ( .A1(n524), .A2(n475), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n476), .B(G22GAT), .ZN(G1327GAT) );
  XNOR2_X1 U537 ( .A(KEYINPUT39), .B(KEYINPUT105), .ZN(n485) );
  NAND2_X1 U538 ( .A1(n477), .A2(n574), .ZN(n478) );
  NOR2_X1 U539 ( .A1(n578), .A2(n478), .ZN(n480) );
  XNOR2_X1 U540 ( .A(KEYINPUT37), .B(KEYINPUT104), .ZN(n479) );
  XNOR2_X1 U541 ( .A(n480), .B(n479), .ZN(n508) );
  NOR2_X1 U542 ( .A1(n508), .A2(n481), .ZN(n482) );
  XOR2_X1 U543 ( .A(KEYINPUT38), .B(n482), .Z(n493) );
  NOR2_X1 U544 ( .A1(n483), .A2(n493), .ZN(n484) );
  XNOR2_X1 U545 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U546 ( .A(G29GAT), .B(n486), .Z(G1328GAT) );
  NOR2_X1 U547 ( .A1(n487), .A2(n493), .ZN(n488) );
  XOR2_X1 U548 ( .A(G36GAT), .B(n488), .Z(G1329GAT) );
  XOR2_X1 U549 ( .A(KEYINPUT107), .B(KEYINPUT106), .Z(n490) );
  XNOR2_X1 U550 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n490), .B(n489), .ZN(n492) );
  NOR2_X1 U552 ( .A1(n548), .A2(n493), .ZN(n491) );
  XOR2_X1 U553 ( .A(n492), .B(n491), .Z(G1330GAT) );
  NOR2_X1 U554 ( .A1(n494), .A2(n493), .ZN(n495) );
  XOR2_X1 U555 ( .A(G50GAT), .B(n495), .Z(G1331GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n499) );
  INV_X1 U557 ( .A(n549), .ZN(n569) );
  NAND2_X1 U558 ( .A1(n554), .A2(n569), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n496), .B(KEYINPUT108), .ZN(n507) );
  NOR2_X1 U560 ( .A1(n507), .A2(n497), .ZN(n504) );
  NAND2_X1 U561 ( .A1(n504), .A2(n520), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U563 ( .A(G57GAT), .B(n500), .ZN(G1332GAT) );
  NAND2_X1 U564 ( .A1(n511), .A2(n504), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n501), .B(KEYINPUT110), .ZN(n502) );
  XNOR2_X1 U566 ( .A(G64GAT), .B(n502), .ZN(G1333GAT) );
  NAND2_X1 U567 ( .A1(n562), .A2(n504), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n503), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U569 ( .A(G78GAT), .B(KEYINPUT43), .Z(n506) );
  NAND2_X1 U570 ( .A1(n504), .A2(n524), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n506), .B(n505), .ZN(G1335GAT) );
  NOR2_X1 U572 ( .A1(n508), .A2(n507), .ZN(n509) );
  XOR2_X1 U573 ( .A(KEYINPUT111), .B(n509), .Z(n514) );
  NAND2_X1 U574 ( .A1(n520), .A2(n514), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n510), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U576 ( .A1(n514), .A2(n511), .ZN(n512) );
  XNOR2_X1 U577 ( .A(G92GAT), .B(n512), .ZN(G1337GAT) );
  NAND2_X1 U578 ( .A1(n562), .A2(n514), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n513), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT44), .B(KEYINPUT112), .Z(n516) );
  NAND2_X1 U581 ( .A1(n514), .A2(n524), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U583 ( .A(G106GAT), .B(n517), .Z(G1339GAT) );
  NOR2_X1 U584 ( .A1(n519), .A2(n518), .ZN(n521) );
  NAND2_X1 U585 ( .A1(n521), .A2(n520), .ZN(n535) );
  NOR2_X1 U586 ( .A1(n548), .A2(n535), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n522), .B(KEYINPUT113), .ZN(n523) );
  NOR2_X1 U588 ( .A1(n524), .A2(n523), .ZN(n532) );
  NAND2_X1 U589 ( .A1(n532), .A2(n549), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n525), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n527) );
  NAND2_X1 U592 ( .A1(n532), .A2(n554), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U594 ( .A(G120GAT), .B(n528), .ZN(G1341GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n530) );
  NAND2_X1 U596 ( .A1(n532), .A2(n557), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U598 ( .A(G127GAT), .B(n531), .ZN(G1342GAT) );
  XOR2_X1 U599 ( .A(G134GAT), .B(KEYINPUT51), .Z(n534) );
  NAND2_X1 U600 ( .A1(n532), .A2(n561), .ZN(n533) );
  XNOR2_X1 U601 ( .A(n534), .B(n533), .ZN(G1343GAT) );
  NOR2_X1 U602 ( .A1(n536), .A2(n535), .ZN(n543) );
  NAND2_X1 U603 ( .A1(n549), .A2(n543), .ZN(n537) );
  XNOR2_X1 U604 ( .A(G141GAT), .B(n537), .ZN(G1344GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n539) );
  NAND2_X1 U606 ( .A1(n543), .A2(n554), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U608 ( .A(G148GAT), .B(n540), .ZN(G1345GAT) );
  NAND2_X1 U609 ( .A1(n543), .A2(n557), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n541), .B(KEYINPUT116), .ZN(n542) );
  XNOR2_X1 U611 ( .A(G155GAT), .B(n542), .ZN(G1346GAT) );
  NAND2_X1 U612 ( .A1(n561), .A2(n543), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n544), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U614 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n547), .B(KEYINPUT55), .ZN(n564) );
  NOR2_X1 U616 ( .A1(n548), .A2(n564), .ZN(n558) );
  NAND2_X1 U617 ( .A1(n558), .A2(n549), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n550), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT57), .B(KEYINPUT118), .Z(n552) );
  XNOR2_X1 U620 ( .A(G176GAT), .B(KEYINPUT117), .ZN(n551) );
  XNOR2_X1 U621 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U622 ( .A(KEYINPUT56), .B(n553), .Z(n556) );
  NAND2_X1 U623 ( .A1(n558), .A2(n554), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(G1349GAT) );
  XOR2_X1 U625 ( .A(G183GAT), .B(KEYINPUT119), .Z(n560) );
  NAND2_X1 U626 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1350GAT) );
  XNOR2_X1 U628 ( .A(G190GAT), .B(KEYINPUT120), .ZN(n568) );
  XOR2_X1 U629 ( .A(KEYINPUT121), .B(KEYINPUT58), .Z(n566) );
  NAND2_X1 U630 ( .A1(n562), .A2(n561), .ZN(n563) );
  OR2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(G1351GAT) );
  NOR2_X1 U634 ( .A1(n569), .A2(n579), .ZN(n573) );
  XOR2_X1 U635 ( .A(KEYINPUT59), .B(KEYINPUT123), .Z(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  NOR2_X1 U639 ( .A1(n579), .A2(n574), .ZN(n575) );
  XOR2_X1 U640 ( .A(G211GAT), .B(n575), .Z(G1354GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT125), .B(KEYINPUT62), .Z(n577) );
  XNOR2_X1 U642 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n581) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U645 ( .A(n581), .B(n580), .Z(G1355GAT) );
endmodule

