//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1287, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n206), .A2(new_n207), .ZN(new_n218));
  NAND4_X1  g0018(.A1(new_n218), .A2(G1), .A3(G13), .A4(G20), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G107), .ZN(new_n223));
  INV_X1    g0023(.A(G264), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n214), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n217), .B(new_n219), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  NAND2_X1  g0040(.A1(new_n207), .A2(G68), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n202), .A2(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT65), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G97), .B(G107), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  XNOR2_X1  g0050(.A(KEYINPUT3), .B(G33), .ZN(new_n251));
  INV_X1    g0051(.A(G1698), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n251), .A2(G222), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(G223), .A3(G1698), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n253), .B(new_n254), .C1(new_n221), .C2(new_n251), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G1), .A2(G13), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n256), .B1(G33), .B2(G41), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT66), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT66), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G41), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n211), .B(G274), .C1(new_n263), .C2(G45), .ZN(new_n264));
  INV_X1    g0064(.A(G226), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G41), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(G1), .A3(G13), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n264), .B1(new_n265), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n258), .A2(new_n271), .A3(G190), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n270), .B1(new_n257), .B2(new_n255), .ZN(new_n273));
  INV_X1    g0073(.A(G200), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n256), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n211), .A2(G20), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G50), .ZN(new_n283));
  OAI22_X1  g0083(.A1(new_n281), .A2(new_n283), .B1(G50), .B2(new_n276), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n208), .A2(G20), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT68), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT68), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n208), .A2(new_n287), .A3(G20), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n212), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT67), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n290), .B(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT8), .B(G58), .ZN(new_n293));
  INV_X1    g0093(.A(G150), .ZN(new_n294));
  NOR2_X1   g0094(.A1(G20), .A2(G33), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  OAI22_X1  g0096(.A1(new_n292), .A2(new_n293), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n289), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n284), .B1(new_n299), .B2(new_n279), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n275), .B1(new_n300), .B2(KEYINPUT9), .ZN(new_n301));
  INV_X1    g0101(.A(new_n284), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n297), .B1(new_n286), .B2(new_n288), .ZN(new_n303));
  INV_X1    g0103(.A(new_n279), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT9), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n305), .A2(KEYINPUT71), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT71), .B1(new_n305), .B2(new_n306), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n301), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT10), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT10), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n301), .B(new_n312), .C1(new_n308), .C2(new_n309), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G179), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n273), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n316), .B1(G169), .B2(new_n273), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n317), .A2(new_n300), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G274), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT66), .B(G41), .ZN(new_n321));
  INV_X1    g0121(.A(G45), .ZN(new_n322));
  AOI211_X1 g0122(.A(G1), .B(new_n320), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n269), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n323), .B1(G244), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n251), .A2(G238), .A3(G1698), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(new_n223), .B2(new_n251), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT3), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G33), .ZN(new_n329));
  INV_X1    g0129(.A(G33), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT3), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n332), .A2(new_n233), .A3(G1698), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n257), .B1(new_n327), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(G169), .B1(new_n325), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT70), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n325), .A2(new_n334), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n335), .A2(new_n336), .B1(new_n337), .B2(G179), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n325), .A2(new_n334), .A3(KEYINPUT70), .A4(new_n315), .ZN(new_n339));
  OAI22_X1  g0139(.A1(new_n293), .A2(new_n296), .B1(new_n212), .B2(new_n221), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT15), .B(G87), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n341), .A2(new_n290), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n279), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT69), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n276), .B(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n304), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n282), .A2(G77), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n343), .B1(G77), .B2(new_n345), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n339), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n348), .B1(G200), .B2(new_n337), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n325), .A2(new_n334), .A3(G190), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n338), .A2(new_n349), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n314), .A2(new_n319), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT72), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT72), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n314), .A2(new_n355), .A3(new_n319), .A4(new_n352), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g0157(.A(new_n290), .B(KEYINPUT67), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G77), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n295), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n304), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT11), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT12), .ZN(new_n363));
  INV_X1    g0163(.A(new_n345), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n363), .B1(new_n364), .B2(new_n202), .ZN(new_n365));
  INV_X1    g0165(.A(G13), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n366), .A2(G1), .ZN(new_n367));
  AND4_X1   g0167(.A1(new_n363), .A2(new_n367), .A3(G20), .A4(new_n202), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n362), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n282), .A2(G68), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n361), .A2(KEYINPUT11), .B1(new_n346), .B2(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n324), .A2(G238), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n373), .A2(new_n264), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n251), .A2(G232), .A3(G1698), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n251), .A2(G226), .A3(new_n252), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G33), .A2(G97), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n257), .ZN(new_n379));
  XNOR2_X1  g0179(.A(KEYINPUT73), .B(KEYINPUT13), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n374), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n374), .A2(new_n379), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT13), .ZN(new_n384));
  OAI211_X1 g0184(.A(G190), .B(new_n381), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  AND3_X1   g0185(.A1(new_n374), .A2(new_n379), .A3(new_n380), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n380), .B1(new_n374), .B2(new_n379), .ZN(new_n387));
  OAI21_X1  g0187(.A(G200), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n372), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n372), .ZN(new_n391));
  OAI21_X1  g0191(.A(G169), .B1(new_n386), .B2(new_n387), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT14), .ZN(new_n393));
  INV_X1    g0193(.A(new_n380), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n382), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n381), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT14), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n396), .A2(new_n397), .A3(G169), .ZN(new_n398));
  OAI211_X1 g0198(.A(G179), .B(new_n381), .C1(new_n383), .C2(new_n384), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n393), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n390), .B1(new_n391), .B2(new_n400), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n203), .B(new_n205), .C1(new_n201), .C2(new_n202), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n402), .A2(G20), .B1(G159), .B2(new_n295), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT7), .ZN(new_n404));
  AND2_X1   g0204(.A1(KEYINPUT74), .A2(G33), .ZN(new_n405));
  NOR2_X1   g0205(.A1(KEYINPUT74), .A2(G33), .ZN(new_n406));
  NOR3_X1   g0206(.A1(new_n405), .A2(new_n406), .A3(new_n328), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT75), .B1(new_n330), .B2(KEYINPUT3), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT75), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n409), .A2(new_n328), .A3(G33), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n404), .B(new_n212), .C1(new_n407), .C2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(G68), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT74), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n330), .ZN(new_n415));
  NAND2_X1  g0215(.A1(KEYINPUT74), .A2(G33), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n415), .A2(KEYINPUT3), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(new_n408), .A3(new_n410), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n404), .B1(new_n418), .B2(new_n212), .ZN(new_n419));
  OAI211_X1 g0219(.A(KEYINPUT16), .B(new_n403), .C1(new_n413), .C2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT16), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n404), .A2(G20), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT3), .B1(new_n415), .B2(new_n416), .ZN(new_n423));
  INV_X1    g0223(.A(new_n331), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n404), .B1(new_n251), .B2(G20), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n202), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n403), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n421), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n420), .A2(new_n429), .A3(new_n279), .ZN(new_n430));
  INV_X1    g0230(.A(new_n293), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n282), .ZN(new_n432));
  OAI22_X1  g0232(.A1(new_n281), .A2(new_n432), .B1(new_n276), .B2(new_n431), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n264), .B1(new_n233), .B2(new_n269), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n407), .A2(new_n411), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n437), .A2(KEYINPUT76), .A3(G223), .A4(new_n252), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n265), .A2(new_n252), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n417), .A2(new_n408), .A3(new_n410), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(G33), .A2(G87), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT76), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n417), .A2(new_n252), .A3(new_n408), .A4(new_n410), .ZN(new_n444));
  INV_X1    g0244(.A(G223), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n438), .A2(new_n442), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n436), .B1(new_n447), .B2(new_n257), .ZN(new_n448));
  INV_X1    g0248(.A(G169), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI211_X1 g0250(.A(new_n315), .B(new_n436), .C1(new_n447), .C2(new_n257), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n435), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT18), .ZN(new_n453));
  INV_X1    g0253(.A(new_n422), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n328), .B1(new_n405), .B2(new_n406), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n454), .B1(new_n455), .B2(new_n331), .ZN(new_n456));
  AOI21_X1  g0256(.A(KEYINPUT7), .B1(new_n332), .B2(new_n212), .ZN(new_n457));
  OAI21_X1  g0257(.A(G68), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n403), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n304), .B1(new_n459), .B2(new_n421), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n433), .B1(new_n460), .B2(new_n420), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n447), .A2(new_n257), .ZN(new_n462));
  INV_X1    g0262(.A(new_n436), .ZN(new_n463));
  AOI21_X1  g0263(.A(G200), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AOI211_X1 g0264(.A(G190), .B(new_n436), .C1(new_n447), .C2(new_n257), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT17), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n462), .A2(G179), .A3(new_n463), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(new_n449), .B2(new_n448), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT18), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n470), .A2(new_n471), .A3(new_n435), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n461), .B(KEYINPUT17), .C1(new_n464), .C2(new_n465), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n453), .A2(new_n468), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  XOR2_X1   g0274(.A(new_n474), .B(KEYINPUT77), .Z(new_n475));
  AND3_X1   g0275(.A1(new_n357), .A2(new_n401), .A3(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT83), .ZN(new_n477));
  INV_X1    g0277(.A(G116), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n478), .B1(new_n211), .B2(G33), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT69), .B1(new_n367), .B2(G20), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n276), .A2(new_n344), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n304), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(G116), .B2(new_n345), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G283), .ZN(new_n484));
  INV_X1    g0284(.A(G97), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n484), .B(new_n212), .C1(G33), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n478), .A2(G20), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n279), .A2(KEYINPUT82), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT82), .B1(new_n279), .B2(new_n487), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT20), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(KEYINPUT20), .B(new_n486), .C1(new_n488), .C2(new_n489), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n483), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n408), .A2(new_n410), .ZN(new_n495));
  NOR2_X1   g0295(.A1(G257), .A2(G1698), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n496), .B1(new_n224), .B2(G1698), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n417), .A3(new_n497), .ZN(new_n498));
  XNOR2_X1  g0298(.A(KEYINPUT81), .B(G303), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n332), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n267), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n263), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n211), .B(G45), .C1(new_n502), .C2(G41), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n503), .A2(new_n505), .A3(G274), .A4(new_n267), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT5), .B1(new_n260), .B2(new_n262), .ZN(new_n507));
  OAI211_X1 g0307(.A(G270), .B(new_n267), .C1(new_n507), .C2(new_n504), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(G169), .B1(new_n501), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n477), .B1(new_n494), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT21), .ZN(new_n512));
  INV_X1    g0312(.A(new_n494), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n501), .A2(new_n509), .A3(new_n315), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT21), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n477), .B(new_n516), .C1(new_n494), .C2(new_n510), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n501), .A2(new_n509), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G190), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n519), .B(new_n494), .C1(new_n274), .C2(new_n518), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n512), .A2(new_n515), .A3(new_n517), .A4(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(G250), .A2(G1698), .ZN(new_n522));
  INV_X1    g0322(.A(G257), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n522), .B1(new_n523), .B2(G1698), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n524), .A2(new_n417), .A3(new_n408), .A4(new_n410), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n415), .A2(new_n416), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G294), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n257), .ZN(new_n529));
  INV_X1    g0329(.A(G190), .ZN(new_n530));
  OAI211_X1 g0330(.A(G264), .B(new_n267), .C1(new_n507), .C2(new_n504), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n529), .A2(new_n530), .A3(new_n506), .A4(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n267), .B1(new_n525), .B2(new_n527), .ZN(new_n533));
  INV_X1    g0333(.A(new_n531), .ZN(new_n534));
  NOR4_X1   g0334(.A1(new_n507), .A2(new_n257), .A3(new_n504), .A4(new_n320), .ZN(new_n535));
  NOR3_X1   g0335(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n532), .B1(new_n536), .B2(G200), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT22), .ZN(new_n538));
  INV_X1    g0338(.A(G87), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(G20), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n538), .B1(new_n332), .B2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n212), .B(G116), .C1(new_n405), .C2(new_n406), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT84), .ZN(new_n544));
  OAI22_X1  g0344(.A1(new_n544), .A2(KEYINPUT23), .B1(new_n212), .B2(G107), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n212), .A2(G107), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n544), .A2(KEYINPUT23), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT23), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n548), .A2(KEYINPUT84), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n546), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n542), .A2(new_n543), .A3(new_n545), .A4(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n417), .A2(new_n212), .A3(new_n408), .A4(new_n410), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n538), .A2(new_n539), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NOR3_X1   g0355(.A1(new_n551), .A2(new_n555), .A3(KEYINPUT24), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT24), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n550), .A2(new_n543), .A3(new_n545), .ZN(new_n558));
  AOI21_X1  g0358(.A(KEYINPUT22), .B1(new_n251), .B2(new_n540), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n437), .A2(new_n212), .A3(new_n553), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n557), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n279), .B1(new_n556), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n277), .A2(new_n223), .ZN(new_n564));
  XNOR2_X1  g0364(.A(new_n564), .B(KEYINPUT25), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n211), .A2(G33), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n276), .A2(new_n566), .A3(new_n256), .A4(new_n278), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n567), .A2(new_n223), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n537), .A2(new_n563), .A3(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n495), .A2(G244), .A3(new_n252), .A4(new_n417), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT4), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n251), .A2(KEYINPUT4), .A3(G244), .A4(new_n252), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n251), .A2(G250), .A3(G1698), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n574), .A2(new_n484), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n267), .B1(new_n573), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n267), .B1(new_n507), .B2(new_n504), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n506), .B1(new_n523), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n449), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n579), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n574), .A2(new_n484), .A3(new_n575), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(new_n572), .B2(new_n571), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n581), .B(new_n315), .C1(new_n583), .C2(new_n267), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n223), .B1(new_n425), .B2(new_n426), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT6), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n586), .A2(new_n485), .A3(G107), .ZN(new_n587));
  XNOR2_X1  g0387(.A(G97), .B(G107), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n587), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  OAI22_X1  g0389(.A1(new_n589), .A2(new_n212), .B1(new_n221), .B2(new_n296), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n279), .B1(new_n585), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n567), .A2(G97), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(G97), .B2(new_n277), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT78), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n592), .B(KEYINPUT78), .C1(G97), .C2(new_n277), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n591), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n580), .A2(new_n584), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(G200), .B1(new_n577), .B2(new_n579), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n581), .B(G190), .C1(new_n583), .C2(new_n267), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n588), .A2(new_n586), .ZN(new_n602));
  INV_X1    g0402(.A(new_n587), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n604), .A2(G20), .B1(G77), .B2(new_n295), .ZN(new_n605));
  OAI21_X1  g0405(.A(G107), .B1(new_n456), .B2(new_n457), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n607), .A2(new_n279), .B1(new_n595), .B2(new_n596), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n600), .A2(new_n601), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n570), .A2(new_n599), .A3(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(G238), .A2(G1698), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n611), .B1(new_n222), .B2(G1698), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n495), .A2(new_n417), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n526), .A2(G116), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n267), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(G250), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(new_n322), .B2(G1), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n211), .A2(new_n320), .A3(G45), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n267), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g0419(.A(new_n619), .B(KEYINPUT79), .ZN(new_n620));
  OAI21_X1  g0420(.A(G200), .B1(new_n615), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT79), .ZN(new_n622));
  XNOR2_X1  g0422(.A(new_n619), .B(new_n622), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n437), .A2(new_n612), .B1(G116), .B2(new_n526), .ZN(new_n624));
  OAI211_X1 g0424(.A(G190), .B(new_n623), .C1(new_n624), .C2(new_n267), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n495), .A2(new_n212), .A3(G68), .A4(new_n417), .ZN(new_n626));
  OR2_X1    g0426(.A1(KEYINPUT80), .A2(G87), .ZN(new_n627));
  NOR2_X1   g0427(.A1(G97), .A2(G107), .ZN(new_n628));
  NAND2_X1  g0428(.A1(KEYINPUT80), .A2(G87), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT19), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n377), .B2(new_n212), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n212), .A2(G33), .A3(G97), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n630), .A2(new_n632), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n304), .B1(new_n626), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n341), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n345), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n567), .A2(new_n539), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n621), .A2(new_n625), .A3(new_n638), .A4(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n634), .B1(new_n552), .B2(new_n202), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n279), .ZN(new_n643));
  INV_X1    g0443(.A(new_n637), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n567), .A2(new_n341), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n449), .B1(new_n615), .B2(new_n620), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n315), .B(new_n623), .C1(new_n624), .C2(new_n267), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n569), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT24), .B1(new_n551), .B2(new_n555), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n560), .A2(new_n557), .A3(new_n561), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n650), .B1(new_n653), .B2(new_n279), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n529), .A2(new_n315), .A3(new_n506), .A4(new_n531), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n536), .B2(G169), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n641), .B(new_n649), .C1(new_n654), .C2(new_n656), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n521), .A2(new_n610), .A3(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n476), .A2(new_n658), .ZN(G372));
  AND3_X1   g0459(.A1(new_n580), .A2(new_n598), .A3(new_n584), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n625), .A2(new_n621), .ZN(new_n661));
  AOI21_X1  g0461(.A(KEYINPUT85), .B1(new_n638), .B2(new_n640), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT85), .ZN(new_n663));
  NOR4_X1   g0463(.A1(new_n635), .A2(new_n637), .A3(new_n663), .A4(new_n639), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n661), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n660), .A2(new_n665), .A3(new_n666), .A4(new_n649), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n641), .A2(new_n649), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT26), .B1(new_n668), .B2(new_n599), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n667), .A2(new_n649), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n563), .A2(new_n569), .ZN(new_n671));
  INV_X1    g0471(.A(new_n536), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n449), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n671), .A2(new_n655), .A3(new_n673), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n674), .A2(new_n517), .A3(new_n515), .A4(new_n512), .ZN(new_n675));
  INV_X1    g0475(.A(new_n610), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n665), .A2(new_n649), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n670), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n476), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n468), .A2(new_n389), .A3(new_n473), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n338), .A2(new_n349), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n399), .B1(new_n392), .B2(KEYINPUT14), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n397), .B1(new_n396), .B2(G169), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n391), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n681), .B1(new_n682), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n453), .A2(new_n472), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n314), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n319), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n680), .A2(new_n690), .ZN(G369));
  AND2_X1   g0491(.A1(new_n512), .A2(new_n515), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n517), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n367), .A2(new_n212), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G213), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G343), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n494), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n693), .A2(new_n701), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n521), .A2(new_n701), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT86), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT86), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n702), .A2(new_n706), .A3(new_n703), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n674), .A2(new_n699), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n671), .A2(new_n699), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n570), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n708), .B1(new_n674), .B2(new_n710), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n705), .A2(G330), .A3(new_n707), .A4(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n699), .B1(new_n692), .B2(new_n517), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n710), .A2(new_n674), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n708), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n712), .A2(new_n715), .ZN(G399));
  INV_X1    g0516(.A(new_n215), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(new_n263), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n218), .ZN(new_n719));
  INV_X1    g0519(.A(new_n718), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G1), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n630), .A2(G116), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT28), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n660), .A2(new_n665), .A3(KEYINPUT26), .A4(new_n649), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT89), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n727), .B(new_n666), .C1(new_n668), .C2(new_n599), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n573), .A2(new_n576), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n579), .B1(new_n730), .B2(new_n257), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n731), .A2(new_n315), .B1(new_n591), .B2(new_n597), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n732), .A2(new_n580), .A3(new_n641), .A4(new_n649), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n727), .B1(new_n733), .B2(new_n666), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n649), .B1(new_n729), .B2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT90), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n725), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI211_X1 g0537(.A(KEYINPUT90), .B(new_n649), .C1(new_n729), .C2(new_n734), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n699), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT29), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(G330), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n610), .A2(new_n657), .ZN(new_n743));
  INV_X1    g0543(.A(new_n521), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n743), .A2(new_n744), .A3(new_n700), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT88), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n658), .A2(KEYINPUT88), .A3(new_n700), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT87), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT30), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n533), .A2(new_n534), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n615), .A2(new_n620), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n514), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n731), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n750), .B(new_n751), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  NOR3_X1   g0556(.A1(new_n518), .A2(new_n753), .A3(G179), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(new_n755), .A3(new_n672), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n753), .A2(new_n752), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n750), .A2(new_n751), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n759), .A2(new_n514), .A3(new_n731), .A4(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n756), .A2(new_n758), .A3(new_n761), .ZN(new_n762));
  AND3_X1   g0562(.A1(new_n762), .A2(KEYINPUT31), .A3(new_n699), .ZN(new_n763));
  AOI21_X1  g0563(.A(KEYINPUT31), .B1(new_n762), .B2(new_n699), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n742), .B1(new_n749), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n699), .B1(new_n670), .B2(new_n678), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n767), .A2(new_n740), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n741), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n724), .B1(new_n769), .B2(G1), .ZN(G364));
  NOR2_X1   g0570(.A1(new_n366), .A2(G20), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n211), .B1(new_n771), .B2(G45), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n718), .A2(new_n773), .ZN(new_n774));
  XOR2_X1   g0574(.A(new_n774), .B(KEYINPUT91), .Z(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n212), .B1(KEYINPUT93), .B2(new_n449), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n449), .A2(KEYINPUT93), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n256), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n530), .A2(G179), .A3(G200), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n212), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n485), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n212), .A2(new_n315), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G190), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G200), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT32), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n212), .A2(G179), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G190), .A2(G200), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(KEYINPUT94), .B(G159), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n787), .A2(new_n201), .B1(new_n788), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n785), .A2(new_n274), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n783), .B(new_n794), .C1(G50), .C2(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n789), .A2(G190), .A3(G200), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(new_n627), .B2(new_n629), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n274), .A2(G190), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n789), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n223), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n798), .A2(new_n332), .A3(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT95), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n784), .A2(new_n799), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n784), .A2(new_n790), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n202), .A2(new_n804), .B1(new_n805), .B2(new_n221), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(new_n788), .B2(new_n793), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n796), .A2(new_n803), .A3(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n797), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n809), .A2(G303), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n251), .B(new_n810), .C1(G326), .C2(new_n795), .ZN(new_n811));
  INV_X1    g0611(.A(new_n800), .ZN(new_n812));
  INV_X1    g0612(.A(new_n791), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n812), .A2(G283), .B1(new_n813), .B2(G329), .ZN(new_n814));
  INV_X1    g0614(.A(new_n804), .ZN(new_n815));
  XNOR2_X1  g0615(.A(KEYINPUT33), .B(G317), .ZN(new_n816));
  INV_X1    g0616(.A(new_n805), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n815), .A2(new_n816), .B1(new_n817), .B2(G311), .ZN(new_n818));
  INV_X1    g0618(.A(new_n782), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G294), .A2(new_n819), .B1(new_n786), .B2(G322), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n811), .A2(new_n814), .A3(new_n818), .A4(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n780), .B1(new_n808), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(G13), .A2(G33), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(G20), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n779), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n717), .A2(new_n332), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n827), .A2(G355), .B1(new_n478), .B2(new_n717), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n418), .A2(new_n215), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT92), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n218), .A2(new_n322), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n245), .B2(new_n322), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n828), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n776), .B(new_n822), .C1(new_n826), .C2(new_n834), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n705), .A2(new_n707), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n825), .B(KEYINPUT96), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n836), .A2(G330), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n718), .B2(new_n773), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n836), .A2(G330), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n838), .B1(new_n840), .B2(new_n841), .ZN(G396));
  INV_X1    g0642(.A(KEYINPUT99), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n682), .B2(new_n700), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n338), .A2(new_n349), .A3(KEYINPUT99), .A4(new_n699), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n348), .A2(new_n699), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT98), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n846), .B(new_n847), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n844), .A2(new_n845), .B1(new_n352), .B2(new_n848), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n699), .B(new_n849), .C1(new_n678), .C2(new_n670), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n849), .B(KEYINPUT100), .Z(new_n852));
  OAI21_X1  g0652(.A(new_n851), .B1(new_n767), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n766), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n774), .B1(new_n853), .B2(new_n854), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n849), .A2(new_n823), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n780), .A2(new_n824), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT97), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n775), .B1(new_n860), .B2(G77), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n786), .A2(G143), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n862), .B1(new_n294), .B2(new_n804), .C1(new_n792), .C2(new_n805), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(G137), .B2(new_n795), .ZN(new_n864));
  OR2_X1    g0664(.A1(new_n864), .A2(KEYINPUT34), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(KEYINPUT34), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n812), .A2(G68), .ZN(new_n867));
  INV_X1    g0667(.A(G132), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n867), .B1(new_n207), .B2(new_n797), .C1(new_n868), .C2(new_n791), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n418), .B(new_n869), .C1(G58), .C2(new_n819), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n865), .A2(new_n866), .A3(new_n870), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n251), .B(new_n783), .C1(G107), .C2(new_n809), .ZN(new_n872));
  AOI22_X1  g0672(.A1(G283), .A2(new_n815), .B1(new_n813), .B2(G311), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n800), .A2(new_n539), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(G116), .B2(new_n817), .ZN(new_n875));
  AOI22_X1  g0675(.A1(G294), .A2(new_n786), .B1(new_n795), .B2(G303), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n872), .A2(new_n873), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n871), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n861), .B1(new_n878), .B2(new_n779), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n856), .A2(new_n857), .B1(new_n858), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(G384));
  NOR3_X1   g0681(.A1(new_n256), .A2(new_n212), .A3(new_n478), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n589), .B(KEYINPUT101), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT35), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n886), .B1(new_n885), .B2(new_n884), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(KEYINPUT36), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n218), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n889));
  AOI211_X1 g0689(.A(new_n211), .B(G13), .C1(new_n889), .C2(new_n241), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n476), .B1(new_n741), .B2(new_n768), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n690), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n682), .A2(new_n699), .ZN(new_n894));
  INV_X1    g0694(.A(new_n849), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n894), .B1(new_n767), .B2(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n391), .B(new_n699), .C1(new_n390), .C2(new_n400), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n391), .A2(new_n699), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n685), .A2(new_n389), .A3(new_n898), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  XOR2_X1   g0701(.A(KEYINPUT103), .B(KEYINPUT37), .Z(new_n902));
  INV_X1    g0702(.A(new_n697), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n435), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n452), .A2(new_n466), .A3(new_n902), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n448), .A2(new_n530), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n440), .A2(new_n441), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n495), .A2(G223), .A3(new_n252), .A4(new_n417), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n907), .B1(new_n443), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n267), .B1(new_n909), .B2(new_n438), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n274), .B1(new_n910), .B2(new_n436), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n435), .B1(new_n906), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n403), .B1(new_n413), .B2(new_n419), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n304), .B1(new_n913), .B2(new_n421), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT102), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n420), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI211_X1 g0716(.A(KEYINPUT102), .B(new_n304), .C1(new_n913), .C2(new_n421), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n434), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n469), .B(new_n697), .C1(new_n449), .C2(new_n448), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n912), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT37), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n905), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n918), .A2(new_n903), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n474), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT38), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n922), .A2(new_n924), .A3(KEYINPUT38), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n901), .A2(new_n929), .B1(new_n687), .B2(new_n697), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT39), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n922), .A2(new_n924), .A3(KEYINPUT38), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT104), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n905), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n435), .B1(new_n470), .B2(new_n903), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n935), .A2(KEYINPUT104), .A3(new_n466), .A4(new_n902), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n452), .A2(new_n466), .A3(new_n904), .ZN(new_n937));
  INV_X1    g0737(.A(new_n902), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n934), .A2(new_n936), .A3(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n904), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n474), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT38), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n931), .B1(new_n932), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n927), .A2(KEYINPUT39), .A3(new_n928), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n400), .A2(new_n391), .A3(new_n700), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n944), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n930), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n893), .B(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(KEYINPUT88), .B1(new_n658), .B2(new_n700), .ZN(new_n951));
  AND4_X1   g0751(.A1(KEYINPUT88), .A2(new_n743), .A3(new_n744), .A4(new_n700), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n765), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n476), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n932), .A2(new_n943), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n897), .A2(new_n899), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n895), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n953), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(KEYINPUT40), .B1(new_n955), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT40), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n957), .B1(new_n749), .B2(new_n765), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n929), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n742), .B1(new_n954), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n954), .B2(new_n964), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n950), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n211), .B2(new_n771), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n950), .A2(new_n966), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n891), .B1(new_n968), .B2(new_n969), .ZN(G367));
  AND2_X1   g0770(.A1(new_n609), .A2(new_n599), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n598), .A2(new_n699), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(KEYINPUT105), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n660), .A2(new_n699), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT105), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n971), .A2(new_n976), .A3(new_n972), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n974), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT106), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n599), .B1(new_n980), .B2(new_n674), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n700), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n978), .A2(new_n711), .A3(new_n713), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT42), .Z(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  OR3_X1    g0785(.A1(new_n662), .A2(new_n664), .A3(new_n700), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n677), .A2(new_n986), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n986), .A2(new_n649), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT43), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n989), .A2(KEYINPUT43), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n985), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n980), .A2(new_n712), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n982), .A2(new_n991), .A3(new_n990), .A4(new_n984), .ZN(new_n996));
  AND3_X1   g0796(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n995), .B1(new_n994), .B2(new_n996), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n718), .B(KEYINPUT41), .Z(new_n1000));
  INV_X1    g0800(.A(KEYINPUT108), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n769), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n711), .A2(new_n713), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n711), .A2(new_n713), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n839), .B(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1001), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n839), .B(new_n1005), .Z(new_n1008));
  NAND3_X1  g0808(.A1(new_n1008), .A2(KEYINPUT108), .A3(new_n769), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n978), .A2(new_n715), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT45), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT44), .ZN(new_n1013));
  OR3_X1    g0813(.A1(new_n978), .A2(new_n715), .A3(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1013), .B1(new_n978), .B2(new_n715), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1012), .A2(new_n1016), .A3(new_n712), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT107), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n712), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1020), .A2(new_n1018), .A3(new_n1017), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1007), .A2(new_n1009), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1000), .B1(new_n1024), .B2(new_n769), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n999), .B1(new_n1025), .B2(new_n773), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n826), .B1(new_n215), .B2(new_n341), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n830), .B2(new_n239), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n809), .A2(G58), .B1(new_n813), .B2(G137), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n207), .B2(new_n805), .C1(new_n792), .C2(new_n804), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n782), .A2(new_n202), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n332), .B(new_n1031), .C1(G77), .C2(new_n812), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(G143), .A2(new_n795), .B1(new_n786), .B2(G150), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n809), .A2(G116), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT46), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G283), .A2(new_n817), .B1(new_n815), .B2(G294), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n800), .A2(new_n485), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(G317), .B2(new_n813), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1036), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n437), .B1(new_n499), .B2(new_n786), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G107), .A2(new_n819), .B1(new_n795), .B2(G311), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n1030), .A2(new_n1034), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT47), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n776), .B(new_n1028), .C1(new_n1045), .C2(new_n779), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n989), .B2(new_n837), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1026), .A2(new_n1047), .ZN(G387));
  NOR2_X1   g0848(.A1(new_n1006), .A2(new_n772), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT109), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n819), .A2(G283), .B1(new_n809), .B2(G294), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n499), .A2(new_n817), .B1(new_n815), .B2(G311), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n786), .A2(G317), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n795), .A2(G322), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT48), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1051), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT111), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1058), .A2(KEYINPUT49), .A3(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n812), .A2(G116), .B1(new_n813), .B2(G326), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1060), .A2(new_n418), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(KEYINPUT49), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n782), .A2(new_n341), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G159), .B2(new_n795), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n207), .B2(new_n787), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1038), .B(new_n418), .C1(G77), .C2(new_n809), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n817), .A2(G68), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n431), .A2(new_n815), .B1(new_n813), .B2(G150), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n1062), .A2(new_n1063), .B1(new_n1066), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT112), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n780), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n1072), .B2(new_n1071), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n831), .B1(G45), .B2(new_n236), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n722), .B2(new_n827), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n293), .A2(G50), .ZN(new_n1077));
  XOR2_X1   g0877(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n1078));
  XNOR2_X1  g0878(.A(new_n1077), .B(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n322), .B1(new_n202), .B2(new_n221), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n1079), .A2(new_n722), .A3(new_n1080), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n1076), .A2(new_n1081), .B1(G107), .B2(new_n215), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n776), .B1(new_n1082), .B2(new_n826), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1074), .B(new_n1083), .C1(new_n711), .C2(new_n837), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n718), .B1(new_n1008), .B2(new_n769), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1050), .B(new_n1084), .C1(new_n1085), .C2(new_n1086), .ZN(G393));
  AND2_X1   g0887(.A1(new_n1021), .A2(new_n1017), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n718), .B(new_n1024), .C1(new_n1085), .C2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n874), .B1(G143), .B2(new_n813), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n202), .B2(new_n797), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n418), .B(new_n1091), .C1(G77), .C2(new_n819), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G150), .A2(new_n795), .B1(new_n786), .B2(G159), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT51), .Z(new_n1094));
  OAI22_X1  g0894(.A1(new_n207), .A2(new_n804), .B1(new_n805), .B2(new_n293), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT113), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1092), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G311), .A2(new_n786), .B1(new_n795), .B2(G317), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT52), .Z(new_n1099));
  AOI22_X1  g0899(.A1(new_n499), .A2(new_n815), .B1(new_n817), .B2(G294), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n809), .A2(G283), .B1(new_n813), .B2(G322), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n251), .B(new_n801), .C1(G116), .C2(new_n819), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n780), .B1(new_n1097), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n830), .A2(new_n249), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1105), .B(new_n826), .C1(new_n485), .C2(new_n215), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n775), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1104), .B(new_n1107), .C1(new_n980), .C2(new_n825), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(new_n1088), .B2(new_n773), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1089), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT114), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1089), .A2(KEYINPUT114), .A3(new_n1109), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(G390));
  INV_X1    g0914(.A(new_n943), .ZN(new_n1115));
  AOI21_X1  g0915(.A(KEYINPUT39), .B1(new_n1115), .B2(new_n928), .ZN(new_n1116));
  AOI21_X1  g0916(.A(KEYINPUT38), .B1(new_n922), .B2(new_n924), .ZN(new_n1117));
  NOR3_X1   g0917(.A1(new_n932), .A2(new_n1117), .A3(new_n931), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n823), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n775), .B1(new_n860), .B2(new_n431), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n797), .A2(new_n294), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1121), .B(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT54), .B(G143), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(G137), .A2(new_n815), .B1(new_n817), .B2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1123), .B(new_n1126), .C1(new_n207), .C2(new_n800), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(G159), .A2(new_n819), .B1(new_n795), .B2(G128), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n332), .B1(new_n813), .B2(G125), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1128), .B(new_n1129), .C1(new_n868), .C2(new_n787), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(G107), .A2(new_n815), .B1(new_n813), .B2(G294), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1131), .B1(new_n539), .B2(new_n797), .C1(new_n485), .C2(new_n805), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(G116), .A2(new_n786), .B1(new_n795), .B2(G283), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n819), .A2(G77), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1133), .A2(new_n332), .A3(new_n867), .A4(new_n1134), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n1127), .A2(new_n1130), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1120), .B1(new_n1136), .B2(new_n779), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1119), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n946), .B1(new_n932), .B2(new_n943), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n894), .B1(new_n739), .B2(new_n895), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1140), .B1(new_n1141), .B2(new_n900), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n1116), .A2(new_n1118), .B1(new_n901), .B2(new_n947), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n953), .A2(new_n958), .A3(G330), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n735), .A2(new_n736), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1146), .A2(new_n678), .A3(new_n738), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1147), .A2(new_n700), .A3(new_n895), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n894), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1139), .B1(new_n1150), .B2(new_n956), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n956), .B1(new_n850), .B2(new_n894), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n944), .A2(new_n945), .B1(new_n1152), .B2(new_n946), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT115), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1144), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n766), .A2(KEYINPUT115), .A3(new_n958), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1145), .B1(new_n1154), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1138), .B1(new_n1159), .B2(new_n772), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT116), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n476), .A2(new_n766), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n892), .A2(new_n690), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n766), .A2(new_n852), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n900), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1166), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n766), .A2(new_n895), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1156), .A2(new_n1157), .B1(new_n1168), .B2(new_n900), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1167), .B1(new_n1169), .B2(new_n896), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1162), .B1(new_n1164), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n1159), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n718), .B1(new_n1171), .B2(new_n1159), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1161), .B1(new_n1173), .B2(new_n1174), .ZN(G378));
  OAI21_X1  g0975(.A(new_n774), .B1(new_n860), .B2(G50), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n300), .A2(new_n697), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n314), .B2(new_n319), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n318), .B(new_n1179), .C1(new_n311), .C2(new_n313), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1178), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n309), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n307), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n312), .B1(new_n1185), .B2(new_n301), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n313), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n319), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n1179), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n314), .A2(new_n319), .A3(new_n1180), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1189), .A2(new_n1190), .A3(new_n1177), .ZN(new_n1191));
  AND2_X1   g0991(.A1(new_n1183), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1193), .A2(new_n824), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n330), .B(new_n259), .C1(new_n800), .C2(new_n792), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(G150), .A2(new_n819), .B1(new_n795), .B2(G125), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT119), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(G132), .A2(new_n815), .B1(new_n817), .B2(G137), .ZN(new_n1198));
  INV_X1    g0998(.A(G128), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1198), .B1(new_n797), .B2(new_n1124), .C1(new_n1199), .C2(new_n787), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT120), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n1202), .A2(KEYINPUT59), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1195), .B(new_n1203), .C1(G124), .C2(new_n813), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(KEYINPUT59), .B2(new_n1202), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n804), .A2(new_n485), .B1(new_n800), .B2(new_n201), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n418), .A2(new_n321), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(new_n636), .C2(new_n817), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n786), .A2(G107), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT118), .ZN(new_n1210));
  INV_X1    g1010(.A(G283), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n797), .A2(new_n221), .B1(new_n791), .B2(new_n1211), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1031), .B(new_n1212), .C1(G116), .C2(new_n795), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1208), .A2(new_n1210), .A3(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT58), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1207), .B(new_n207), .C1(G33), .C2(G41), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1205), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1176), .B(new_n1194), .C1(new_n779), .C2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1193), .B1(new_n964), .B2(G330), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n742), .B(new_n1192), .C1(new_n960), .C2(new_n963), .ZN(new_n1222));
  OAI21_X1  g1022(.A(KEYINPUT121), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n949), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n953), .B(new_n958), .C1(new_n932), .C2(new_n943), .ZN(new_n1226));
  AOI21_X1  g1026(.A(KEYINPUT40), .B1(new_n927), .B2(new_n928), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(KEYINPUT40), .A2(new_n1226), .B1(new_n1227), .B2(new_n962), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1192), .B1(new_n1228), .B2(new_n742), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n964), .A2(G330), .A3(new_n1193), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1231), .A2(KEYINPUT121), .A3(new_n949), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1225), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1220), .B1(new_n1233), .B2(new_n773), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1168), .A2(new_n900), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1158), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n896), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1144), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n900), .B2(new_n1165), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n1236), .A2(new_n1237), .B1(new_n1239), .B2(new_n1141), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1164), .B1(new_n1159), .B2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(KEYINPUT57), .B1(new_n1233), .B2(new_n1241), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1229), .A2(new_n1230), .A3(new_n1224), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1224), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1244));
  OAI21_X1  g1044(.A(KEYINPUT57), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n892), .A2(new_n690), .A3(new_n1163), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(new_n1151), .A2(new_n1153), .A3(new_n1238), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1158), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1246), .B1(new_n1249), .B2(new_n1170), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n718), .B1(new_n1245), .B2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1234), .B1(new_n1242), .B2(new_n1251), .ZN(G375));
  NAND2_X1  g1052(.A1(new_n1240), .A2(new_n1246), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1000), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1164), .A2(new_n1170), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n900), .A2(new_n823), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n775), .B1(new_n860), .B2(G68), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1064), .B1(G294), .B2(new_n795), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(G107), .A2(new_n817), .B1(new_n815), .B2(G116), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n809), .A2(G97), .B1(new_n813), .B2(G303), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n786), .A2(G283), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .A4(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n332), .B1(new_n800), .B2(new_n221), .ZN(new_n1264));
  XOR2_X1   g1064(.A(new_n1264), .B(KEYINPUT122), .Z(new_n1265));
  AOI22_X1  g1065(.A1(G132), .A2(new_n795), .B1(new_n786), .B2(G137), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1266), .B1(new_n207), .B2(new_n782), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(G150), .A2(new_n817), .B1(new_n812), .B2(G58), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n809), .A2(G159), .B1(new_n813), .B2(G128), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n815), .A2(new_n1125), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1268), .A2(new_n1269), .A3(new_n437), .A4(new_n1270), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n1263), .A2(new_n1265), .B1(new_n1267), .B2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1258), .B1(new_n1272), .B2(new_n779), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1170), .A2(new_n773), .B1(new_n1257), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1256), .A2(new_n1274), .ZN(G381));
  INV_X1    g1075(.A(new_n1113), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT114), .B1(new_n1089), .B2(new_n1109), .ZN(new_n1277));
  NOR3_X1   g1077(.A1(G387), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(G393), .A2(G396), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NOR3_X1   g1080(.A1(new_n1280), .A2(G384), .A3(G381), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1255), .A2(KEYINPUT116), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n720), .B1(new_n1282), .B2(new_n1249), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1160), .B1(new_n1283), .B2(new_n1172), .ZN(new_n1284));
  INV_X1    g1084(.A(G375), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1278), .A2(new_n1281), .A3(new_n1284), .A4(new_n1285), .ZN(G407));
  NAND3_X1  g1086(.A1(new_n1285), .A2(new_n698), .A3(new_n1284), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(G407), .A2(new_n1287), .A3(G213), .ZN(G409));
  INV_X1    g1088(.A(KEYINPUT124), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(G393), .A2(G396), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1291), .A2(new_n1279), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(new_n1112), .A2(new_n1113), .B1(new_n1026), .B2(new_n1047), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1289), .B(new_n1292), .C1(new_n1278), .C2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1280), .A2(new_n1289), .A3(new_n1290), .ZN(new_n1295));
  OAI21_X1  g1095(.A(G387), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1296));
  OAI21_X1  g1096(.A(KEYINPUT124), .B1(new_n1291), .B2(new_n1279), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1112), .A2(new_n1026), .A3(new_n1047), .A4(new_n1113), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1295), .A2(new_n1296), .A3(new_n1297), .A4(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1294), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT61), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1240), .A2(KEYINPUT60), .A3(new_n1246), .ZN(new_n1302));
  AND2_X1   g1102(.A1(new_n1302), .A2(new_n718), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1255), .A2(KEYINPUT60), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1253), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(G384), .B1(new_n1306), .B2(new_n1274), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1274), .ZN(new_n1309));
  AOI211_X1 g1109(.A(new_n880), .B(new_n1309), .C1(new_n1303), .C2(new_n1305), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n698), .A2(G213), .A3(G2897), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1308), .A2(new_n1311), .A3(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1312), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1314), .B1(new_n1307), .B2(new_n1310), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1313), .A2(new_n1315), .ZN(new_n1316));
  OAI211_X1 g1116(.A(G378), .B(new_n1234), .C1(new_n1242), .C2(new_n1251), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n949), .B1(new_n1231), .B2(KEYINPUT121), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1241), .B(new_n1254), .C1(new_n1318), .C2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1231), .A2(new_n949), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1229), .A2(new_n1230), .A3(new_n1224), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1220), .B1(new_n1323), .B2(new_n773), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1320), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n1284), .ZN(new_n1326));
  AOI22_X1  g1126(.A1(new_n1317), .A2(new_n1326), .B1(G213), .B2(new_n698), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1301), .B1(new_n1316), .B2(new_n1327), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1300), .A2(new_n1328), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1307), .A2(new_n1310), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1327), .A2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT63), .ZN(new_n1332));
  OAI21_X1  g1132(.A(KEYINPUT125), .B1(new_n1331), .B2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT125), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1327), .A2(new_n1334), .A3(KEYINPUT63), .A4(new_n1330), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1333), .A2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1331), .A2(KEYINPUT123), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT123), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1327), .A2(new_n1338), .A3(new_n1330), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1337), .A2(new_n1332), .A3(new_n1339), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1329), .A2(new_n1336), .A3(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1317), .A2(new_n1326), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n698), .A2(G213), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1342), .A2(KEYINPUT62), .A3(new_n1343), .A4(new_n1330), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT126), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  NAND4_X1  g1146(.A1(new_n1327), .A2(KEYINPUT126), .A3(KEYINPUT62), .A4(new_n1330), .ZN(new_n1347));
  AND2_X1   g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT62), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1337), .A2(new_n1349), .A3(new_n1339), .ZN(new_n1350));
  AOI21_X1  g1150(.A(new_n1328), .B1(new_n1348), .B2(new_n1350), .ZN(new_n1351));
  AND2_X1   g1151(.A1(new_n1294), .A2(new_n1299), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1341), .B1(new_n1351), .B2(new_n1352), .ZN(G405));
  NAND2_X1  g1153(.A1(G375), .A2(new_n1284), .ZN(new_n1354));
  AOI21_X1  g1154(.A(KEYINPUT127), .B1(new_n1354), .B2(new_n1317), .ZN(new_n1355));
  INV_X1    g1155(.A(new_n1355), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1354), .A2(KEYINPUT127), .A3(new_n1317), .ZN(new_n1357));
  OAI211_X1 g1157(.A(new_n1356), .B(new_n1357), .C1(new_n1307), .C2(new_n1310), .ZN(new_n1358));
  INV_X1    g1158(.A(new_n1357), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1330), .B1(new_n1359), .B2(new_n1355), .ZN(new_n1360));
  AND3_X1   g1160(.A1(new_n1352), .A2(new_n1358), .A3(new_n1360), .ZN(new_n1361));
  AOI21_X1  g1161(.A(new_n1352), .B1(new_n1360), .B2(new_n1358), .ZN(new_n1362));
  NOR2_X1   g1162(.A1(new_n1361), .A2(new_n1362), .ZN(G402));
endmodule


