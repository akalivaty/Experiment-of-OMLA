//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 1 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 1 0 1 0 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n772,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  OAI21_X1  g001(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT90), .ZN(new_n204));
  OR2_X1    g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n204), .ZN(new_n206));
  NOR2_X1   g005(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n207));
  INV_X1    g006(.A(G36gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AND3_X1   g008(.A1(new_n205), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT91), .B(G29gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(new_n208), .ZN(new_n212));
  OAI211_X1 g011(.A(KEYINPUT15), .B(new_n202), .C1(new_n210), .C2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT15), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n202), .B(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n209), .A2(KEYINPUT92), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT92), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n207), .A2(new_n217), .A3(new_n208), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n218), .A3(new_n203), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n212), .A2(KEYINPUT93), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT93), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(new_n211), .B2(new_n208), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n215), .A2(new_n219), .A3(new_n220), .A4(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n213), .A2(new_n223), .A3(KEYINPUT17), .ZN(new_n224));
  XNOR2_X1  g023(.A(G15gat), .B(G22gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT16), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n225), .B1(new_n226), .B2(G1gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(G1gat), .B2(new_n225), .ZN(new_n228));
  INV_X1    g027(.A(G8gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n228), .B(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n224), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT17), .B1(new_n213), .B2(new_n223), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n213), .A2(new_n223), .ZN(new_n234));
  INV_X1    g033(.A(new_n230), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G229gat), .A2(G233gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT18), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n236), .A2(KEYINPUT18), .A3(new_n237), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n230), .B(new_n234), .Z(new_n242));
  XOR2_X1   g041(.A(new_n237), .B(KEYINPUT13), .Z(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n240), .A2(new_n241), .A3(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G169gat), .B(G197gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(KEYINPUT89), .ZN(new_n247));
  INV_X1    g046(.A(G113gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n250));
  INV_X1    g049(.A(G141gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n249), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT12), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n245), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n240), .A2(new_n241), .A3(new_n244), .A4(new_n254), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AND2_X1   g057(.A1(G71gat), .A2(G78gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(G71gat), .A2(G78gat), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n259), .B1(KEYINPUT9), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(G57gat), .ZN(new_n262));
  INV_X1    g061(.A(G64gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G57gat), .A2(G64gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT95), .B1(new_n261), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT95), .ZN(new_n268));
  AND2_X1   g067(.A1(G57gat), .A2(G64gat), .ZN(new_n269));
  NOR2_X1   g068(.A1(G57gat), .A2(G64gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n260), .A2(KEYINPUT9), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n268), .B(new_n271), .C1(new_n272), .C2(new_n259), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT94), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n274), .B1(new_n269), .B2(new_n270), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n264), .A2(KEYINPUT94), .A3(new_n265), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(new_n276), .A3(KEYINPUT9), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n259), .A2(new_n260), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n267), .A2(new_n273), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n279), .A2(KEYINPUT21), .ZN(new_n280));
  NAND2_X1  g079(.A1(G231gat), .A2(G233gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G127gat), .B(G155gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT20), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n282), .B(new_n284), .ZN(new_n285));
  XOR2_X1   g084(.A(G183gat), .B(G211gat), .Z(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n235), .B1(KEYINPUT21), .B2(new_n279), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  OR2_X1    g089(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n287), .A2(new_n290), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  OR2_X1    g093(.A1(G99gat), .A2(G106gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(G99gat), .A2(G106gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(KEYINPUT97), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT97), .ZN(new_n298));
  AND2_X1   g097(.A1(G99gat), .A2(G106gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(G99gat), .A2(G106gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G85gat), .A2(G92gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT7), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT7), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(G85gat), .A3(G92gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G85gat), .ZN(new_n308));
  INV_X1    g107(.A(G92gat), .ZN(new_n309));
  AOI22_X1  g108(.A1(KEYINPUT8), .A2(new_n296), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n302), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n301), .A2(new_n297), .A3(new_n307), .A4(new_n310), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AND2_X1   g113(.A1(G232gat), .A2(G233gat), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n234), .A2(new_n314), .B1(KEYINPUT41), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n314), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n224), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n316), .B1(new_n318), .B2(new_n232), .ZN(new_n319));
  XNOR2_X1  g118(.A(G190gat), .B(G218gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n319), .B(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n315), .A2(KEYINPUT41), .ZN(new_n322));
  XNOR2_X1  g121(.A(G134gat), .B(G162gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n322), .B(new_n323), .ZN(new_n324));
  OR2_X1    g123(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n321), .A2(new_n324), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(G230gat), .A2(G233gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n267), .A2(new_n273), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n297), .A2(new_n301), .A3(KEYINPUT98), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n331), .A2(new_n307), .A3(new_n310), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n311), .A2(KEYINPUT98), .A3(new_n301), .A4(new_n297), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n277), .A2(new_n278), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n330), .A2(new_n332), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n335), .B(KEYINPUT99), .C1(new_n279), .C2(new_n314), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT99), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n279), .A2(new_n337), .A3(new_n333), .A4(new_n332), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT10), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n279), .A2(KEYINPUT10), .A3(new_n314), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n329), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n335), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT99), .B1(new_n279), .B2(new_n314), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n338), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n342), .B1(new_n329), .B2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G120gat), .B(G148gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(G176gat), .B(G204gat), .ZN(new_n348));
  XOR2_X1   g147(.A(new_n347), .B(new_n348), .Z(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  OR2_X1    g149(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n346), .A2(new_n350), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NOR3_X1   g153(.A1(new_n294), .A2(new_n328), .A3(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G197gat), .B(G204gat), .ZN(new_n356));
  INV_X1    g155(.A(G211gat), .ZN(new_n357));
  INV_X1    g156(.A(G218gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n356), .B1(KEYINPUT22), .B2(new_n359), .ZN(new_n360));
  XOR2_X1   g159(.A(G211gat), .B(G218gat), .Z(new_n361));
  XOR2_X1   g160(.A(new_n360), .B(new_n361), .Z(new_n362));
  AND3_X1   g161(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(G190gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT66), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT66), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(G190gat), .ZN(new_n369));
  INV_X1    g168(.A(G183gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n367), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(G169gat), .A2(G176gat), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT65), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(KEYINPUT23), .A3(new_n376), .ZN(new_n377));
  AND2_X1   g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n373), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT23), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n372), .A2(new_n377), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT25), .B1(G169gat), .B2(G176gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n373), .A2(KEYINPUT23), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n383), .B1(new_n384), .B2(KEYINPUT64), .ZN(new_n385));
  NOR2_X1   g184(.A1(G183gat), .A2(G190gat), .ZN(new_n386));
  NOR3_X1   g185(.A1(new_n363), .A2(new_n364), .A3(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n373), .A2(KEYINPUT23), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n384), .B1(new_n389), .B2(KEYINPUT64), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n382), .A2(KEYINPUT25), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n370), .A2(KEYINPUT27), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT27), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(G183gat), .ZN(new_n394));
  AND3_X1   g193(.A1(new_n392), .A2(new_n394), .A3(KEYINPUT68), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT68), .B1(new_n392), .B2(new_n394), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n367), .A2(new_n369), .A3(KEYINPUT28), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n367), .A2(new_n369), .A3(new_n392), .A4(new_n394), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT28), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT67), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n399), .A2(KEYINPUT67), .A3(new_n400), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n398), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n378), .B1(new_n379), .B2(KEYINPUT26), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n375), .A2(new_n376), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n406), .B1(new_n407), .B2(KEYINPUT26), .ZN(new_n408));
  NAND2_X1  g207(.A1(G183gat), .A2(G190gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n391), .B1(new_n405), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(G226gat), .A2(G233gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT75), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n411), .A2(KEYINPUT75), .A3(new_n413), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT66), .B(G190gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT27), .B(G183gat), .ZN(new_n419));
  AOI211_X1 g218(.A(new_n402), .B(KEYINPUT28), .C1(new_n418), .C2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT67), .B1(new_n399), .B2(new_n400), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n392), .A2(new_n394), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT68), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n419), .A2(KEYINPUT68), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI22_X1  g225(.A1(new_n420), .A2(new_n421), .B1(new_n426), .B2(new_n397), .ZN(new_n427));
  INV_X1    g226(.A(new_n410), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n427), .A2(KEYINPUT69), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT69), .B1(new_n427), .B2(new_n428), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n391), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT29), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n413), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n362), .B1(new_n417), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n431), .A2(new_n413), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n411), .A2(new_n432), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT76), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(new_n437), .A3(new_n412), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n427), .A2(new_n428), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT29), .B1(new_n439), .B2(new_n391), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT76), .B1(new_n440), .B2(new_n413), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n360), .B(new_n361), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n435), .A2(new_n438), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(G8gat), .B(G36gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(G64gat), .B(G92gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(KEYINPUT78), .B(KEYINPUT79), .ZN(new_n447));
  XOR2_X1   g246(.A(new_n446), .B(new_n447), .Z(new_n448));
  NAND3_X1  g247(.A1(new_n434), .A2(new_n443), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT30), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n443), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n382), .A2(KEYINPUT25), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n388), .A2(new_n390), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT69), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n456), .B1(new_n405), .B2(new_n410), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n427), .A2(new_n428), .A3(KEYINPUT69), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n455), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n412), .B1(new_n459), .B2(KEYINPUT29), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT75), .ZN(new_n461));
  AOI211_X1 g260(.A(new_n461), .B(new_n412), .C1(new_n439), .C2(new_n391), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n462), .A2(new_n414), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n442), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT77), .B1(new_n452), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT77), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n434), .A2(new_n466), .A3(new_n443), .ZN(new_n467));
  INV_X1    g266(.A(new_n448), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n449), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n451), .B1(new_n470), .B2(KEYINPUT30), .ZN(new_n471));
  XNOR2_X1  g270(.A(G113gat), .B(G120gat), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n472), .A2(KEYINPUT1), .ZN(new_n473));
  XNOR2_X1  g272(.A(G127gat), .B(G134gat), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n472), .A2(KEYINPUT70), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT1), .ZN(new_n477));
  INV_X1    g276(.A(G120gat), .ZN(new_n478));
  OR3_X1    g277(.A1(new_n478), .A2(KEYINPUT70), .A3(G113gat), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n476), .A2(new_n477), .A3(new_n474), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT71), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT71), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n475), .A2(new_n483), .A3(new_n480), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n431), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n485), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n459), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(G227gat), .A2(G233gat), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n486), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT34), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT34), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n486), .A2(new_n488), .A3(new_n492), .A4(new_n489), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT73), .ZN(new_n495));
  XNOR2_X1  g294(.A(G15gat), .B(G43gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n496), .B(KEYINPUT72), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(G71gat), .ZN(new_n498));
  INV_X1    g297(.A(G99gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n498), .B(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n489), .B1(new_n486), .B2(new_n488), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n500), .B1(new_n501), .B2(KEYINPUT33), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT32), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n486), .A2(new_n488), .ZN(new_n506));
  INV_X1    g305(.A(new_n489), .ZN(new_n507));
  AOI221_X4 g306(.A(new_n503), .B1(KEYINPUT33), .B2(new_n500), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n495), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n431), .A2(new_n485), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n459), .A2(new_n487), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT32), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT33), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n515), .A3(new_n500), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n502), .A2(new_n504), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT73), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n518), .B1(new_n491), .B2(new_n493), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(KEYINPUT84), .B(G22gat), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G78gat), .B(G106gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(G155gat), .A2(G162gat), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT2), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(G155gat), .A2(G162gat), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n251), .A2(G148gat), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n526), .A2(new_n527), .B1(new_n528), .B2(KEYINPUT80), .ZN(new_n529));
  XNOR2_X1  g328(.A(G141gat), .B(G148gat), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT80), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT81), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n529), .A2(KEYINPUT81), .A3(new_n532), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT3), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n530), .A2(KEYINPUT2), .ZN(new_n539));
  INV_X1    g338(.A(new_n524), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n527), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n537), .A2(new_n538), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n442), .B1(new_n544), .B2(new_n432), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n542), .B1(new_n535), .B2(new_n536), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n442), .A2(new_n432), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n546), .B1(new_n547), .B2(new_n538), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n523), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  AOI211_X1 g348(.A(KEYINPUT3), .B(new_n542), .C1(new_n535), .C2(new_n536), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n362), .B1(new_n550), .B2(KEYINPUT29), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n547), .A2(new_n538), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n543), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n523), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n551), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT31), .B(G50gat), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n549), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n557), .B1(new_n549), .B2(new_n556), .ZN(new_n560));
  INV_X1    g359(.A(G228gat), .ZN(new_n561));
  INV_X1    g360(.A(G233gat), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NOR3_X1   g362(.A1(new_n559), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n563), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n556), .ZN(new_n566));
  INV_X1    g365(.A(new_n557), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n565), .B1(new_n568), .B2(new_n558), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n522), .B1(new_n564), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n563), .B1(new_n559), .B2(new_n560), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n568), .A2(new_n565), .A3(new_n558), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n571), .A2(new_n521), .A3(new_n572), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n509), .A2(new_n520), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G1gat), .B(G29gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT0), .ZN(new_n576));
  XNOR2_X1  g375(.A(G57gat), .B(G85gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  NAND2_X1  g377(.A1(G225gat), .A2(G233gat), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n481), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n546), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n546), .A2(new_n581), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n580), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n482), .A2(new_n546), .A3(KEYINPUT4), .A4(new_n484), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n586), .B(new_n579), .C1(new_n583), .C2(KEYINPUT4), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n481), .B1(new_n546), .B2(new_n538), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n588), .A2(new_n550), .ZN(new_n589));
  OAI211_X1 g388(.A(KEYINPUT5), .B(new_n585), .C1(new_n587), .C2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT4), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n482), .A2(new_n546), .A3(new_n591), .A4(new_n484), .ZN(new_n592));
  OAI211_X1 g391(.A(KEYINPUT82), .B(new_n592), .C1(new_n583), .C2(new_n591), .ZN(new_n593));
  INV_X1    g392(.A(new_n589), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT82), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n582), .A2(new_n595), .A3(KEYINPUT4), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n580), .A2(KEYINPUT5), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n593), .A2(new_n594), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n578), .B1(new_n590), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n590), .A2(new_n598), .A3(new_n578), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT6), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n599), .B1(new_n602), .B2(KEYINPUT83), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT83), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n600), .A2(new_n604), .A3(new_n601), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n599), .A2(KEYINPUT6), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n471), .A2(new_n574), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT35), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n491), .B(new_n493), .C1(new_n505), .C2(new_n508), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n516), .A2(new_n517), .A3(new_n494), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n570), .A2(new_n573), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n590), .A2(new_n598), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n578), .B(KEYINPUT85), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n617), .A2(new_n601), .A3(new_n600), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT35), .B1(new_n618), .B2(new_n607), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n471), .A2(new_n613), .A3(new_n614), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n610), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT87), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n623));
  NOR3_X1   g422(.A1(new_n583), .A2(new_n580), .A3(new_n584), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n593), .A2(new_n594), .A3(new_n596), .ZN(new_n625));
  AOI211_X1 g424(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n580), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n625), .A2(new_n623), .A3(new_n580), .ZN(new_n627));
  INV_X1    g426(.A(new_n616), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT40), .ZN(new_n630));
  OR3_X1    g429(.A1(new_n626), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n630), .B1(new_n626), .B2(new_n629), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n631), .A2(new_n617), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n614), .B1(new_n471), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n465), .A2(KEYINPUT37), .A3(new_n467), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n468), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(KEYINPUT86), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT86), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n635), .A2(new_n638), .A3(new_n468), .ZN(new_n639));
  OR3_X1    g438(.A1(new_n452), .A2(new_n464), .A3(KEYINPUT37), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n637), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT38), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n442), .B1(new_n417), .B2(new_n433), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n435), .A2(new_n438), .A3(new_n441), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n643), .B(KEYINPUT37), .C1(new_n644), .C2(new_n442), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n448), .A2(KEYINPUT38), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n640), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n647), .A2(new_n607), .A3(new_n618), .A4(new_n449), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n634), .B1(new_n642), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT36), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n509), .A2(new_n520), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n612), .A2(KEYINPUT74), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(KEYINPUT74), .A2(KEYINPUT36), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n611), .A2(new_n612), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n607), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n658), .B1(new_n603), .B2(new_n605), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n450), .B1(new_n469), .B2(new_n449), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n659), .A2(new_n660), .A3(new_n451), .ZN(new_n661));
  OAI22_X1  g460(.A1(new_n654), .A2(new_n657), .B1(new_n661), .B2(new_n614), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n621), .B(new_n622), .C1(new_n650), .C2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n614), .ZN(new_n665));
  INV_X1    g464(.A(new_n471), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n665), .B1(new_n666), .B2(new_n659), .ZN(new_n667));
  INV_X1    g466(.A(new_n653), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n509), .A2(new_n520), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT36), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(new_n656), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n648), .B1(new_n641), .B2(KEYINPUT38), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n667), .B(new_n671), .C1(new_n672), .C2(new_n634), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n622), .B1(new_n673), .B2(new_n621), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n258), .B(new_n355), .C1(new_n664), .C2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT100), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n673), .A2(new_n621), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(KEYINPUT87), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(new_n663), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n680), .A2(KEYINPUT100), .A3(new_n258), .A4(new_n355), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n659), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g483(.A(new_n229), .B1(new_n682), .B2(new_n666), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT101), .B(KEYINPUT16), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(G8gat), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  AOI211_X1 g487(.A(new_n471), .B(new_n688), .C1(new_n677), .C2(new_n681), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT42), .B1(new_n685), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n682), .A2(new_n666), .A3(new_n687), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT42), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n690), .A2(new_n693), .ZN(G1325gat));
  AOI21_X1  g493(.A(new_n671), .B1(new_n677), .B2(new_n681), .ZN(new_n695));
  INV_X1    g494(.A(G15gat), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n613), .ZN(new_n698));
  AOI211_X1 g497(.A(G15gat), .B(new_n698), .C1(new_n677), .C2(new_n681), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT102), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n682), .A2(new_n696), .A3(new_n613), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT102), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n701), .B(new_n702), .C1(new_n696), .C2(new_n695), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n700), .A2(new_n703), .ZN(G1326gat));
  NAND2_X1  g503(.A1(new_n682), .A2(new_n665), .ZN(new_n705));
  XNOR2_X1  g504(.A(KEYINPUT43), .B(G22gat), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1327gat));
  NOR3_X1   g506(.A1(new_n293), .A2(new_n327), .A3(new_n354), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n258), .B(new_n708), .C1(new_n664), .C2(new_n674), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n659), .A2(new_n211), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT45), .Z(new_n712));
  AOI21_X1  g511(.A(new_n327), .B1(new_n673), .B2(new_n621), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(KEYINPUT44), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n327), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n714), .B1(new_n680), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n293), .B(KEYINPUT103), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n258), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n720), .A2(new_n721), .A3(new_n354), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n718), .A2(new_n608), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n712), .B1(new_n211), .B2(new_n724), .ZN(G1328gat));
  NAND2_X1  g524(.A1(new_n666), .A2(new_n208), .ZN(new_n726));
  OAI21_X1  g525(.A(KEYINPUT46), .B1(new_n709), .B2(new_n726), .ZN(new_n727));
  OR3_X1    g526(.A1(new_n709), .A2(KEYINPUT46), .A3(new_n726), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n718), .A2(new_n471), .A3(new_n723), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n727), .B(new_n728), .C1(new_n729), .C2(new_n208), .ZN(G1329gat));
  INV_X1    g529(.A(G43gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(new_n709), .B2(new_n698), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT104), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n716), .B1(new_n664), .B2(new_n674), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n678), .A2(new_n328), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n715), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n671), .A2(new_n731), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n734), .A2(new_n736), .A3(new_n722), .A4(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n732), .A2(new_n733), .A3(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT105), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT47), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n739), .A2(new_n740), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n732), .A2(KEYINPUT105), .A3(new_n738), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n744), .A2(KEYINPUT47), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n742), .B1(new_n743), .B2(new_n745), .ZN(G1330gat));
  NAND4_X1  g545(.A1(new_n717), .A2(G50gat), .A3(new_n665), .A4(new_n722), .ZN(new_n747));
  INV_X1    g546(.A(G50gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n709), .B2(new_n614), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT106), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT48), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n747), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n750), .A2(KEYINPUT48), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1331gat));
  NAND3_X1  g553(.A1(new_n721), .A2(new_n293), .A3(new_n327), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(new_n353), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT107), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n678), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n659), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G57gat), .ZN(G1332gat));
  INV_X1    g559(.A(KEYINPUT49), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n666), .B1(new_n761), .B2(new_n263), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT108), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n758), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n761), .A2(new_n263), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(G1333gat));
  INV_X1    g565(.A(new_n671), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n758), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n698), .A2(G71gat), .ZN(new_n769));
  AOI22_X1  g568(.A1(new_n768), .A2(G71gat), .B1(new_n758), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g570(.A1(new_n758), .A2(new_n665), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G78gat), .ZN(G1335gat));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n293), .A2(new_n258), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n678), .A2(new_n328), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n774), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n713), .A2(KEYINPUT109), .A3(KEYINPUT51), .A4(new_n775), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n776), .A2(new_n777), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT110), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT110), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n608), .A2(G85gat), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n783), .A2(new_n354), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n293), .A2(new_n258), .A3(new_n353), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n717), .A2(new_n659), .A3(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n787), .B1(new_n308), .B2(new_n789), .ZN(G1336gat));
  NAND3_X1  g589(.A1(new_n717), .A2(new_n666), .A3(new_n788), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G92gat), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n471), .A2(G92gat), .A3(new_n353), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n792), .B(new_n793), .C1(new_n782), .C2(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n776), .B(KEYINPUT51), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(new_n795), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n798), .B1(G92gat), .B2(new_n791), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n796), .B1(new_n793), .B2(new_n799), .ZN(G1337gat));
  NAND3_X1  g599(.A1(new_n717), .A2(new_n767), .A3(new_n788), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT111), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n499), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n803), .B1(new_n802), .B2(new_n801), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n698), .A2(G99gat), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n783), .A2(new_n354), .A3(new_n785), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(G1338gat));
  NAND4_X1  g606(.A1(new_n734), .A2(new_n736), .A3(new_n665), .A4(new_n788), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(G106gat), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n614), .A2(G106gat), .A3(new_n353), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n809), .B1(new_n797), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT53), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n808), .A2(KEYINPUT113), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(G106gat), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n808), .A2(KEYINPUT113), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n814), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT112), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n781), .A2(new_n819), .A3(new_n810), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n781), .B2(new_n810), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n813), .B1(new_n818), .B2(new_n822), .ZN(G1339gat));
  OAI21_X1  g622(.A(new_n350), .B1(new_n342), .B2(KEYINPUT54), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT10), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n341), .B1(new_n345), .B2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n329), .ZN(new_n828));
  OAI21_X1  g627(.A(KEYINPUT54), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT114), .B1(new_n827), .B2(new_n828), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI211_X1 g630(.A(new_n329), .B(new_n341), .C1(new_n345), .C2(new_n826), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT114), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT115), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n345), .A2(new_n826), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n340), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n835), .B1(new_n837), .B2(new_n329), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n836), .A2(new_n828), .A3(new_n340), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AND4_X1   g640(.A1(KEYINPUT115), .A2(new_n838), .A3(new_n833), .A4(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n825), .B1(new_n834), .B2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g644(.A(KEYINPUT55), .B(new_n825), .C1(new_n834), .C2(new_n842), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n845), .A2(new_n258), .A3(new_n351), .A4(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n236), .A2(new_n237), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n242), .A2(new_n243), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n253), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n354), .A2(new_n257), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n328), .B1(new_n847), .B2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n853));
  OAI211_X1 g652(.A(KEYINPUT54), .B(new_n342), .C1(new_n832), .C2(KEYINPUT114), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n840), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n838), .A2(new_n833), .A3(new_n841), .A4(KEYINPUT115), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n824), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n351), .B1(new_n858), .B2(KEYINPUT55), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n328), .A2(new_n257), .A3(new_n850), .ZN(new_n860));
  AOI211_X1 g659(.A(new_n844), .B(new_n824), .C1(new_n856), .C2(new_n857), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n719), .B1(new_n852), .B2(new_n862), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n755), .A2(new_n354), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n608), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n865), .A2(new_n614), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n666), .A2(new_n698), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n868), .A2(new_n248), .A3(new_n721), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n866), .A2(new_n471), .A3(new_n669), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n870), .A2(new_n721), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n869), .B1(new_n871), .B2(new_n248), .ZN(G1340gat));
  NOR3_X1   g671(.A1(new_n868), .A2(new_n478), .A3(new_n353), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n870), .A2(new_n353), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n873), .B1(new_n874), .B2(new_n478), .ZN(G1341gat));
  OAI21_X1  g674(.A(G127gat), .B1(new_n868), .B2(new_n719), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n294), .A2(G127gat), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n870), .B2(new_n877), .ZN(G1342gat));
  OR2_X1    g677(.A1(new_n327), .A2(G134gat), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n880));
  OAI22_X1  g679(.A1(new_n870), .A2(new_n879), .B1(new_n880), .B2(KEYINPUT56), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT56), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(KEYINPUT117), .B2(new_n882), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n880), .B(KEYINPUT56), .C1(new_n870), .C2(new_n879), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n866), .A2(new_n867), .A3(new_n328), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n885), .A2(KEYINPUT116), .A3(G134gat), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT116), .B1(new_n885), .B2(G134gat), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n883), .B(new_n884), .C1(new_n886), .C2(new_n887), .ZN(G1343gat));
  NAND2_X1  g687(.A1(new_n671), .A2(new_n665), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n889), .A2(new_n666), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n865), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n251), .B1(new_n891), .B2(new_n721), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n671), .A2(new_n659), .A3(new_n471), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n614), .B1(new_n863), .B2(new_n864), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT57), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(KEYINPUT118), .B1(new_n859), .B2(new_n861), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n845), .A2(new_n898), .A3(new_n351), .A4(new_n846), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n897), .A2(new_n899), .A3(new_n258), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n328), .B1(new_n900), .B2(new_n851), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n294), .B1(new_n901), .B2(new_n862), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n614), .B1(new_n902), .B2(new_n864), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n896), .B1(new_n903), .B2(new_n895), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n258), .A2(G141gat), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n892), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(KEYINPUT119), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT58), .ZN(G1344gat));
  NAND2_X1  g707(.A1(new_n902), .A2(new_n864), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n895), .A3(new_n665), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n863), .A2(new_n864), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n895), .B1(new_n911), .B2(new_n665), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n893), .A2(new_n353), .ZN(new_n915));
  OAI21_X1  g714(.A(G148gat), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n916), .A2(KEYINPUT59), .ZN(new_n917));
  INV_X1    g716(.A(G148gat), .ZN(new_n918));
  INV_X1    g717(.A(new_n904), .ZN(new_n919));
  AOI211_X1 g718(.A(KEYINPUT59), .B(new_n918), .C1(new_n919), .C2(new_n354), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n354), .A2(new_n918), .ZN(new_n921));
  OAI22_X1  g720(.A1(new_n917), .A2(new_n920), .B1(new_n891), .B2(new_n921), .ZN(G1345gat));
  OAI21_X1  g721(.A(G155gat), .B1(new_n904), .B2(new_n719), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n294), .A2(G155gat), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n891), .B2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT120), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n925), .B(new_n926), .ZN(G1346gat));
  OAI21_X1  g726(.A(G162gat), .B1(new_n904), .B2(new_n327), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n327), .A2(G162gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n928), .B1(new_n891), .B2(new_n929), .ZN(G1347gat));
  NOR2_X1   g729(.A1(new_n471), .A2(new_n659), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT122), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n911), .A2(new_n614), .A3(new_n613), .A4(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(G169gat), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n933), .A2(new_n934), .A3(new_n721), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n911), .A2(new_n931), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n574), .ZN(new_n937));
  XOR2_X1   g736(.A(new_n937), .B(KEYINPUT121), .Z(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(new_n258), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n935), .B1(new_n939), .B2(new_n934), .ZN(G1348gat));
  INV_X1    g739(.A(G176gat), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n938), .A2(new_n941), .A3(new_n354), .ZN(new_n942));
  OAI21_X1  g741(.A(G176gat), .B1(new_n933), .B2(new_n353), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1349gat));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n945), .B1(new_n933), .B2(new_n719), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(G183gat), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n933), .A2(new_n945), .A3(new_n719), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n293), .A2(new_n424), .A3(new_n425), .ZN(new_n949));
  OAI22_X1  g748(.A1(new_n947), .A2(new_n948), .B1(new_n937), .B2(new_n949), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g750(.A1(new_n938), .A2(new_n418), .A3(new_n328), .ZN(new_n952));
  OAI21_X1  g751(.A(G190gat), .B1(new_n933), .B2(new_n327), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT61), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(G1351gat));
  INV_X1    g754(.A(new_n889), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n936), .A2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(G197gat), .B1(new_n958), .B2(new_n258), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n932), .A2(new_n671), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT125), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT124), .ZN(new_n962));
  AOI211_X1 g761(.A(new_n962), .B(new_n912), .C1(new_n903), .C2(new_n895), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT124), .B1(new_n910), .B2(new_n913), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n258), .A2(G197gat), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n959), .B1(new_n966), .B2(new_n967), .ZN(G1352gat));
  OAI21_X1  g767(.A(G204gat), .B1(new_n965), .B2(new_n353), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n957), .A2(G204gat), .A3(new_n353), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n970), .B(KEYINPUT62), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n969), .A2(new_n971), .ZN(G1353gat));
  NAND3_X1  g771(.A1(new_n958), .A2(new_n357), .A3(new_n293), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n932), .A2(new_n671), .A3(new_n293), .ZN(new_n974));
  OAI21_X1  g773(.A(G211gat), .B1(new_n914), .B2(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT63), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n975), .A2(new_n976), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n973), .B1(new_n977), .B2(new_n978), .ZN(G1354gat));
  OAI21_X1  g778(.A(new_n358), .B1(new_n957), .B2(new_n327), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT126), .ZN(new_n981));
  XNOR2_X1  g780(.A(new_n980), .B(new_n981), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n328), .A2(G218gat), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n983), .B1(new_n965), .B2(KEYINPUT127), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT127), .ZN(new_n985));
  OAI211_X1 g784(.A(new_n985), .B(new_n961), .C1(new_n963), .C2(new_n964), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n982), .B1(new_n984), .B2(new_n986), .ZN(G1355gat));
endmodule


