

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742;

  AND2_X1 U370 ( .A1(n548), .A2(n578), .ZN(n350) );
  XNOR2_X1 U371 ( .A(n536), .B(n477), .ZN(n726) );
  XNOR2_X2 U372 ( .A(n486), .B(n476), .ZN(n536) );
  OR2_X2 U373 ( .A1(n701), .A2(G902), .ZN(n439) );
  NOR2_X2 U374 ( .A1(G953), .A2(G237), .ZN(n538) );
  XNOR2_X1 U375 ( .A(G122), .B(G143), .ZN(n499) );
  XNOR2_X1 U376 ( .A(n421), .B(G472), .ZN(n667) );
  INV_X1 U377 ( .A(G953), .ZN(n720) );
  AND2_X4 U378 ( .A1(n616), .A2(n615), .ZN(n454) );
  XOR2_X2 U379 ( .A(G101), .B(G119), .Z(n357) );
  NOR2_X1 U380 ( .A1(n740), .A2(n742), .ZN(n450) );
  INV_X1 U381 ( .A(G469), .ZN(n438) );
  INV_X1 U382 ( .A(KEYINPUT35), .ZN(n349) );
  NAND2_X1 U383 ( .A1(n385), .A2(n382), .ZN(n626) );
  NOR2_X1 U384 ( .A1(n376), .A2(n737), .ZN(n404) );
  AND2_X1 U385 ( .A1(n386), .A2(n387), .ZN(n385) );
  XNOR2_X1 U386 ( .A(n350), .B(n349), .ZN(n737) );
  XNOR2_X1 U387 ( .A(n414), .B(n569), .ZN(n674) );
  NOR2_X1 U388 ( .A1(n685), .A2(n351), .ZN(n435) );
  NOR2_X1 U389 ( .A1(n681), .A2(n679), .ZN(n414) );
  XNOR2_X1 U390 ( .A(n605), .B(KEYINPUT38), .ZN(n675) );
  INV_X1 U391 ( .A(n511), .ZN(n445) );
  XNOR2_X1 U392 ( .A(n441), .B(G110), .ZN(n511) );
  INV_X1 U393 ( .A(KEYINPUT73), .ZN(n398) );
  XNOR2_X1 U394 ( .A(G125), .B(G146), .ZN(n455) );
  XNOR2_X1 U395 ( .A(G113), .B(KEYINPUT3), .ZN(n510) );
  XNOR2_X1 U396 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n464) );
  XNOR2_X1 U397 ( .A(n534), .B(n448), .ZN(n351) );
  XNOR2_X1 U398 ( .A(n534), .B(n448), .ZN(n552) );
  XNOR2_X1 U399 ( .A(n546), .B(n377), .ZN(n376) );
  NOR2_X1 U400 ( .A1(n611), .A2(n356), .ZN(n400) );
  XNOR2_X1 U401 ( .A(n527), .B(n526), .ZN(n582) );
  XNOR2_X1 U402 ( .A(n407), .B(n362), .ZN(n544) );
  NOR2_X1 U403 ( .A1(n552), .A2(n447), .ZN(n407) );
  XNOR2_X1 U404 ( .A(n446), .B(n445), .ZN(n514) );
  XNOR2_X2 U405 ( .A(n370), .B(n474), .ZN(n564) );
  XNOR2_X2 U406 ( .A(n410), .B(n395), .ZN(n411) );
  INV_X1 U407 ( .A(G134), .ZN(n475) );
  XNOR2_X1 U408 ( .A(n373), .B(n372), .ZN(n590) );
  INV_X1 U409 ( .A(KEYINPUT69), .ZN(n372) );
  NOR2_X1 U410 ( .A1(n564), .A2(n374), .ZN(n373) );
  NAND2_X1 U411 ( .A1(n664), .A2(n355), .ZN(n374) );
  NAND2_X1 U412 ( .A1(n675), .A2(n676), .ZN(n681) );
  XNOR2_X1 U413 ( .A(n667), .B(n420), .ZN(n589) );
  XNOR2_X1 U414 ( .A(KEYINPUT99), .B(KEYINPUT6), .ZN(n420) );
  NAND2_X1 U415 ( .A1(n568), .A2(n676), .ZN(n527) );
  XNOR2_X1 U416 ( .A(n541), .B(n540), .ZN(n618) );
  XNOR2_X1 U417 ( .A(n417), .B(n415), .ZN(n539) );
  INV_X1 U418 ( .A(KEYINPUT45), .ZN(n395) );
  NOR2_X2 U419 ( .A1(n544), .A2(n589), .ZN(n549) );
  INV_X1 U420 ( .A(n667), .ZN(n402) );
  NAND2_X1 U421 ( .A1(n680), .A2(KEYINPUT66), .ZN(n594) );
  XNOR2_X1 U422 ( .A(n485), .B(G116), .ZN(n512) );
  XNOR2_X1 U423 ( .A(G107), .B(G122), .ZN(n485) );
  NAND2_X1 U424 ( .A1(n564), .A2(n664), .ZN(n660) );
  XNOR2_X1 U425 ( .A(n549), .B(KEYINPUT80), .ZN(n390) );
  XNOR2_X1 U426 ( .A(G137), .B(G140), .ZN(n477) );
  INV_X1 U427 ( .A(KEYINPUT24), .ZN(n456) );
  XNOR2_X1 U428 ( .A(n492), .B(n491), .ZN(n711) );
  XOR2_X1 U429 ( .A(n504), .B(n725), .Z(n708) );
  NAND2_X1 U430 ( .A1(n425), .A2(n424), .ZN(n429) );
  XOR2_X1 U431 ( .A(KEYINPUT87), .B(n525), .Z(n676) );
  XNOR2_X1 U432 ( .A(n575), .B(KEYINPUT39), .ZN(n608) );
  INV_X1 U433 ( .A(KEYINPUT1), .ZN(n437) );
  BUF_X1 U434 ( .A(n659), .Z(n396) );
  OR2_X1 U435 ( .A1(n618), .A2(G902), .ZN(n421) );
  NOR2_X1 U436 ( .A1(n389), .A2(n388), .ZN(n387) );
  INV_X1 U437 ( .A(n663), .ZN(n388) );
  NOR2_X1 U438 ( .A1(n396), .A2(KEYINPUT81), .ZN(n389) );
  INV_X1 U439 ( .A(n711), .ZN(n394) );
  NAND2_X1 U440 ( .A1(n413), .A2(n363), .ZN(n615) );
  XNOR2_X1 U441 ( .A(n557), .B(KEYINPUT98), .ZN(n680) );
  XNOR2_X1 U442 ( .A(n419), .B(n418), .ZN(n417) );
  XNOR2_X1 U443 ( .A(KEYINPUT72), .B(KEYINPUT5), .ZN(n418) );
  XNOR2_X1 U444 ( .A(n537), .B(n416), .ZN(n415) );
  XNOR2_X1 U445 ( .A(G116), .B(G146), .ZN(n537) );
  XNOR2_X1 U446 ( .A(KEYINPUT92), .B(G137), .ZN(n416) );
  XNOR2_X1 U447 ( .A(KEYINPUT4), .B(G131), .ZN(n476) );
  XNOR2_X1 U448 ( .A(n512), .B(n487), .ZN(n406) );
  XOR2_X1 U449 ( .A(KEYINPUT93), .B(KEYINPUT11), .Z(n497) );
  INV_X1 U450 ( .A(G131), .ZN(n498) );
  XNOR2_X1 U451 ( .A(G113), .B(G104), .ZN(n494) );
  INV_X1 U452 ( .A(G104), .ZN(n441) );
  XNOR2_X1 U453 ( .A(n481), .B(G107), .ZN(n440) );
  INV_X1 U454 ( .A(G146), .ZN(n481) );
  INV_X1 U455 ( .A(G101), .ZN(n478) );
  INV_X1 U456 ( .A(n455), .ZN(n518) );
  NAND2_X1 U457 ( .A1(G237), .A2(G234), .ZN(n528) );
  OR2_X1 U458 ( .A1(G902), .A2(G237), .ZN(n524) );
  INV_X1 U459 ( .A(KEYINPUT104), .ZN(n434) );
  NOR2_X1 U460 ( .A1(n605), .A2(n428), .ZN(n427) );
  INV_X1 U461 ( .A(n676), .ZN(n428) );
  NAND2_X1 U462 ( .A1(n432), .A2(n433), .ZN(n426) );
  NAND2_X1 U463 ( .A1(n591), .A2(n434), .ZN(n433) );
  NAND2_X1 U464 ( .A1(n641), .A2(n434), .ZN(n432) );
  XNOR2_X1 U465 ( .A(n726), .B(n453), .ZN(n701) );
  XNOR2_X1 U466 ( .A(n482), .B(n480), .ZN(n453) );
  XNOR2_X1 U467 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U468 ( .A(n511), .B(n440), .ZN(n482) );
  NAND2_X1 U469 ( .A1(n375), .A2(n567), .ZN(n583) );
  XNOR2_X1 U470 ( .A(n565), .B(KEYINPUT28), .ZN(n375) );
  NOR2_X1 U471 ( .A1(n641), .A2(n434), .ZN(n430) );
  NAND2_X1 U472 ( .A1(n426), .A2(n427), .ZN(n423) );
  XNOR2_X1 U473 ( .A(KEYINPUT33), .B(KEYINPUT71), .ZN(n547) );
  NOR2_X1 U474 ( .A1(n574), .A2(n573), .ZN(n579) );
  XNOR2_X1 U475 ( .A(n452), .B(KEYINPUT74), .ZN(n574) );
  OR2_X1 U476 ( .A1(n583), .A2(n582), .ZN(n595) );
  NOR2_X1 U477 ( .A1(n660), .A2(n566), .ZN(n571) );
  INV_X1 U478 ( .A(KEYINPUT0), .ZN(n448) );
  XNOR2_X1 U479 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U480 ( .A(n477), .B(n456), .ZN(n457) );
  NAND2_X1 U481 ( .A1(n429), .A2(n676), .ZN(n602) );
  XNOR2_X1 U482 ( .A(KEYINPUT105), .B(KEYINPUT40), .ZN(n576) );
  XNOR2_X1 U483 ( .A(n543), .B(KEYINPUT32), .ZN(n739) );
  NOR2_X1 U484 ( .A1(n556), .A2(n555), .ZN(n636) );
  INV_X1 U485 ( .A(n595), .ZN(n637) );
  INV_X1 U486 ( .A(KEYINPUT102), .ZN(n377) );
  NAND2_X1 U487 ( .A1(n403), .A2(n401), .ZN(n546) );
  AND2_X1 U488 ( .A1(n545), .A2(n402), .ZN(n401) );
  INV_X1 U489 ( .A(n636), .ZN(n641) );
  NAND2_X1 U490 ( .A1(n384), .A2(n383), .ZN(n382) );
  INV_X1 U491 ( .A(KEYINPUT81), .ZN(n383) );
  XNOR2_X1 U492 ( .A(n369), .B(n368), .ZN(G63) );
  INV_X1 U493 ( .A(KEYINPUT122), .ZN(n368) );
  XNOR2_X1 U494 ( .A(n367), .B(n366), .ZN(G60) );
  XOR2_X1 U495 ( .A(n523), .B(KEYINPUT86), .Z(n352) );
  OR2_X1 U496 ( .A1(n352), .A2(n613), .ZN(n353) );
  AND2_X1 U497 ( .A1(n411), .A2(n613), .ZN(n354) );
  OR2_X1 U498 ( .A1(n563), .A2(n562), .ZN(n355) );
  XNOR2_X1 U499 ( .A(KEYINPUT78), .B(n609), .ZN(n356) );
  AND2_X1 U500 ( .A1(n411), .A2(n360), .ZN(n358) );
  AND2_X1 U501 ( .A1(n431), .A2(n427), .ZN(n359) );
  AND2_X1 U502 ( .A1(n412), .A2(n610), .ZN(n360) );
  AND2_X1 U503 ( .A1(n396), .A2(KEYINPUT81), .ZN(n361) );
  XOR2_X1 U504 ( .A(KEYINPUT64), .B(KEYINPUT22), .Z(n362) );
  XOR2_X1 U505 ( .A(n614), .B(KEYINPUT65), .Z(n363) );
  XNOR2_X1 U506 ( .A(G902), .B(KEYINPUT15), .ZN(n612) );
  INV_X1 U507 ( .A(n612), .ZN(n613) );
  XOR2_X1 U508 ( .A(n698), .B(n697), .Z(n364) );
  XOR2_X1 U509 ( .A(n708), .B(n707), .Z(n365) );
  XNOR2_X1 U510 ( .A(KEYINPUT84), .B(n621), .ZN(n715) );
  INV_X1 U511 ( .A(n715), .ZN(n392) );
  XNOR2_X1 U512 ( .A(KEYINPUT60), .B(KEYINPUT121), .ZN(n366) );
  NAND2_X1 U513 ( .A1(n352), .A2(n613), .ZN(n380) );
  NAND2_X1 U514 ( .A1(n411), .A2(n400), .ZN(n399) );
  NAND2_X1 U515 ( .A1(n391), .A2(n392), .ZN(n367) );
  NAND2_X1 U516 ( .A1(n393), .A2(n392), .ZN(n369) );
  NOR2_X1 U517 ( .A1(n713), .A2(G902), .ZN(n370) );
  XNOR2_X1 U518 ( .A(n371), .B(n601), .ZN(n607) );
  NAND2_X1 U519 ( .A1(n449), .A2(n451), .ZN(n371) );
  XNOR2_X1 U520 ( .A(n376), .B(G110), .ZN(n738) );
  OR2_X2 U521 ( .A1(n379), .A2(n378), .ZN(n568) );
  NOR2_X1 U522 ( .A1(n696), .A2(n353), .ZN(n378) );
  NAND2_X1 U523 ( .A1(n381), .A2(n380), .ZN(n379) );
  NAND2_X1 U524 ( .A1(n696), .A2(n352), .ZN(n381) );
  XNOR2_X2 U525 ( .A(n409), .B(n522), .ZN(n696) );
  INV_X1 U526 ( .A(n390), .ZN(n384) );
  NAND2_X1 U527 ( .A1(n390), .A2(n361), .ZN(n386) );
  XNOR2_X1 U528 ( .A(n709), .B(n365), .ZN(n391) );
  INV_X1 U529 ( .A(n611), .ZN(n412) );
  XNOR2_X1 U530 ( .A(n450), .B(KEYINPUT46), .ZN(n449) );
  NAND2_X1 U531 ( .A1(n354), .A2(n360), .ZN(n413) );
  XNOR2_X1 U532 ( .A(n710), .B(n394), .ZN(n393) );
  XNOR2_X2 U533 ( .A(n397), .B(n517), .ZN(n409) );
  XNOR2_X1 U534 ( .A(n397), .B(KEYINPUT123), .ZN(n722) );
  XNOR2_X2 U535 ( .A(n514), .B(n513), .ZN(n397) );
  INV_X1 U536 ( .A(n616), .ZN(n656) );
  XNOR2_X2 U537 ( .A(n399), .B(n398), .ZN(n616) );
  INV_X1 U538 ( .A(n544), .ZN(n403) );
  NAND2_X1 U539 ( .A1(n404), .A2(n739), .ZN(n444) );
  NAND2_X1 U540 ( .A1(n405), .A2(n586), .ZN(n587) );
  NAND2_X1 U541 ( .A1(n585), .A2(KEYINPUT47), .ZN(n405) );
  AND2_X1 U542 ( .A1(n600), .A2(n588), .ZN(n451) );
  XNOR2_X1 U543 ( .A(n486), .B(n406), .ZN(n488) );
  NAND2_X1 U544 ( .A1(n626), .A2(n559), .ZN(n442) );
  NAND2_X1 U545 ( .A1(n454), .A2(G478), .ZN(n710) );
  XNOR2_X1 U546 ( .A(n444), .B(KEYINPUT44), .ZN(n443) );
  XNOR2_X1 U547 ( .A(n408), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U548 ( .A1(n700), .A2(n715), .ZN(n408) );
  NOR2_X2 U549 ( .A1(n622), .A2(n715), .ZN(n625) );
  NOR2_X2 U550 ( .A1(n443), .A2(n442), .ZN(n410) );
  NAND2_X1 U551 ( .A1(n538), .A2(G210), .ZN(n419) );
  NAND2_X1 U552 ( .A1(n423), .A2(n422), .ZN(n592) );
  NAND2_X1 U553 ( .A1(n359), .A2(n430), .ZN(n422) );
  NAND2_X1 U554 ( .A1(n430), .A2(n431), .ZN(n424) );
  INV_X1 U555 ( .A(n426), .ZN(n425) );
  INV_X1 U556 ( .A(n591), .ZN(n431) );
  NAND2_X1 U557 ( .A1(n535), .A2(n664), .ZN(n447) );
  XNOR2_X1 U558 ( .A(n446), .B(n539), .ZN(n540) );
  XNOR2_X1 U559 ( .A(n435), .B(KEYINPUT34), .ZN(n548) );
  XNOR2_X2 U560 ( .A(n436), .B(n547), .ZN(n685) );
  NAND2_X1 U561 ( .A1(n551), .A2(n589), .ZN(n436) );
  XNOR2_X2 U562 ( .A(n566), .B(n437), .ZN(n603) );
  XNOR2_X2 U563 ( .A(n439), .B(n438), .ZN(n566) );
  XNOR2_X2 U564 ( .A(n357), .B(n510), .ZN(n446) );
  NAND2_X1 U565 ( .A1(n571), .A2(n355), .ZN(n452) );
  XNOR2_X1 U566 ( .A(n699), .B(n364), .ZN(n700) );
  NAND2_X1 U567 ( .A1(n454), .A2(G210), .ZN(n699) );
  NAND2_X1 U568 ( .A1(n454), .A2(G475), .ZN(n709) );
  XNOR2_X1 U569 ( .A(n577), .B(n576), .ZN(n740) );
  NOR2_X2 U570 ( .A1(n659), .A2(n660), .ZN(n551) );
  XNOR2_X2 U571 ( .A(n516), .B(n475), .ZN(n486) );
  INV_X1 U572 ( .A(n648), .ZN(n599) );
  XNOR2_X1 U573 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U574 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U575 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U576 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U577 ( .A(KEYINPUT75), .B(KEYINPUT19), .ZN(n526) );
  XNOR2_X1 U578 ( .A(n725), .B(n457), .ZN(n469) );
  XNOR2_X1 U579 ( .A(n620), .B(n619), .ZN(n622) );
  XNOR2_X1 U580 ( .A(KEYINPUT10), .B(n455), .ZN(n725) );
  XOR2_X1 U581 ( .A(KEYINPUT70), .B(G110), .Z(n459) );
  XNOR2_X1 U582 ( .A(G128), .B(G119), .ZN(n458) );
  XNOR2_X1 U583 ( .A(n459), .B(n458), .ZN(n463) );
  XOR2_X1 U584 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n461) );
  XNOR2_X1 U585 ( .A(KEYINPUT89), .B(KEYINPUT23), .ZN(n460) );
  XNOR2_X1 U586 ( .A(n461), .B(n460), .ZN(n462) );
  XOR2_X1 U587 ( .A(n463), .B(n462), .Z(n467) );
  NAND2_X1 U588 ( .A1(n720), .A2(G234), .ZN(n465) );
  XNOR2_X1 U589 ( .A(n465), .B(n464), .ZN(n490) );
  NAND2_X1 U590 ( .A1(G221), .A2(n490), .ZN(n466) );
  XNOR2_X1 U591 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U592 ( .A(n469), .B(n468), .ZN(n713) );
  XOR2_X1 U593 ( .A(KEYINPUT25), .B(KEYINPUT76), .Z(n472) );
  NAND2_X1 U594 ( .A1(n612), .A2(G234), .ZN(n470) );
  XNOR2_X1 U595 ( .A(n470), .B(KEYINPUT20), .ZN(n508) );
  NAND2_X1 U596 ( .A1(n508), .A2(G217), .ZN(n471) );
  XNOR2_X1 U597 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U598 ( .A(KEYINPUT77), .B(n473), .ZN(n474) );
  XNOR2_X1 U599 ( .A(n564), .B(KEYINPUT100), .ZN(n663) );
  XOR2_X2 U600 ( .A(G143), .B(G128), .Z(n516) );
  NAND2_X1 U601 ( .A1(G227), .A2(n720), .ZN(n479) );
  INV_X1 U602 ( .A(n603), .ZN(n659) );
  OR2_X1 U603 ( .A1(n663), .A2(n396), .ZN(n483) );
  XNOR2_X1 U604 ( .A(KEYINPUT101), .B(n483), .ZN(n542) );
  XNOR2_X1 U605 ( .A(KEYINPUT97), .B(KEYINPUT95), .ZN(n484) );
  XNOR2_X1 U606 ( .A(n484), .B(KEYINPUT96), .ZN(n489) );
  XOR2_X1 U607 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n487) );
  XOR2_X1 U608 ( .A(n489), .B(n488), .Z(n492) );
  NAND2_X1 U609 ( .A1(G217), .A2(n490), .ZN(n491) );
  NOR2_X1 U610 ( .A1(G902), .A2(n711), .ZN(n493) );
  XNOR2_X1 U611 ( .A(n493), .B(G478), .ZN(n554) );
  XOR2_X1 U612 ( .A(KEYINPUT12), .B(G140), .Z(n495) );
  XNOR2_X1 U613 ( .A(n495), .B(n494), .ZN(n503) );
  NAND2_X1 U614 ( .A1(n538), .A2(G214), .ZN(n496) );
  XNOR2_X1 U615 ( .A(n497), .B(n496), .ZN(n501) );
  XNOR2_X1 U616 ( .A(n503), .B(n502), .ZN(n504) );
  NOR2_X1 U617 ( .A1(G902), .A2(n708), .ZN(n506) );
  XNOR2_X1 U618 ( .A(KEYINPUT94), .B(KEYINPUT13), .ZN(n505) );
  XNOR2_X1 U619 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X2 U620 ( .A(G475), .B(n507), .Z(n555) );
  NAND2_X1 U621 ( .A1(n554), .A2(n555), .ZN(n679) );
  INV_X1 U622 ( .A(n679), .ZN(n535) );
  NAND2_X1 U623 ( .A1(G221), .A2(n508), .ZN(n509) );
  XOR2_X1 U624 ( .A(KEYINPUT21), .B(n509), .Z(n664) );
  XNOR2_X1 U625 ( .A(n512), .B(KEYINPUT16), .ZN(n513) );
  AND2_X1 U626 ( .A1(G224), .A2(n720), .ZN(n515) );
  XNOR2_X1 U627 ( .A(n518), .B(KEYINPUT18), .ZN(n519) );
  XOR2_X1 U628 ( .A(n519), .B(KEYINPUT4), .Z(n521) );
  XNOR2_X1 U629 ( .A(KEYINPUT85), .B(KEYINPUT17), .ZN(n520) );
  NAND2_X1 U630 ( .A1(G210), .A2(n524), .ZN(n523) );
  NAND2_X1 U631 ( .A1(G214), .A2(n524), .ZN(n525) );
  XNOR2_X1 U632 ( .A(KEYINPUT14), .B(n528), .ZN(n530) );
  NAND2_X1 U633 ( .A1(n530), .A2(G952), .ZN(n529) );
  XNOR2_X1 U634 ( .A(n529), .B(KEYINPUT88), .ZN(n691) );
  NOR2_X1 U635 ( .A1(G953), .A2(n691), .ZN(n563) );
  AND2_X1 U636 ( .A1(G953), .A2(n530), .ZN(n531) );
  NAND2_X1 U637 ( .A1(G902), .A2(n531), .ZN(n560) );
  NOR2_X1 U638 ( .A1(G898), .A2(n560), .ZN(n532) );
  NOR2_X1 U639 ( .A1(n563), .A2(n532), .ZN(n533) );
  NOR2_X2 U640 ( .A1(n582), .A2(n533), .ZN(n534) );
  INV_X1 U641 ( .A(n536), .ZN(n541) );
  NAND2_X1 U642 ( .A1(n542), .A2(n549), .ZN(n543) );
  NOR2_X1 U643 ( .A1(n603), .A2(n564), .ZN(n545) );
  NOR2_X1 U644 ( .A1(n555), .A2(n554), .ZN(n578) );
  NOR2_X1 U645 ( .A1(n667), .A2(n351), .ZN(n550) );
  NAND2_X1 U646 ( .A1(n571), .A2(n550), .ZN(n628) );
  NAND2_X1 U647 ( .A1(n667), .A2(n551), .ZN(n670) );
  NOR2_X1 U648 ( .A1(n670), .A2(n351), .ZN(n553) );
  XNOR2_X1 U649 ( .A(n553), .B(KEYINPUT31), .ZN(n643) );
  NAND2_X1 U650 ( .A1(n628), .A2(n643), .ZN(n558) );
  INV_X1 U651 ( .A(n554), .ZN(n556) );
  NAND2_X1 U652 ( .A1(n556), .A2(n555), .ZN(n644) );
  NAND2_X1 U653 ( .A1(n641), .A2(n644), .ZN(n557) );
  NAND2_X1 U654 ( .A1(n558), .A2(n680), .ZN(n559) );
  XOR2_X1 U655 ( .A(KEYINPUT68), .B(KEYINPUT48), .Z(n601) );
  XOR2_X1 U656 ( .A(n560), .B(KEYINPUT103), .Z(n561) );
  NOR2_X1 U657 ( .A1(G900), .A2(n561), .ZN(n562) );
  AND2_X1 U658 ( .A1(n590), .A2(n667), .ZN(n565) );
  INV_X1 U659 ( .A(n566), .ZN(n567) );
  INV_X1 U660 ( .A(n568), .ZN(n605) );
  XNOR2_X1 U661 ( .A(KEYINPUT41), .B(KEYINPUT106), .ZN(n569) );
  NOR2_X1 U662 ( .A1(n583), .A2(n674), .ZN(n570) );
  XNOR2_X1 U663 ( .A(n570), .B(KEYINPUT42), .ZN(n742) );
  AND2_X1 U664 ( .A1(n676), .A2(n667), .ZN(n572) );
  XOR2_X1 U665 ( .A(KEYINPUT30), .B(n572), .Z(n573) );
  NAND2_X1 U666 ( .A1(n675), .A2(n579), .ZN(n575) );
  NAND2_X1 U667 ( .A1(n608), .A2(n636), .ZN(n577) );
  NAND2_X1 U668 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U669 ( .A1(n605), .A2(n580), .ZN(n635) );
  NAND2_X1 U670 ( .A1(KEYINPUT79), .A2(n680), .ZN(n586) );
  INV_X1 U671 ( .A(KEYINPUT79), .ZN(n581) );
  NAND2_X1 U672 ( .A1(n594), .A2(n581), .ZN(n584) );
  NAND2_X1 U673 ( .A1(n584), .A2(n637), .ZN(n585) );
  NOR2_X1 U674 ( .A1(n635), .A2(n587), .ZN(n588) );
  NAND2_X1 U675 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U676 ( .A(n592), .B(KEYINPUT36), .ZN(n593) );
  NAND2_X1 U677 ( .A1(n593), .A2(n603), .ZN(n648) );
  NOR2_X1 U678 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U679 ( .A1(n596), .A2(KEYINPUT79), .ZN(n597) );
  NOR2_X1 U680 ( .A1(KEYINPUT47), .A2(n597), .ZN(n598) );
  NOR2_X1 U681 ( .A1(n599), .A2(n598), .ZN(n600) );
  OR2_X1 U682 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U683 ( .A(KEYINPUT43), .B(n604), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n606), .A2(n605), .ZN(n651) );
  NAND2_X1 U685 ( .A1(n607), .A2(n651), .ZN(n611) );
  INV_X1 U686 ( .A(n644), .ZN(n632) );
  NAND2_X1 U687 ( .A1(n608), .A2(n632), .ZN(n610) );
  NAND2_X1 U688 ( .A1(KEYINPUT2), .A2(n610), .ZN(n609) );
  INV_X1 U689 ( .A(n610), .ZN(n649) );
  NAND2_X1 U690 ( .A1(n613), .A2(KEYINPUT2), .ZN(n614) );
  NAND2_X1 U691 ( .A1(n454), .A2(G472), .ZN(n620) );
  XOR2_X1 U692 ( .A(KEYINPUT62), .B(KEYINPUT107), .Z(n617) );
  NOR2_X1 U693 ( .A1(G952), .A2(n720), .ZN(n621) );
  XOR2_X1 U694 ( .A(KEYINPUT63), .B(KEYINPUT108), .Z(n623) );
  XNOR2_X1 U695 ( .A(KEYINPUT82), .B(n623), .ZN(n624) );
  XNOR2_X1 U696 ( .A(n625), .B(n624), .ZN(G57) );
  XNOR2_X1 U697 ( .A(n626), .B(G101), .ZN(G3) );
  NOR2_X1 U698 ( .A1(n641), .A2(n628), .ZN(n627) );
  XOR2_X1 U699 ( .A(G104), .B(n627), .Z(G6) );
  NOR2_X1 U700 ( .A1(n644), .A2(n628), .ZN(n630) );
  XNOR2_X1 U701 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n629) );
  XNOR2_X1 U702 ( .A(n630), .B(n629), .ZN(n631) );
  XNOR2_X1 U703 ( .A(G107), .B(n631), .ZN(G9) );
  XOR2_X1 U704 ( .A(G128), .B(KEYINPUT29), .Z(n634) );
  NAND2_X1 U705 ( .A1(n632), .A2(n637), .ZN(n633) );
  XNOR2_X1 U706 ( .A(n634), .B(n633), .ZN(G30) );
  XOR2_X1 U707 ( .A(G143), .B(n635), .Z(G45) );
  XOR2_X1 U708 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n639) );
  NAND2_X1 U709 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U710 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U711 ( .A(G146), .B(n640), .ZN(G48) );
  NOR2_X1 U712 ( .A1(n641), .A2(n643), .ZN(n642) );
  XOR2_X1 U713 ( .A(G113), .B(n642), .Z(G15) );
  NOR2_X1 U714 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U715 ( .A(KEYINPUT112), .B(n645), .Z(n646) );
  XNOR2_X1 U716 ( .A(G116), .B(n646), .ZN(G18) );
  XOR2_X1 U717 ( .A(G125), .B(KEYINPUT37), .Z(n647) );
  XNOR2_X1 U718 ( .A(n648), .B(n647), .ZN(G27) );
  XNOR2_X1 U719 ( .A(G134), .B(n649), .ZN(n650) );
  XNOR2_X1 U720 ( .A(n650), .B(KEYINPUT113), .ZN(G36) );
  XNOR2_X1 U721 ( .A(G140), .B(KEYINPUT114), .ZN(n652) );
  XNOR2_X1 U722 ( .A(n652), .B(n651), .ZN(G42) );
  NOR2_X1 U723 ( .A1(n685), .A2(n674), .ZN(n653) );
  XOR2_X1 U724 ( .A(KEYINPUT118), .B(n653), .Z(n654) );
  NAND2_X1 U725 ( .A1(n720), .A2(n654), .ZN(n658) );
  NOR2_X1 U726 ( .A1(n358), .A2(KEYINPUT2), .ZN(n655) );
  NOR2_X1 U727 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U728 ( .A1(n658), .A2(n657), .ZN(n694) );
  NAND2_X1 U729 ( .A1(n660), .A2(n396), .ZN(n661) );
  XOR2_X1 U730 ( .A(KEYINPUT50), .B(n661), .Z(n662) );
  XNOR2_X1 U731 ( .A(n662), .B(KEYINPUT115), .ZN(n669) );
  NOR2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U733 ( .A(KEYINPUT49), .B(n665), .Z(n666) );
  NOR2_X1 U734 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U735 ( .A1(n669), .A2(n668), .ZN(n671) );
  NAND2_X1 U736 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U737 ( .A(KEYINPUT51), .B(n672), .ZN(n673) );
  NOR2_X1 U738 ( .A1(n674), .A2(n673), .ZN(n688) );
  NOR2_X1 U739 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U740 ( .A(n677), .B(KEYINPUT116), .ZN(n678) );
  NOR2_X1 U741 ( .A1(n679), .A2(n678), .ZN(n684) );
  INV_X1 U742 ( .A(n680), .ZN(n682) );
  NOR2_X1 U743 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U744 ( .A1(n684), .A2(n683), .ZN(n686) );
  NOR2_X1 U745 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U746 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U747 ( .A(KEYINPUT52), .B(n689), .ZN(n690) );
  NOR2_X1 U748 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U749 ( .A(n692), .B(KEYINPUT117), .ZN(n693) );
  NAND2_X1 U750 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U751 ( .A(KEYINPUT53), .B(n695), .Z(G75) );
  XOR2_X1 U752 ( .A(KEYINPUT83), .B(KEYINPUT55), .Z(n698) );
  XNOR2_X1 U753 ( .A(n696), .B(KEYINPUT54), .ZN(n697) );
  XOR2_X1 U754 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n703) );
  XNOR2_X1 U755 ( .A(n701), .B(KEYINPUT119), .ZN(n702) );
  XNOR2_X1 U756 ( .A(n703), .B(n702), .ZN(n705) );
  NAND2_X1 U757 ( .A1(n454), .A2(G469), .ZN(n704) );
  XOR2_X1 U758 ( .A(n705), .B(n704), .Z(n706) );
  NOR2_X1 U759 ( .A1(n715), .A2(n706), .ZN(G54) );
  XOR2_X1 U760 ( .A(KEYINPUT120), .B(KEYINPUT59), .Z(n707) );
  NAND2_X1 U761 ( .A1(G217), .A2(n454), .ZN(n712) );
  XNOR2_X1 U762 ( .A(n713), .B(n712), .ZN(n714) );
  NOR2_X1 U763 ( .A1(n715), .A2(n714), .ZN(G66) );
  NAND2_X1 U764 ( .A1(n720), .A2(n411), .ZN(n719) );
  NAND2_X1 U765 ( .A1(G953), .A2(G224), .ZN(n716) );
  XNOR2_X1 U766 ( .A(KEYINPUT61), .B(n716), .ZN(n717) );
  NAND2_X1 U767 ( .A1(n717), .A2(G898), .ZN(n718) );
  NAND2_X1 U768 ( .A1(n719), .A2(n718), .ZN(n724) );
  NOR2_X1 U769 ( .A1(n720), .A2(G898), .ZN(n721) );
  NOR2_X1 U770 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U771 ( .A(n724), .B(n723), .ZN(G69) );
  XNOR2_X1 U772 ( .A(n726), .B(n725), .ZN(n727) );
  XNOR2_X1 U773 ( .A(n727), .B(KEYINPUT124), .ZN(n732) );
  INV_X1 U774 ( .A(n732), .ZN(n728) );
  XNOR2_X1 U775 ( .A(KEYINPUT126), .B(n728), .ZN(n729) );
  XNOR2_X1 U776 ( .A(G227), .B(n729), .ZN(n730) );
  NAND2_X1 U777 ( .A1(n730), .A2(G900), .ZN(n731) );
  NAND2_X1 U778 ( .A1(n731), .A2(G953), .ZN(n736) );
  XOR2_X1 U779 ( .A(n360), .B(n732), .Z(n733) );
  NOR2_X1 U780 ( .A1(G953), .A2(n733), .ZN(n734) );
  XNOR2_X1 U781 ( .A(KEYINPUT125), .B(n734), .ZN(n735) );
  NAND2_X1 U782 ( .A1(n736), .A2(n735), .ZN(G72) );
  XOR2_X1 U783 ( .A(n737), .B(G122), .Z(G24) );
  XNOR2_X1 U784 ( .A(KEYINPUT109), .B(n738), .ZN(G12) );
  XNOR2_X1 U785 ( .A(n739), .B(G119), .ZN(G21) );
  XNOR2_X1 U786 ( .A(G131), .B(KEYINPUT127), .ZN(n741) );
  XNOR2_X1 U787 ( .A(n741), .B(n740), .ZN(G33) );
  XOR2_X1 U788 ( .A(G137), .B(n742), .Z(G39) );
endmodule

