

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U548 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U549 ( .A1(n774), .A2(n691), .ZN(n735) );
  AND2_X1 U550 ( .A1(n690), .A2(n689), .ZN(n697) );
  XOR2_X1 U551 ( .A(G2104), .B(KEYINPUT64), .Z(n515) );
  XNOR2_X1 U552 ( .A(KEYINPUT23), .B(KEYINPUT65), .ZN(n535) );
  XNOR2_X1 U553 ( .A(n688), .B(n687), .ZN(n690) );
  NOR2_X1 U554 ( .A1(n542), .A2(n541), .ZN(G160) );
  INV_X1 U555 ( .A(G168), .ZN(n689) );
  INV_X1 U556 ( .A(n773), .ZN(n691) );
  NOR2_X1 U557 ( .A1(G651), .A2(G543), .ZN(n642) );
  NOR2_X1 U558 ( .A1(G651), .A2(n638), .ZN(n647) );
  XNOR2_X1 U559 ( .A(n536), .B(n535), .ZN(n538) );
  AND2_X1 U560 ( .A1(G2105), .A2(G2104), .ZN(n889) );
  NAND2_X1 U561 ( .A1(G114), .A2(n889), .ZN(n513) );
  AND2_X1 U562 ( .A1(G2105), .A2(n515), .ZN(n886) );
  NAND2_X1 U563 ( .A1(G126), .A2(n886), .ZN(n512) );
  AND2_X1 U564 ( .A1(n513), .A2(n512), .ZN(n520) );
  NOR2_X1 U565 ( .A1(G2105), .A2(G2104), .ZN(n514) );
  XOR2_X2 U566 ( .A(KEYINPUT17), .B(n514), .Z(n882) );
  NAND2_X1 U567 ( .A1(n882), .A2(G138), .ZN(n517) );
  NOR2_X4 U568 ( .A1(n515), .A2(G2105), .ZN(n881) );
  NAND2_X1 U569 ( .A1(n881), .A2(G102), .ZN(n516) );
  NAND2_X1 U570 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U571 ( .A(KEYINPUT87), .B(n518), .ZN(n519) );
  AND2_X2 U572 ( .A1(n520), .A2(n519), .ZN(G164) );
  INV_X1 U573 ( .A(G651), .ZN(n527) );
  NOR2_X1 U574 ( .A1(G543), .A2(n527), .ZN(n521) );
  XOR2_X1 U575 ( .A(KEYINPUT1), .B(n521), .Z(n646) );
  NAND2_X1 U576 ( .A1(G63), .A2(n646), .ZN(n523) );
  XOR2_X1 U577 ( .A(KEYINPUT0), .B(G543), .Z(n638) );
  NAND2_X1 U578 ( .A1(G51), .A2(n647), .ZN(n522) );
  NAND2_X1 U579 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U580 ( .A(KEYINPUT6), .B(n524), .ZN(n533) );
  NAND2_X1 U581 ( .A1(G89), .A2(n642), .ZN(n525) );
  XNOR2_X1 U582 ( .A(n525), .B(KEYINPUT4), .ZN(n526) );
  XNOR2_X1 U583 ( .A(n526), .B(KEYINPUT74), .ZN(n529) );
  NOR2_X1 U584 ( .A1(n638), .A2(n527), .ZN(n643) );
  NAND2_X1 U585 ( .A1(G76), .A2(n643), .ZN(n528) );
  NAND2_X1 U586 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U587 ( .A(KEYINPUT5), .B(n530), .ZN(n531) );
  XNOR2_X1 U588 ( .A(KEYINPUT75), .B(n531), .ZN(n532) );
  NOR2_X1 U589 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U590 ( .A(KEYINPUT7), .B(n534), .Z(G168) );
  NAND2_X1 U591 ( .A1(G101), .A2(n881), .ZN(n536) );
  NAND2_X1 U592 ( .A1(G113), .A2(n889), .ZN(n537) );
  NAND2_X1 U593 ( .A1(n538), .A2(n537), .ZN(n542) );
  NAND2_X1 U594 ( .A1(G137), .A2(n882), .ZN(n540) );
  NAND2_X1 U595 ( .A1(G125), .A2(n886), .ZN(n539) );
  NAND2_X1 U596 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U597 ( .A1(G65), .A2(n646), .ZN(n544) );
  NAND2_X1 U598 ( .A1(G91), .A2(n642), .ZN(n543) );
  NAND2_X1 U599 ( .A1(n544), .A2(n543), .ZN(n548) );
  NAND2_X1 U600 ( .A1(G78), .A2(n643), .ZN(n546) );
  NAND2_X1 U601 ( .A1(G53), .A2(n647), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n546), .A2(n545), .ZN(n547) );
  OR2_X1 U603 ( .A1(n548), .A2(n547), .ZN(G299) );
  NAND2_X1 U604 ( .A1(G85), .A2(n642), .ZN(n550) );
  NAND2_X1 U605 ( .A1(G72), .A2(n643), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U607 ( .A1(G60), .A2(n646), .ZN(n552) );
  NAND2_X1 U608 ( .A1(G47), .A2(n647), .ZN(n551) );
  NAND2_X1 U609 ( .A1(n552), .A2(n551), .ZN(n553) );
  OR2_X1 U610 ( .A1(n554), .A2(n553), .ZN(G290) );
  XOR2_X1 U611 ( .A(G2443), .B(G2451), .Z(n556) );
  XNOR2_X1 U612 ( .A(G2430), .B(G2427), .ZN(n555) );
  XNOR2_X1 U613 ( .A(n556), .B(n555), .ZN(n560) );
  XOR2_X1 U614 ( .A(KEYINPUT110), .B(G2438), .Z(n558) );
  XNOR2_X1 U615 ( .A(G2435), .B(G2454), .ZN(n557) );
  XNOR2_X1 U616 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U617 ( .A(n560), .B(n559), .Z(n562) );
  XNOR2_X1 U618 ( .A(G2446), .B(KEYINPUT108), .ZN(n561) );
  XNOR2_X1 U619 ( .A(n562), .B(n561), .ZN(n565) );
  XOR2_X1 U620 ( .A(G1341), .B(G1348), .Z(n563) );
  XNOR2_X1 U621 ( .A(KEYINPUT109), .B(n563), .ZN(n564) );
  XOR2_X1 U622 ( .A(n565), .B(n564), .Z(n566) );
  AND2_X1 U623 ( .A1(G14), .A2(n566), .ZN(G401) );
  NAND2_X1 U624 ( .A1(G64), .A2(n646), .ZN(n568) );
  NAND2_X1 U625 ( .A1(G52), .A2(n647), .ZN(n567) );
  NAND2_X1 U626 ( .A1(n568), .A2(n567), .ZN(n573) );
  NAND2_X1 U627 ( .A1(G90), .A2(n642), .ZN(n570) );
  NAND2_X1 U628 ( .A1(G77), .A2(n643), .ZN(n569) );
  NAND2_X1 U629 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U630 ( .A(KEYINPUT9), .B(n571), .Z(n572) );
  NOR2_X1 U631 ( .A1(n573), .A2(n572), .ZN(G171) );
  AND2_X1 U632 ( .A1(G452), .A2(G94), .ZN(G173) );
  XOR2_X1 U633 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U634 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n575) );
  NAND2_X1 U635 ( .A1(G7), .A2(G661), .ZN(n574) );
  XNOR2_X1 U636 ( .A(n575), .B(n574), .ZN(G223) );
  XOR2_X1 U637 ( .A(G223), .B(KEYINPUT70), .Z(n826) );
  NAND2_X1 U638 ( .A1(n826), .A2(G567), .ZN(n576) );
  XNOR2_X1 U639 ( .A(n576), .B(KEYINPUT71), .ZN(n577) );
  XNOR2_X1 U640 ( .A(KEYINPUT11), .B(n577), .ZN(G234) );
  XOR2_X1 U641 ( .A(KEYINPUT72), .B(KEYINPUT14), .Z(n579) );
  NAND2_X1 U642 ( .A1(G56), .A2(n646), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(n585) );
  NAND2_X1 U644 ( .A1(n642), .A2(G81), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(KEYINPUT12), .ZN(n582) );
  NAND2_X1 U646 ( .A1(G68), .A2(n643), .ZN(n581) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U648 ( .A(KEYINPUT13), .B(n583), .Z(n584) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n587) );
  NAND2_X1 U650 ( .A1(n647), .A2(G43), .ZN(n586) );
  NAND2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n943) );
  INV_X1 U652 ( .A(G860), .ZN(n600) );
  OR2_X1 U653 ( .A1(n943), .A2(n600), .ZN(G153) );
  INV_X1 U654 ( .A(G868), .ZN(n661) );
  NOR2_X1 U655 ( .A1(n661), .A2(G171), .ZN(n588) );
  XNOR2_X1 U656 ( .A(n588), .B(KEYINPUT73), .ZN(n597) );
  NAND2_X1 U657 ( .A1(G79), .A2(n643), .ZN(n590) );
  NAND2_X1 U658 ( .A1(G54), .A2(n647), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U660 ( .A1(G66), .A2(n646), .ZN(n592) );
  NAND2_X1 U661 ( .A1(G92), .A2(n642), .ZN(n591) );
  NAND2_X1 U662 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U663 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U664 ( .A(n595), .B(KEYINPUT15), .ZN(n940) );
  NAND2_X1 U665 ( .A1(n661), .A2(n940), .ZN(n596) );
  NAND2_X1 U666 ( .A1(n597), .A2(n596), .ZN(G284) );
  NOR2_X1 U667 ( .A1(G286), .A2(n661), .ZN(n599) );
  NOR2_X1 U668 ( .A1(G868), .A2(G299), .ZN(n598) );
  NOR2_X1 U669 ( .A1(n599), .A2(n598), .ZN(G297) );
  NAND2_X1 U670 ( .A1(n600), .A2(G559), .ZN(n601) );
  INV_X1 U671 ( .A(n940), .ZN(n897) );
  NAND2_X1 U672 ( .A1(n601), .A2(n897), .ZN(n602) );
  XNOR2_X1 U673 ( .A(n602), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U674 ( .A1(G868), .A2(n943), .ZN(n603) );
  XNOR2_X1 U675 ( .A(KEYINPUT76), .B(n603), .ZN(n606) );
  NAND2_X1 U676 ( .A1(G868), .A2(n897), .ZN(n604) );
  NOR2_X1 U677 ( .A1(G559), .A2(n604), .ZN(n605) );
  NOR2_X1 U678 ( .A1(n606), .A2(n605), .ZN(G282) );
  NAND2_X1 U679 ( .A1(G111), .A2(n889), .ZN(n613) );
  NAND2_X1 U680 ( .A1(G99), .A2(n881), .ZN(n608) );
  NAND2_X1 U681 ( .A1(G135), .A2(n882), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U683 ( .A1(n886), .A2(G123), .ZN(n609) );
  XOR2_X1 U684 ( .A(KEYINPUT18), .B(n609), .Z(n610) );
  NOR2_X1 U685 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U687 ( .A(n614), .B(KEYINPUT77), .ZN(n919) );
  XNOR2_X1 U688 ( .A(n919), .B(G2096), .ZN(n616) );
  INV_X1 U689 ( .A(G2100), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n616), .A2(n615), .ZN(G156) );
  NAND2_X1 U691 ( .A1(G93), .A2(n642), .ZN(n617) );
  XNOR2_X1 U692 ( .A(n617), .B(KEYINPUT78), .ZN(n624) );
  NAND2_X1 U693 ( .A1(G80), .A2(n643), .ZN(n619) );
  NAND2_X1 U694 ( .A1(G55), .A2(n647), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U696 ( .A1(G67), .A2(n646), .ZN(n620) );
  XNOR2_X1 U697 ( .A(KEYINPUT79), .B(n620), .ZN(n621) );
  NOR2_X1 U698 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U699 ( .A1(n624), .A2(n623), .ZN(n662) );
  NAND2_X1 U700 ( .A1(n897), .A2(G559), .ZN(n658) );
  XNOR2_X1 U701 ( .A(n943), .B(n658), .ZN(n625) );
  NOR2_X1 U702 ( .A1(G860), .A2(n625), .ZN(n626) );
  XOR2_X1 U703 ( .A(n662), .B(n626), .Z(G145) );
  NAND2_X1 U704 ( .A1(G61), .A2(n646), .ZN(n628) );
  NAND2_X1 U705 ( .A1(G86), .A2(n642), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U707 ( .A1(n643), .A2(G73), .ZN(n629) );
  XOR2_X1 U708 ( .A(KEYINPUT2), .B(n629), .Z(n630) );
  NOR2_X1 U709 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n647), .A2(G48), .ZN(n632) );
  NAND2_X1 U711 ( .A1(n633), .A2(n632), .ZN(G305) );
  NAND2_X1 U712 ( .A1(G49), .A2(n647), .ZN(n635) );
  NAND2_X1 U713 ( .A1(G74), .A2(G651), .ZN(n634) );
  NAND2_X1 U714 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U715 ( .A1(n646), .A2(n636), .ZN(n637) );
  XNOR2_X1 U716 ( .A(n637), .B(KEYINPUT80), .ZN(n640) );
  NAND2_X1 U717 ( .A1(G87), .A2(n638), .ZN(n639) );
  NAND2_X1 U718 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U719 ( .A(KEYINPUT81), .B(n641), .Z(G288) );
  NAND2_X1 U720 ( .A1(G88), .A2(n642), .ZN(n645) );
  NAND2_X1 U721 ( .A1(G75), .A2(n643), .ZN(n644) );
  NAND2_X1 U722 ( .A1(n645), .A2(n644), .ZN(n651) );
  NAND2_X1 U723 ( .A1(G62), .A2(n646), .ZN(n649) );
  NAND2_X1 U724 ( .A1(G50), .A2(n647), .ZN(n648) );
  NAND2_X1 U725 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U726 ( .A1(n651), .A2(n650), .ZN(G166) );
  XNOR2_X1 U727 ( .A(KEYINPUT19), .B(G290), .ZN(n652) );
  XNOR2_X1 U728 ( .A(n652), .B(G299), .ZN(n655) );
  XOR2_X1 U729 ( .A(G305), .B(G288), .Z(n653) );
  XNOR2_X1 U730 ( .A(n662), .B(n653), .ZN(n654) );
  XNOR2_X1 U731 ( .A(n655), .B(n654), .ZN(n657) );
  XNOR2_X1 U732 ( .A(n943), .B(G166), .ZN(n656) );
  XNOR2_X1 U733 ( .A(n657), .B(n656), .ZN(n899) );
  XOR2_X1 U734 ( .A(n899), .B(n658), .Z(n659) );
  NAND2_X1 U735 ( .A1(G868), .A2(n659), .ZN(n660) );
  XNOR2_X1 U736 ( .A(KEYINPUT82), .B(n660), .ZN(n665) );
  NAND2_X1 U737 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U738 ( .A(KEYINPUT83), .B(n663), .Z(n664) );
  NAND2_X1 U739 ( .A1(n665), .A2(n664), .ZN(G295) );
  NAND2_X1 U740 ( .A1(G2084), .A2(G2078), .ZN(n667) );
  XOR2_X1 U741 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n666) );
  XNOR2_X1 U742 ( .A(n667), .B(n666), .ZN(n668) );
  NAND2_X1 U743 ( .A1(G2090), .A2(n668), .ZN(n669) );
  XNOR2_X1 U744 ( .A(KEYINPUT21), .B(n669), .ZN(n670) );
  NAND2_X1 U745 ( .A1(n670), .A2(G2072), .ZN(G158) );
  XOR2_X1 U746 ( .A(KEYINPUT66), .B(G57), .Z(G237) );
  XNOR2_X1 U747 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U748 ( .A(KEYINPUT68), .B(G82), .Z(G220) );
  XNOR2_X1 U749 ( .A(KEYINPUT67), .B(G132), .ZN(G219) );
  NAND2_X1 U750 ( .A1(G108), .A2(G120), .ZN(n671) );
  NOR2_X1 U751 ( .A1(G237), .A2(n671), .ZN(n672) );
  NAND2_X1 U752 ( .A1(G69), .A2(n672), .ZN(n909) );
  NAND2_X1 U753 ( .A1(n909), .A2(G567), .ZN(n677) );
  NOR2_X1 U754 ( .A1(G220), .A2(G219), .ZN(n673) );
  XOR2_X1 U755 ( .A(KEYINPUT22), .B(n673), .Z(n674) );
  NOR2_X1 U756 ( .A1(G218), .A2(n674), .ZN(n675) );
  NAND2_X1 U757 ( .A1(G96), .A2(n675), .ZN(n910) );
  NAND2_X1 U758 ( .A1(n910), .A2(G2106), .ZN(n676) );
  NAND2_X1 U759 ( .A1(n677), .A2(n676), .ZN(n832) );
  NAND2_X1 U760 ( .A1(G483), .A2(G661), .ZN(n678) );
  NOR2_X1 U761 ( .A1(n832), .A2(n678), .ZN(n679) );
  XOR2_X1 U762 ( .A(KEYINPUT85), .B(n679), .Z(n831) );
  NAND2_X1 U763 ( .A1(G36), .A2(n831), .ZN(n680) );
  XNOR2_X1 U764 ( .A(n680), .B(KEYINPUT86), .ZN(G176) );
  INV_X1 U765 ( .A(G166), .ZN(G303) );
  NOR2_X1 U766 ( .A1(G164), .A2(G1384), .ZN(n774) );
  NAND2_X1 U767 ( .A1(G160), .A2(G40), .ZN(n773) );
  NAND2_X2 U768 ( .A1(G8), .A2(n735), .ZN(n769) );
  NOR2_X1 U769 ( .A1(G1981), .A2(G305), .ZN(n681) );
  XOR2_X1 U770 ( .A(n681), .B(KEYINPUT24), .Z(n682) );
  NOR2_X1 U771 ( .A1(n769), .A2(n682), .ZN(n764) );
  NOR2_X1 U772 ( .A1(G1966), .A2(n769), .ZN(n683) );
  XOR2_X1 U773 ( .A(n683), .B(KEYINPUT93), .Z(n730) );
  NOR2_X1 U774 ( .A1(G2084), .A2(n735), .ZN(n728) );
  INV_X1 U775 ( .A(G8), .ZN(n684) );
  OR2_X1 U776 ( .A1(n728), .A2(n684), .ZN(n685) );
  OR2_X2 U777 ( .A1(n730), .A2(n685), .ZN(n688) );
  XNOR2_X1 U778 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n686) );
  XNOR2_X1 U779 ( .A(n686), .B(KEYINPUT30), .ZN(n687) );
  AND2_X1 U780 ( .A1(n774), .A2(n691), .ZN(n710) );
  NOR2_X1 U781 ( .A1(n710), .A2(G1961), .ZN(n692) );
  XNOR2_X1 U782 ( .A(n692), .B(KEYINPUT94), .ZN(n694) );
  XOR2_X1 U783 ( .A(G2078), .B(KEYINPUT25), .Z(n992) );
  NOR2_X1 U784 ( .A1(n735), .A2(n992), .ZN(n693) );
  NOR2_X1 U785 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U786 ( .A(KEYINPUT95), .B(n695), .ZN(n723) );
  NOR2_X1 U787 ( .A1(G171), .A2(n723), .ZN(n696) );
  OR2_X1 U788 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U789 ( .A(n698), .B(KEYINPUT31), .ZN(n727) );
  NAND2_X1 U790 ( .A1(G1348), .A2(n735), .ZN(n700) );
  NAND2_X1 U791 ( .A1(G2067), .A2(n710), .ZN(n699) );
  NAND2_X1 U792 ( .A1(n700), .A2(n699), .ZN(n707) );
  NOR2_X1 U793 ( .A1(n940), .A2(n707), .ZN(n706) );
  AND2_X1 U794 ( .A1(n710), .A2(G1996), .ZN(n701) );
  XOR2_X1 U795 ( .A(n701), .B(KEYINPUT26), .Z(n703) );
  NAND2_X1 U796 ( .A1(n735), .A2(G1341), .ZN(n702) );
  NAND2_X1 U797 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U798 ( .A1(n704), .A2(n943), .ZN(n705) );
  NOR2_X1 U799 ( .A1(n706), .A2(n705), .ZN(n709) );
  AND2_X1 U800 ( .A1(n940), .A2(n707), .ZN(n708) );
  NOR2_X1 U801 ( .A1(n709), .A2(n708), .ZN(n716) );
  NAND2_X1 U802 ( .A1(n710), .A2(G2072), .ZN(n711) );
  XOR2_X1 U803 ( .A(KEYINPUT27), .B(n711), .Z(n713) );
  XNOR2_X1 U804 ( .A(G1956), .B(KEYINPUT96), .ZN(n965) );
  NAND2_X1 U805 ( .A1(n735), .A2(n965), .ZN(n712) );
  NAND2_X1 U806 ( .A1(n713), .A2(n712), .ZN(n717) );
  NOR2_X1 U807 ( .A1(G299), .A2(n717), .ZN(n714) );
  XNOR2_X1 U808 ( .A(n714), .B(KEYINPUT98), .ZN(n715) );
  NOR2_X1 U809 ( .A1(n716), .A2(n715), .ZN(n721) );
  NAND2_X1 U810 ( .A1(n717), .A2(G299), .ZN(n718) );
  XNOR2_X1 U811 ( .A(n718), .B(KEYINPUT97), .ZN(n719) );
  XNOR2_X1 U812 ( .A(n719), .B(KEYINPUT28), .ZN(n720) );
  XNOR2_X1 U813 ( .A(n722), .B(KEYINPUT29), .ZN(n725) );
  NAND2_X1 U814 ( .A1(G171), .A2(n723), .ZN(n724) );
  NAND2_X1 U815 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U816 ( .A1(n727), .A2(n726), .ZN(n734) );
  XNOR2_X1 U817 ( .A(n734), .B(KEYINPUT101), .ZN(n732) );
  AND2_X1 U818 ( .A1(G8), .A2(n728), .ZN(n729) );
  OR2_X1 U819 ( .A1(n730), .A2(n729), .ZN(n731) );
  OR2_X1 U820 ( .A1(n732), .A2(n731), .ZN(n744) );
  AND2_X1 U821 ( .A1(G286), .A2(G8), .ZN(n733) );
  NAND2_X1 U822 ( .A1(n734), .A2(n733), .ZN(n741) );
  NOR2_X1 U823 ( .A1(G1971), .A2(n769), .ZN(n737) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n735), .ZN(n736) );
  NOR2_X1 U825 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U826 ( .A1(n738), .A2(G303), .ZN(n739) );
  OR2_X1 U827 ( .A1(n684), .A2(n739), .ZN(n740) );
  AND2_X1 U828 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U829 ( .A(n742), .B(KEYINPUT32), .ZN(n743) );
  NAND2_X1 U830 ( .A1(n744), .A2(n743), .ZN(n767) );
  NOR2_X1 U831 ( .A1(G1976), .A2(G288), .ZN(n749) );
  NOR2_X1 U832 ( .A1(G1971), .A2(G303), .ZN(n745) );
  NOR2_X1 U833 ( .A1(n749), .A2(n745), .ZN(n746) );
  XNOR2_X1 U834 ( .A(KEYINPUT102), .B(n746), .ZN(n747) );
  AND2_X1 U835 ( .A1(n767), .A2(n747), .ZN(n748) );
  NOR2_X1 U836 ( .A1(n748), .A2(n769), .ZN(n755) );
  NAND2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n948) );
  INV_X1 U838 ( .A(KEYINPUT33), .ZN(n757) );
  INV_X1 U839 ( .A(n749), .ZN(n949) );
  OR2_X1 U840 ( .A1(n769), .A2(n949), .ZN(n750) );
  NOR2_X1 U841 ( .A1(n757), .A2(n750), .ZN(n751) );
  XNOR2_X1 U842 ( .A(n751), .B(KEYINPUT103), .ZN(n756) );
  AND2_X1 U843 ( .A1(n948), .A2(n756), .ZN(n753) );
  XNOR2_X1 U844 ( .A(G1981), .B(G305), .ZN(n938) );
  INV_X1 U845 ( .A(n938), .ZN(n752) );
  AND2_X1 U846 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U847 ( .A1(n755), .A2(n754), .ZN(n761) );
  INV_X1 U848 ( .A(n756), .ZN(n758) );
  OR2_X1 U849 ( .A1(n758), .A2(n757), .ZN(n759) );
  OR2_X1 U850 ( .A1(n938), .A2(n759), .ZN(n760) );
  NAND2_X1 U851 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U852 ( .A(n762), .B(KEYINPUT104), .ZN(n763) );
  NOR2_X1 U853 ( .A1(n764), .A2(n763), .ZN(n772) );
  NOR2_X1 U854 ( .A1(G2090), .A2(G303), .ZN(n765) );
  XOR2_X1 U855 ( .A(KEYINPUT105), .B(n765), .Z(n766) );
  NAND2_X1 U856 ( .A1(G8), .A2(n766), .ZN(n768) );
  NAND2_X1 U857 ( .A1(n768), .A2(n767), .ZN(n770) );
  NAND2_X1 U858 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U859 ( .A1(n772), .A2(n771), .ZN(n809) );
  NOR2_X1 U860 ( .A1(n774), .A2(n773), .ZN(n821) );
  XNOR2_X1 U861 ( .A(G1986), .B(G290), .ZN(n942) );
  NAND2_X1 U862 ( .A1(n821), .A2(n942), .ZN(n794) );
  NAND2_X1 U863 ( .A1(G95), .A2(n881), .ZN(n776) );
  NAND2_X1 U864 ( .A1(G107), .A2(n889), .ZN(n775) );
  NAND2_X1 U865 ( .A1(n776), .A2(n775), .ZN(n780) );
  NAND2_X1 U866 ( .A1(G131), .A2(n882), .ZN(n778) );
  NAND2_X1 U867 ( .A1(G119), .A2(n886), .ZN(n777) );
  NAND2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n779) );
  OR2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n864) );
  NAND2_X1 U870 ( .A1(G1991), .A2(n864), .ZN(n791) );
  NAND2_X1 U871 ( .A1(G117), .A2(n889), .ZN(n782) );
  NAND2_X1 U872 ( .A1(G129), .A2(n886), .ZN(n781) );
  NAND2_X1 U873 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U874 ( .A(KEYINPUT90), .B(n783), .ZN(n787) );
  NAND2_X1 U875 ( .A1(G105), .A2(n881), .ZN(n784) );
  XNOR2_X1 U876 ( .A(n784), .B(KEYINPUT91), .ZN(n785) );
  XNOR2_X1 U877 ( .A(n785), .B(KEYINPUT38), .ZN(n786) );
  NOR2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n789) );
  NAND2_X1 U879 ( .A1(n882), .A2(G141), .ZN(n788) );
  NAND2_X1 U880 ( .A1(n789), .A2(n788), .ZN(n863) );
  NAND2_X1 U881 ( .A1(G1996), .A2(n863), .ZN(n790) );
  NAND2_X1 U882 ( .A1(n791), .A2(n790), .ZN(n912) );
  NAND2_X1 U883 ( .A1(n821), .A2(n912), .ZN(n792) );
  XOR2_X1 U884 ( .A(KEYINPUT92), .B(n792), .Z(n813) );
  INV_X1 U885 ( .A(n813), .ZN(n793) );
  NAND2_X1 U886 ( .A1(n794), .A2(n793), .ZN(n807) );
  NAND2_X1 U887 ( .A1(G104), .A2(n881), .ZN(n796) );
  NAND2_X1 U888 ( .A1(G140), .A2(n882), .ZN(n795) );
  NAND2_X1 U889 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U890 ( .A(KEYINPUT34), .B(n797), .ZN(n802) );
  NAND2_X1 U891 ( .A1(G116), .A2(n889), .ZN(n799) );
  NAND2_X1 U892 ( .A1(G128), .A2(n886), .ZN(n798) );
  NAND2_X1 U893 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U894 ( .A(n800), .B(KEYINPUT35), .Z(n801) );
  NOR2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n803) );
  XOR2_X1 U896 ( .A(KEYINPUT36), .B(n803), .Z(n804) );
  XOR2_X1 U897 ( .A(KEYINPUT88), .B(n804), .Z(n867) );
  XNOR2_X1 U898 ( .A(KEYINPUT37), .B(G2067), .ZN(n819) );
  NOR2_X1 U899 ( .A1(n867), .A2(n819), .ZN(n915) );
  NAND2_X1 U900 ( .A1(n915), .A2(n821), .ZN(n805) );
  XOR2_X1 U901 ( .A(KEYINPUT89), .B(n805), .Z(n817) );
  INV_X1 U902 ( .A(n817), .ZN(n806) );
  NOR2_X1 U903 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U905 ( .A(n810), .B(KEYINPUT106), .ZN(n824) );
  NOR2_X1 U906 ( .A1(G1996), .A2(n863), .ZN(n927) );
  NOR2_X1 U907 ( .A1(G1986), .A2(G290), .ZN(n811) );
  NOR2_X1 U908 ( .A1(G1991), .A2(n864), .ZN(n914) );
  NOR2_X1 U909 ( .A1(n811), .A2(n914), .ZN(n812) );
  NOR2_X1 U910 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U911 ( .A1(n927), .A2(n814), .ZN(n815) );
  XOR2_X1 U912 ( .A(n815), .B(KEYINPUT39), .Z(n816) );
  XNOR2_X1 U913 ( .A(KEYINPUT107), .B(n816), .ZN(n818) );
  NAND2_X1 U914 ( .A1(n818), .A2(n817), .ZN(n820) );
  NAND2_X1 U915 ( .A1(n867), .A2(n819), .ZN(n911) );
  NAND2_X1 U916 ( .A1(n820), .A2(n911), .ZN(n822) );
  NAND2_X1 U917 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U918 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U919 ( .A(n825), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n826), .ZN(G217) );
  NAND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n828) );
  INV_X1 U922 ( .A(G661), .ZN(n827) );
  NOR2_X1 U923 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U924 ( .A(n829), .B(KEYINPUT111), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U926 ( .A1(n831), .A2(n830), .ZN(G188) );
  INV_X1 U927 ( .A(n832), .ZN(G319) );
  XNOR2_X1 U928 ( .A(G1991), .B(KEYINPUT41), .ZN(n842) );
  XOR2_X1 U929 ( .A(G1981), .B(G1961), .Z(n834) );
  XNOR2_X1 U930 ( .A(G1996), .B(G1966), .ZN(n833) );
  XNOR2_X1 U931 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U932 ( .A(G1976), .B(G1971), .Z(n836) );
  XNOR2_X1 U933 ( .A(G1986), .B(G1956), .ZN(n835) );
  XNOR2_X1 U934 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U935 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U936 ( .A(KEYINPUT114), .B(G2474), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(G229) );
  XOR2_X1 U939 ( .A(G2100), .B(KEYINPUT113), .Z(n844) );
  XNOR2_X1 U940 ( .A(KEYINPUT112), .B(KEYINPUT43), .ZN(n843) );
  XNOR2_X1 U941 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U942 ( .A(KEYINPUT42), .B(G2090), .Z(n846) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2072), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U945 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U946 ( .A(G2678), .B(G2096), .ZN(n849) );
  XNOR2_X1 U947 ( .A(n850), .B(n849), .ZN(n852) );
  XOR2_X1 U948 ( .A(G2084), .B(G2078), .Z(n851) );
  XNOR2_X1 U949 ( .A(n852), .B(n851), .ZN(G227) );
  NAND2_X1 U950 ( .A1(G124), .A2(n886), .ZN(n853) );
  XOR2_X1 U951 ( .A(KEYINPUT115), .B(n853), .Z(n854) );
  XNOR2_X1 U952 ( .A(n854), .B(KEYINPUT44), .ZN(n856) );
  NAND2_X1 U953 ( .A1(G136), .A2(n882), .ZN(n855) );
  NAND2_X1 U954 ( .A1(n856), .A2(n855), .ZN(n857) );
  XOR2_X1 U955 ( .A(KEYINPUT116), .B(n857), .Z(n859) );
  NAND2_X1 U956 ( .A1(n881), .A2(G100), .ZN(n858) );
  NAND2_X1 U957 ( .A1(n859), .A2(n858), .ZN(n862) );
  NAND2_X1 U958 ( .A1(G112), .A2(n889), .ZN(n860) );
  XNOR2_X1 U959 ( .A(KEYINPUT117), .B(n860), .ZN(n861) );
  NOR2_X1 U960 ( .A1(n862), .A2(n861), .ZN(G162) );
  XNOR2_X1 U961 ( .A(KEYINPUT48), .B(n863), .ZN(n865) );
  XNOR2_X1 U962 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U963 ( .A(n866), .B(KEYINPUT46), .Z(n869) );
  XNOR2_X1 U964 ( .A(n867), .B(G162), .ZN(n868) );
  XNOR2_X1 U965 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U966 ( .A(n870), .B(n919), .Z(n880) );
  NAND2_X1 U967 ( .A1(G103), .A2(n881), .ZN(n872) );
  NAND2_X1 U968 ( .A1(G139), .A2(n882), .ZN(n871) );
  NAND2_X1 U969 ( .A1(n872), .A2(n871), .ZN(n878) );
  NAND2_X1 U970 ( .A1(G115), .A2(n889), .ZN(n874) );
  NAND2_X1 U971 ( .A1(G127), .A2(n886), .ZN(n873) );
  NAND2_X1 U972 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U973 ( .A(KEYINPUT119), .B(n875), .ZN(n876) );
  XNOR2_X1 U974 ( .A(KEYINPUT47), .B(n876), .ZN(n877) );
  NOR2_X1 U975 ( .A1(n878), .A2(n877), .ZN(n922) );
  XNOR2_X1 U976 ( .A(G160), .B(n922), .ZN(n879) );
  XNOR2_X1 U977 ( .A(n880), .B(n879), .ZN(n895) );
  NAND2_X1 U978 ( .A1(G106), .A2(n881), .ZN(n884) );
  NAND2_X1 U979 ( .A1(G142), .A2(n882), .ZN(n883) );
  NAND2_X1 U980 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U981 ( .A(n885), .B(KEYINPUT45), .ZN(n888) );
  NAND2_X1 U982 ( .A1(G130), .A2(n886), .ZN(n887) );
  NAND2_X1 U983 ( .A1(n888), .A2(n887), .ZN(n892) );
  NAND2_X1 U984 ( .A1(n889), .A2(G118), .ZN(n890) );
  XOR2_X1 U985 ( .A(KEYINPUT118), .B(n890), .Z(n891) );
  NOR2_X1 U986 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U987 ( .A(G164), .B(n893), .ZN(n894) );
  XNOR2_X1 U988 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U989 ( .A1(G37), .A2(n896), .ZN(G395) );
  XNOR2_X1 U990 ( .A(G171), .B(n897), .ZN(n898) );
  XNOR2_X1 U991 ( .A(n898), .B(G286), .ZN(n900) );
  XNOR2_X1 U992 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U993 ( .A1(G37), .A2(n901), .ZN(G397) );
  NOR2_X1 U994 ( .A1(G229), .A2(G227), .ZN(n903) );
  XNOR2_X1 U995 ( .A(KEYINPUT49), .B(KEYINPUT120), .ZN(n902) );
  XNOR2_X1 U996 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U997 ( .A1(G401), .A2(n904), .ZN(n905) );
  NAND2_X1 U998 ( .A1(G319), .A2(n905), .ZN(n906) );
  XNOR2_X1 U999 ( .A(KEYINPUT121), .B(n906), .ZN(n908) );
  NOR2_X1 U1000 ( .A1(G395), .A2(G397), .ZN(n907) );
  NAND2_X1 U1001 ( .A1(n908), .A2(n907), .ZN(G225) );
  XOR2_X1 U1002 ( .A(KEYINPUT122), .B(G225), .Z(G308) );
  INV_X1 U1004 ( .A(G120), .ZN(G236) );
  INV_X1 U1005 ( .A(G108), .ZN(G238) );
  INV_X1 U1006 ( .A(G96), .ZN(G221) );
  INV_X1 U1007 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1008 ( .A1(n910), .A2(n909), .ZN(G325) );
  INV_X1 U1009 ( .A(G325), .ZN(G261) );
  INV_X1 U1010 ( .A(G171), .ZN(G301) );
  INV_X1 U1011 ( .A(n911), .ZN(n913) );
  NOR2_X1 U1012 ( .A1(n913), .A2(n912), .ZN(n921) );
  XNOR2_X1 U1013 ( .A(G160), .B(G2084), .ZN(n917) );
  NOR2_X1 U1014 ( .A1(n915), .A2(n914), .ZN(n916) );
  NAND2_X1 U1015 ( .A1(n917), .A2(n916), .ZN(n918) );
  NOR2_X1 U1016 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(n932) );
  XOR2_X1 U1018 ( .A(G2072), .B(n922), .Z(n924) );
  XOR2_X1 U1019 ( .A(G164), .B(G2078), .Z(n923) );
  NOR2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1021 ( .A(KEYINPUT50), .B(n925), .ZN(n930) );
  XOR2_X1 U1022 ( .A(G2090), .B(G162), .Z(n926) );
  NOR2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1024 ( .A(KEYINPUT51), .B(n928), .Z(n929) );
  NAND2_X1 U1025 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1026 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1027 ( .A(KEYINPUT52), .B(n933), .ZN(n935) );
  INV_X1 U1028 ( .A(KEYINPUT55), .ZN(n934) );
  NAND2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1030 ( .A1(n936), .A2(G29), .ZN(n1013) );
  XNOR2_X1 U1031 ( .A(G16), .B(KEYINPUT56), .ZN(n962) );
  XOR2_X1 U1032 ( .A(G1966), .B(G168), .Z(n937) );
  NOR2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1034 ( .A(KEYINPUT57), .B(n939), .Z(n960) );
  XNOR2_X1 U1035 ( .A(G1348), .B(n940), .ZN(n941) );
  NOR2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n947) );
  XNOR2_X1 U1037 ( .A(G301), .B(G1961), .ZN(n945) );
  XNOR2_X1 U1038 ( .A(n943), .B(G1341), .ZN(n944) );
  NOR2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n957) );
  NAND2_X1 U1041 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1042 ( .A(KEYINPUT124), .B(n950), .Z(n954) );
  XNOR2_X1 U1043 ( .A(G299), .B(G1956), .ZN(n952) );
  XNOR2_X1 U1044 ( .A(G303), .B(G1971), .ZN(n951) );
  NOR2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1046 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1047 ( .A(KEYINPUT125), .B(n955), .Z(n956) );
  NOR2_X1 U1048 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1049 ( .A(KEYINPUT126), .B(n958), .ZN(n959) );
  NAND2_X1 U1050 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1051 ( .A1(n962), .A2(n961), .ZN(n988) );
  INV_X1 U1052 ( .A(G16), .ZN(n986) );
  XNOR2_X1 U1053 ( .A(KEYINPUT127), .B(G1341), .ZN(n963) );
  XNOR2_X1 U1054 ( .A(n963), .B(G19), .ZN(n969) );
  XOR2_X1 U1055 ( .A(G1348), .B(KEYINPUT59), .Z(n964) );
  XNOR2_X1 U1056 ( .A(G4), .B(n964), .ZN(n967) );
  XNOR2_X1 U1057 ( .A(G20), .B(n965), .ZN(n966) );
  NOR2_X1 U1058 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1059 ( .A1(n969), .A2(n968), .ZN(n971) );
  XNOR2_X1 U1060 ( .A(G6), .B(G1981), .ZN(n970) );
  NOR2_X1 U1061 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1062 ( .A(KEYINPUT60), .B(n972), .ZN(n976) );
  XNOR2_X1 U1063 ( .A(G1966), .B(G21), .ZN(n974) );
  XNOR2_X1 U1064 ( .A(G5), .B(G1961), .ZN(n973) );
  NOR2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1066 ( .A1(n976), .A2(n975), .ZN(n983) );
  XNOR2_X1 U1067 ( .A(G1971), .B(G22), .ZN(n978) );
  XNOR2_X1 U1068 ( .A(G23), .B(G1976), .ZN(n977) );
  NOR2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n980) );
  XOR2_X1 U1070 ( .A(G1986), .B(G24), .Z(n979) );
  NAND2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(KEYINPUT58), .B(n981), .ZN(n982) );
  NOR2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1074 ( .A(KEYINPUT61), .B(n984), .ZN(n985) );
  NAND2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1076 ( .A1(n988), .A2(n987), .ZN(n1011) );
  XOR2_X1 U1077 ( .A(G1991), .B(G25), .Z(n989) );
  NAND2_X1 U1078 ( .A1(n989), .A2(G28), .ZN(n998) );
  XNOR2_X1 U1079 ( .A(G1996), .B(G32), .ZN(n991) );
  XNOR2_X1 U1080 ( .A(G33), .B(G2072), .ZN(n990) );
  NOR2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n996) );
  XNOR2_X1 U1082 ( .A(G2067), .B(G26), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(G27), .B(n992), .ZN(n993) );
  NOR2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1086 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1087 ( .A(KEYINPUT53), .B(n999), .Z(n1002) );
  XOR2_X1 U1088 ( .A(KEYINPUT54), .B(G34), .Z(n1000) );
  XNOR2_X1 U1089 ( .A(G2084), .B(n1000), .ZN(n1001) );
  NAND2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(G35), .B(G2090), .ZN(n1003) );
  NOR2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(KEYINPUT55), .B(n1005), .ZN(n1007) );
  INV_X1 U1094 ( .A(G29), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1096 ( .A1(n1008), .A2(G11), .ZN(n1009) );
  XOR2_X1 U1097 ( .A(KEYINPUT123), .B(n1009), .Z(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1100 ( .A(KEYINPUT62), .B(n1014), .Z(G311) );
  INV_X1 U1101 ( .A(G311), .ZN(G150) );
endmodule

