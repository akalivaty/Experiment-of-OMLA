

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U551 ( .A1(G651), .A2(n647), .ZN(n659) );
  NAND2_X1 U552 ( .A1(n726), .A2(G1996), .ZN(n711) );
  NOR2_X1 U553 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U554 ( .A(n524), .B(n523), .ZN(n522) );
  INV_X1 U555 ( .A(KEYINPUT99), .ZN(n523) );
  NOR2_X1 U556 ( .A1(G164), .A2(G1384), .ZN(n791) );
  INV_X1 U557 ( .A(G2104), .ZN(n530) );
  AND2_X1 U558 ( .A1(n791), .A2(n700), .ZN(n726) );
  XNOR2_X1 U559 ( .A(n741), .B(n740), .ZN(n742) );
  XNOR2_X1 U560 ( .A(n739), .B(KEYINPUT98), .ZN(n740) );
  INV_X1 U561 ( .A(n726), .ZN(n744) );
  XNOR2_X1 U562 ( .A(n766), .B(KEYINPUT101), .ZN(n532) );
  XNOR2_X1 U563 ( .A(n528), .B(KEYINPUT88), .ZN(n566) );
  AND2_X1 U564 ( .A1(n778), .A2(n518), .ZN(n517) );
  AND2_X1 U565 ( .A1(n566), .A2(n565), .ZN(G164) );
  OR2_X1 U566 ( .A1(n770), .A2(n777), .ZN(n518) );
  NAND2_X1 U567 ( .A1(G303), .A2(n747), .ZN(n519) );
  AND2_X1 U568 ( .A1(n827), .A2(n980), .ZN(n520) );
  NAND2_X1 U569 ( .A1(n521), .A2(G8), .ZN(n748) );
  NAND2_X1 U570 ( .A1(n522), .A2(n519), .ZN(n521) );
  NAND2_X1 U571 ( .A1(n750), .A2(G286), .ZN(n524) );
  XNOR2_X1 U572 ( .A(n525), .B(n829), .ZN(G329) );
  NAND2_X1 U573 ( .A1(n526), .A2(n828), .ZN(n525) );
  XNOR2_X1 U574 ( .A(n814), .B(n527), .ZN(n526) );
  INV_X1 U575 ( .A(KEYINPUT103), .ZN(n527) );
  NAND2_X1 U576 ( .A1(n890), .A2(G138), .ZN(n528) );
  XNOR2_X2 U577 ( .A(n529), .B(KEYINPUT17), .ZN(n890) );
  NAND2_X1 U578 ( .A1(n560), .A2(n530), .ZN(n529) );
  NAND2_X1 U579 ( .A1(n531), .A2(n517), .ZN(n813) );
  NAND2_X1 U580 ( .A1(n532), .A2(n767), .ZN(n531) );
  XNOR2_X1 U581 ( .A(KEYINPUT30), .B(KEYINPUT96), .ZN(n734) );
  XNOR2_X1 U582 ( .A(n735), .B(n734), .ZN(n736) );
  INV_X1 U583 ( .A(KEYINPUT31), .ZN(n739) );
  NAND2_X1 U584 ( .A1(n743), .A2(n742), .ZN(n750) );
  AND2_X1 U585 ( .A1(n698), .A2(n697), .ZN(n700) );
  NAND2_X1 U586 ( .A1(G8), .A2(n744), .ZN(n777) );
  NOR2_X1 U587 ( .A1(n647), .A2(n537), .ZN(n656) );
  AND2_X1 U588 ( .A1(n560), .A2(G2104), .ZN(n891) );
  NOR2_X1 U589 ( .A1(G651), .A2(G543), .ZN(n655) );
  NAND2_X1 U590 ( .A1(n655), .A2(G89), .ZN(n533) );
  XNOR2_X1 U591 ( .A(n533), .B(KEYINPUT4), .ZN(n535) );
  XOR2_X1 U592 ( .A(G543), .B(KEYINPUT0), .Z(n647) );
  INV_X1 U593 ( .A(G651), .ZN(n537) );
  NAND2_X1 U594 ( .A1(G76), .A2(n656), .ZN(n534) );
  NAND2_X1 U595 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U596 ( .A(KEYINPUT5), .B(n536), .ZN(n546) );
  XNOR2_X1 U597 ( .A(KEYINPUT73), .B(KEYINPUT74), .ZN(n544) );
  NAND2_X1 U598 ( .A1(G51), .A2(n659), .ZN(n541) );
  NOR2_X1 U599 ( .A1(G543), .A2(n537), .ZN(n539) );
  XNOR2_X1 U600 ( .A(KEYINPUT1), .B(KEYINPUT65), .ZN(n538) );
  XNOR2_X1 U601 ( .A(n539), .B(n538), .ZN(n653) );
  NAND2_X1 U602 ( .A1(G63), .A2(n653), .ZN(n540) );
  NAND2_X1 U603 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U604 ( .A(n542), .B(KEYINPUT6), .ZN(n543) );
  XNOR2_X1 U605 ( .A(n544), .B(n543), .ZN(n545) );
  NAND2_X1 U606 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U607 ( .A(KEYINPUT7), .B(n547), .ZN(G168) );
  XOR2_X1 U608 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U609 ( .A1(G91), .A2(n655), .ZN(n549) );
  NAND2_X1 U610 ( .A1(G78), .A2(n656), .ZN(n548) );
  NAND2_X1 U611 ( .A1(n549), .A2(n548), .ZN(n553) );
  NAND2_X1 U612 ( .A1(G53), .A2(n659), .ZN(n551) );
  NAND2_X1 U613 ( .A1(G65), .A2(n653), .ZN(n550) );
  NAND2_X1 U614 ( .A1(n551), .A2(n550), .ZN(n552) );
  OR2_X1 U615 ( .A1(n553), .A2(n552), .ZN(G299) );
  INV_X1 U616 ( .A(KEYINPUT23), .ZN(n555) );
  INV_X1 U617 ( .A(G2105), .ZN(n560) );
  NAND2_X1 U618 ( .A1(G101), .A2(n891), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n555), .B(n554), .ZN(n695) );
  INV_X1 U620 ( .A(KEYINPUT64), .ZN(n559) );
  NAND2_X1 U621 ( .A1(n890), .A2(G137), .ZN(n557) );
  AND2_X1 U622 ( .A1(G2105), .A2(G2104), .ZN(n887) );
  NAND2_X1 U623 ( .A1(n887), .A2(G113), .ZN(n556) );
  NAND2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n697) );
  NOR2_X1 U626 ( .A1(G2104), .A2(n560), .ZN(n620) );
  NAND2_X1 U627 ( .A1(n620), .A2(G125), .ZN(n696) );
  AND2_X1 U628 ( .A1(n697), .A2(n696), .ZN(n789) );
  AND2_X1 U629 ( .A1(n695), .A2(n789), .ZN(G160) );
  AND2_X1 U630 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U631 ( .A(G57), .ZN(G237) );
  INV_X1 U632 ( .A(G132), .ZN(G219) );
  INV_X1 U633 ( .A(G82), .ZN(G220) );
  NAND2_X1 U634 ( .A1(G114), .A2(n887), .ZN(n562) );
  NAND2_X1 U635 ( .A1(G102), .A2(n891), .ZN(n561) );
  NAND2_X1 U636 ( .A1(n562), .A2(n561), .ZN(n564) );
  AND2_X1 U637 ( .A1(G126), .A2(n620), .ZN(n563) );
  NOR2_X1 U638 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U639 ( .A1(G90), .A2(n655), .ZN(n568) );
  NAND2_X1 U640 ( .A1(G77), .A2(n656), .ZN(n567) );
  NAND2_X1 U641 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U642 ( .A(KEYINPUT9), .B(n569), .ZN(n573) );
  NAND2_X1 U643 ( .A1(n659), .A2(G52), .ZN(n571) );
  NAND2_X1 U644 ( .A1(G64), .A2(n653), .ZN(n570) );
  AND2_X1 U645 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U646 ( .A1(n573), .A2(n572), .ZN(G301) );
  NAND2_X1 U647 ( .A1(G50), .A2(n659), .ZN(n575) );
  NAND2_X1 U648 ( .A1(G62), .A2(n653), .ZN(n574) );
  NAND2_X1 U649 ( .A1(n575), .A2(n574), .ZN(n579) );
  NAND2_X1 U650 ( .A1(G88), .A2(n655), .ZN(n577) );
  NAND2_X1 U651 ( .A1(G75), .A2(n656), .ZN(n576) );
  NAND2_X1 U652 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U653 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U654 ( .A(n580), .B(KEYINPUT83), .ZN(G303) );
  NAND2_X1 U655 ( .A1(G7), .A2(G661), .ZN(n581) );
  XNOR2_X1 U656 ( .A(n581), .B(KEYINPUT68), .ZN(n582) );
  XNOR2_X1 U657 ( .A(KEYINPUT10), .B(n582), .ZN(G223) );
  INV_X1 U658 ( .A(G223), .ZN(n830) );
  NAND2_X1 U659 ( .A1(n830), .A2(G567), .ZN(n583) );
  XOR2_X1 U660 ( .A(KEYINPUT11), .B(n583), .Z(G234) );
  XNOR2_X1 U661 ( .A(KEYINPUT13), .B(KEYINPUT69), .ZN(n588) );
  NAND2_X1 U662 ( .A1(n655), .A2(G81), .ZN(n584) );
  XNOR2_X1 U663 ( .A(n584), .B(KEYINPUT12), .ZN(n586) );
  NAND2_X1 U664 ( .A1(G68), .A2(n656), .ZN(n585) );
  NAND2_X1 U665 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U666 ( .A(n588), .B(n587), .ZN(n591) );
  NAND2_X1 U667 ( .A1(n653), .A2(G56), .ZN(n589) );
  XOR2_X1 U668 ( .A(KEYINPUT14), .B(n589), .Z(n590) );
  NOR2_X1 U669 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U670 ( .A(n592), .B(KEYINPUT70), .ZN(n594) );
  NAND2_X1 U671 ( .A1(G43), .A2(n659), .ZN(n593) );
  NAND2_X1 U672 ( .A1(n594), .A2(n593), .ZN(n992) );
  INV_X1 U673 ( .A(G860), .ZN(n609) );
  OR2_X1 U674 ( .A1(n992), .A2(n609), .ZN(G153) );
  NAND2_X1 U675 ( .A1(n653), .A2(G66), .ZN(n601) );
  NAND2_X1 U676 ( .A1(G54), .A2(n659), .ZN(n595) );
  XNOR2_X1 U677 ( .A(KEYINPUT71), .B(n595), .ZN(n599) );
  NAND2_X1 U678 ( .A1(G79), .A2(n656), .ZN(n597) );
  NAND2_X1 U679 ( .A1(G92), .A2(n655), .ZN(n596) );
  NAND2_X1 U680 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U681 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U682 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U683 ( .A(KEYINPUT15), .B(n602), .Z(n981) );
  NOR2_X1 U684 ( .A1(G868), .A2(n981), .ZN(n604) );
  INV_X1 U685 ( .A(G868), .ZN(n677) );
  NOR2_X1 U686 ( .A1(n677), .A2(G301), .ZN(n603) );
  NOR2_X1 U687 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U688 ( .A(KEYINPUT72), .B(n605), .ZN(G284) );
  XNOR2_X1 U689 ( .A(KEYINPUT75), .B(G868), .ZN(n606) );
  NOR2_X1 U690 ( .A1(G286), .A2(n606), .ZN(n608) );
  NOR2_X1 U691 ( .A1(G868), .A2(G299), .ZN(n607) );
  NOR2_X1 U692 ( .A1(n608), .A2(n607), .ZN(G297) );
  NAND2_X1 U693 ( .A1(n609), .A2(G559), .ZN(n610) );
  INV_X1 U694 ( .A(n981), .ZN(n636) );
  NAND2_X1 U695 ( .A1(n610), .A2(n636), .ZN(n611) );
  XNOR2_X1 U696 ( .A(n611), .B(KEYINPUT16), .ZN(n612) );
  XNOR2_X1 U697 ( .A(KEYINPUT76), .B(n612), .ZN(G148) );
  NOR2_X1 U698 ( .A1(n981), .A2(n677), .ZN(n613) );
  XNOR2_X1 U699 ( .A(n613), .B(KEYINPUT77), .ZN(n614) );
  NOR2_X1 U700 ( .A1(G559), .A2(n614), .ZN(n615) );
  XNOR2_X1 U701 ( .A(n615), .B(KEYINPUT78), .ZN(n617) );
  NOR2_X1 U702 ( .A1(n992), .A2(G868), .ZN(n616) );
  NOR2_X1 U703 ( .A1(n617), .A2(n616), .ZN(G282) );
  NAND2_X1 U704 ( .A1(G111), .A2(n887), .ZN(n619) );
  NAND2_X1 U705 ( .A1(G135), .A2(n890), .ZN(n618) );
  NAND2_X1 U706 ( .A1(n619), .A2(n618), .ZN(n623) );
  NAND2_X1 U707 ( .A1(n620), .A2(G123), .ZN(n621) );
  XOR2_X1 U708 ( .A(KEYINPUT18), .B(n621), .Z(n622) );
  NOR2_X1 U709 ( .A1(n623), .A2(n622), .ZN(n625) );
  NAND2_X1 U710 ( .A1(n891), .A2(G99), .ZN(n624) );
  NAND2_X1 U711 ( .A1(n625), .A2(n624), .ZN(n954) );
  XNOR2_X1 U712 ( .A(G2096), .B(n954), .ZN(n626) );
  NOR2_X1 U713 ( .A1(n626), .A2(G2100), .ZN(n627) );
  XNOR2_X1 U714 ( .A(n627), .B(KEYINPUT79), .ZN(G156) );
  NAND2_X1 U715 ( .A1(G93), .A2(n655), .ZN(n629) );
  NAND2_X1 U716 ( .A1(G80), .A2(n656), .ZN(n628) );
  NAND2_X1 U717 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U718 ( .A(n630), .B(KEYINPUT81), .ZN(n632) );
  NAND2_X1 U719 ( .A1(G67), .A2(n653), .ZN(n631) );
  NAND2_X1 U720 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U721 ( .A1(n659), .A2(G55), .ZN(n633) );
  XOR2_X1 U722 ( .A(KEYINPUT82), .B(n633), .Z(n634) );
  OR2_X1 U723 ( .A1(n635), .A2(n634), .ZN(n676) );
  XNOR2_X1 U724 ( .A(KEYINPUT80), .B(n992), .ZN(n637) );
  NAND2_X1 U725 ( .A1(n636), .A2(G559), .ZN(n674) );
  XNOR2_X1 U726 ( .A(n637), .B(n674), .ZN(n638) );
  NOR2_X1 U727 ( .A1(G860), .A2(n638), .ZN(n639) );
  XOR2_X1 U728 ( .A(n676), .B(n639), .Z(G145) );
  NAND2_X1 U729 ( .A1(G86), .A2(n655), .ZN(n641) );
  NAND2_X1 U730 ( .A1(G61), .A2(n653), .ZN(n640) );
  NAND2_X1 U731 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U732 ( .A1(n656), .A2(G73), .ZN(n642) );
  XOR2_X1 U733 ( .A(KEYINPUT2), .B(n642), .Z(n643) );
  NOR2_X1 U734 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U735 ( .A1(n659), .A2(G48), .ZN(n645) );
  NAND2_X1 U736 ( .A1(n646), .A2(n645), .ZN(G305) );
  NAND2_X1 U737 ( .A1(G49), .A2(n659), .ZN(n649) );
  NAND2_X1 U738 ( .A1(G87), .A2(n647), .ZN(n648) );
  NAND2_X1 U739 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U740 ( .A1(n653), .A2(n650), .ZN(n652) );
  NAND2_X1 U741 ( .A1(G651), .A2(G74), .ZN(n651) );
  NAND2_X1 U742 ( .A1(n652), .A2(n651), .ZN(G288) );
  NAND2_X1 U743 ( .A1(n653), .A2(G60), .ZN(n654) );
  XNOR2_X1 U744 ( .A(n654), .B(KEYINPUT66), .ZN(n664) );
  NAND2_X1 U745 ( .A1(G85), .A2(n655), .ZN(n658) );
  NAND2_X1 U746 ( .A1(G72), .A2(n656), .ZN(n657) );
  NAND2_X1 U747 ( .A1(n658), .A2(n657), .ZN(n662) );
  NAND2_X1 U748 ( .A1(G47), .A2(n659), .ZN(n660) );
  XNOR2_X1 U749 ( .A(KEYINPUT67), .B(n660), .ZN(n661) );
  NOR2_X1 U750 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U751 ( .A1(n664), .A2(n663), .ZN(G290) );
  INV_X1 U752 ( .A(G303), .ZN(G166) );
  XOR2_X1 U753 ( .A(KEYINPUT85), .B(KEYINPUT19), .Z(n665) );
  XNOR2_X1 U754 ( .A(G288), .B(n665), .ZN(n666) );
  XNOR2_X1 U755 ( .A(KEYINPUT84), .B(n666), .ZN(n668) );
  XNOR2_X1 U756 ( .A(G290), .B(KEYINPUT86), .ZN(n667) );
  XNOR2_X1 U757 ( .A(n668), .B(n667), .ZN(n669) );
  XOR2_X1 U758 ( .A(n676), .B(n669), .Z(n671) );
  XNOR2_X1 U759 ( .A(n992), .B(G166), .ZN(n670) );
  XNOR2_X1 U760 ( .A(n671), .B(n670), .ZN(n672) );
  XOR2_X1 U761 ( .A(n672), .B(G299), .Z(n673) );
  XNOR2_X1 U762 ( .A(G305), .B(n673), .ZN(n904) );
  XNOR2_X1 U763 ( .A(n674), .B(n904), .ZN(n675) );
  NAND2_X1 U764 ( .A1(n675), .A2(G868), .ZN(n679) );
  NAND2_X1 U765 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U766 ( .A1(n679), .A2(n678), .ZN(G295) );
  NAND2_X1 U767 ( .A1(G2084), .A2(G2078), .ZN(n680) );
  XOR2_X1 U768 ( .A(KEYINPUT20), .B(n680), .Z(n681) );
  NAND2_X1 U769 ( .A1(G2090), .A2(n681), .ZN(n682) );
  XNOR2_X1 U770 ( .A(KEYINPUT21), .B(n682), .ZN(n683) );
  NAND2_X1 U771 ( .A1(n683), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U772 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U773 ( .A1(G220), .A2(G219), .ZN(n684) );
  XOR2_X1 U774 ( .A(KEYINPUT22), .B(n684), .Z(n685) );
  NOR2_X1 U775 ( .A1(G218), .A2(n685), .ZN(n686) );
  XOR2_X1 U776 ( .A(KEYINPUT87), .B(n686), .Z(n687) );
  NAND2_X1 U777 ( .A1(G96), .A2(n687), .ZN(n834) );
  NAND2_X1 U778 ( .A1(n834), .A2(G2106), .ZN(n691) );
  NAND2_X1 U779 ( .A1(G108), .A2(G120), .ZN(n688) );
  NOR2_X1 U780 ( .A1(G237), .A2(n688), .ZN(n689) );
  NAND2_X1 U781 ( .A1(G69), .A2(n689), .ZN(n835) );
  NAND2_X1 U782 ( .A1(n835), .A2(G567), .ZN(n690) );
  NAND2_X1 U783 ( .A1(n691), .A2(n690), .ZN(n858) );
  NAND2_X1 U784 ( .A1(G483), .A2(G661), .ZN(n692) );
  NOR2_X1 U785 ( .A1(n858), .A2(n692), .ZN(n833) );
  NAND2_X1 U786 ( .A1(n833), .A2(G36), .ZN(G176) );
  XOR2_X1 U787 ( .A(G1981), .B(KEYINPUT102), .Z(n693) );
  XNOR2_X1 U788 ( .A(G305), .B(n693), .ZN(n986) );
  NOR2_X1 U789 ( .A1(G1976), .A2(G288), .ZN(n694) );
  XOR2_X1 U790 ( .A(KEYINPUT100), .B(n694), .Z(n758) );
  AND2_X1 U791 ( .A1(n695), .A2(G40), .ZN(n788) );
  AND2_X1 U792 ( .A1(n788), .A2(n696), .ZN(n698) );
  NOR2_X1 U793 ( .A1(n758), .A2(n777), .ZN(n701) );
  NAND2_X1 U794 ( .A1(KEYINPUT33), .A2(n701), .ZN(n702) );
  AND2_X1 U795 ( .A1(n986), .A2(n702), .ZN(n767) );
  NAND2_X1 U796 ( .A1(G1348), .A2(n744), .ZN(n704) );
  NAND2_X1 U797 ( .A1(G2067), .A2(n726), .ZN(n703) );
  NAND2_X1 U798 ( .A1(n704), .A2(n703), .ZN(n710) );
  NOR2_X1 U799 ( .A1(n981), .A2(n710), .ZN(n709) );
  NAND2_X1 U800 ( .A1(n726), .A2(G2072), .ZN(n705) );
  XOR2_X1 U801 ( .A(KEYINPUT27), .B(n705), .Z(n707) );
  NAND2_X1 U802 ( .A1(G1956), .A2(n744), .ZN(n706) );
  NAND2_X1 U803 ( .A1(n707), .A2(n706), .ZN(n721) );
  NOR2_X1 U804 ( .A1(n721), .A2(G299), .ZN(n708) );
  NOR2_X1 U805 ( .A1(n709), .A2(n708), .ZN(n719) );
  NAND2_X1 U806 ( .A1(n710), .A2(n981), .ZN(n717) );
  XNOR2_X1 U807 ( .A(n711), .B(KEYINPUT26), .ZN(n713) );
  NAND2_X1 U808 ( .A1(G1341), .A2(n744), .ZN(n712) );
  NAND2_X1 U809 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U810 ( .A(KEYINPUT94), .B(n714), .ZN(n715) );
  NOR2_X1 U811 ( .A1(n992), .A2(n715), .ZN(n716) );
  NAND2_X1 U812 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U813 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U814 ( .A(n720), .B(KEYINPUT95), .ZN(n724) );
  NAND2_X1 U815 ( .A1(G299), .A2(n721), .ZN(n722) );
  XOR2_X1 U816 ( .A(KEYINPUT28), .B(n722), .Z(n723) );
  XNOR2_X1 U817 ( .A(n725), .B(KEYINPUT29), .ZN(n730) );
  NAND2_X1 U818 ( .A1(G1961), .A2(n744), .ZN(n728) );
  XOR2_X1 U819 ( .A(G2078), .B(KEYINPUT25), .Z(n934) );
  NAND2_X1 U820 ( .A1(n726), .A2(n934), .ZN(n727) );
  NAND2_X1 U821 ( .A1(n728), .A2(n727), .ZN(n731) );
  OR2_X1 U822 ( .A1(n731), .A2(G301), .ZN(n729) );
  NAND2_X1 U823 ( .A1(n730), .A2(n729), .ZN(n743) );
  NAND2_X1 U824 ( .A1(G301), .A2(n731), .ZN(n732) );
  XNOR2_X1 U825 ( .A(n732), .B(KEYINPUT97), .ZN(n738) );
  NOR2_X1 U826 ( .A1(G1966), .A2(n777), .ZN(n752) );
  NOR2_X1 U827 ( .A1(G2084), .A2(n744), .ZN(n749) );
  NOR2_X1 U828 ( .A1(n752), .A2(n749), .ZN(n733) );
  NAND2_X1 U829 ( .A1(G8), .A2(n733), .ZN(n735) );
  NOR2_X1 U830 ( .A1(n736), .A2(G168), .ZN(n737) );
  NOR2_X1 U831 ( .A1(n738), .A2(n737), .ZN(n741) );
  NOR2_X1 U832 ( .A1(G1971), .A2(n777), .ZN(n746) );
  NOR2_X1 U833 ( .A1(G2090), .A2(n744), .ZN(n745) );
  NOR2_X1 U834 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U835 ( .A(KEYINPUT32), .B(n748), .ZN(n771) );
  NAND2_X1 U836 ( .A1(G8), .A2(n749), .ZN(n754) );
  INV_X1 U837 ( .A(n750), .ZN(n751) );
  NOR2_X1 U838 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U839 ( .A1(n754), .A2(n753), .ZN(n772) );
  NAND2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n974) );
  INV_X1 U841 ( .A(n974), .ZN(n755) );
  OR2_X1 U842 ( .A1(n777), .A2(n755), .ZN(n761) );
  INV_X1 U843 ( .A(n761), .ZN(n756) );
  AND2_X1 U844 ( .A1(n772), .A2(n756), .ZN(n757) );
  AND2_X1 U845 ( .A1(n771), .A2(n757), .ZN(n765) );
  NOR2_X1 U846 ( .A1(G1971), .A2(G303), .ZN(n760) );
  INV_X1 U847 ( .A(n758), .ZN(n759) );
  NOR2_X1 U848 ( .A1(n760), .A2(n759), .ZN(n983) );
  OR2_X1 U849 ( .A1(n761), .A2(n983), .ZN(n763) );
  INV_X1 U850 ( .A(KEYINPUT33), .ZN(n762) );
  NAND2_X1 U851 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U852 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U853 ( .A1(G1981), .A2(G305), .ZN(n768) );
  XNOR2_X1 U854 ( .A(n768), .B(KEYINPUT24), .ZN(n769) );
  XNOR2_X1 U855 ( .A(n769), .B(KEYINPUT93), .ZN(n770) );
  NAND2_X1 U856 ( .A1(n772), .A2(n771), .ZN(n775) );
  NOR2_X1 U857 ( .A1(G2090), .A2(G303), .ZN(n773) );
  NAND2_X1 U858 ( .A1(G8), .A2(n773), .ZN(n774) );
  NAND2_X1 U859 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U860 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U861 ( .A1(G140), .A2(n890), .ZN(n780) );
  NAND2_X1 U862 ( .A1(G104), .A2(n891), .ZN(n779) );
  NAND2_X1 U863 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U864 ( .A(KEYINPUT34), .B(n781), .ZN(n786) );
  NAND2_X1 U865 ( .A1(G116), .A2(n887), .ZN(n783) );
  NAND2_X1 U866 ( .A1(G128), .A2(n620), .ZN(n782) );
  NAND2_X1 U867 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U868 ( .A(KEYINPUT35), .B(n784), .Z(n785) );
  NOR2_X1 U869 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U870 ( .A(KEYINPUT36), .B(n787), .ZN(n901) );
  XNOR2_X1 U871 ( .A(KEYINPUT37), .B(G2067), .ZN(n824) );
  NOR2_X1 U872 ( .A1(n901), .A2(n824), .ZN(n947) );
  NAND2_X1 U873 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U874 ( .A1(n791), .A2(n790), .ZN(n827) );
  NAND2_X1 U875 ( .A1(n947), .A2(n827), .ZN(n792) );
  XNOR2_X1 U876 ( .A(n792), .B(KEYINPUT89), .ZN(n821) );
  NAND2_X1 U877 ( .A1(G107), .A2(n887), .ZN(n794) );
  NAND2_X1 U878 ( .A1(G131), .A2(n890), .ZN(n793) );
  NAND2_X1 U879 ( .A1(n794), .A2(n793), .ZN(n798) );
  NAND2_X1 U880 ( .A1(G95), .A2(n891), .ZN(n796) );
  NAND2_X1 U881 ( .A1(G119), .A2(n620), .ZN(n795) );
  NAND2_X1 U882 ( .A1(n796), .A2(n795), .ZN(n797) );
  NOR2_X1 U883 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U884 ( .A(KEYINPUT90), .B(n799), .Z(n881) );
  NAND2_X1 U885 ( .A1(n881), .A2(G1991), .ZN(n808) );
  NAND2_X1 U886 ( .A1(G117), .A2(n887), .ZN(n801) );
  NAND2_X1 U887 ( .A1(G141), .A2(n890), .ZN(n800) );
  NAND2_X1 U888 ( .A1(n801), .A2(n800), .ZN(n804) );
  NAND2_X1 U889 ( .A1(n891), .A2(G105), .ZN(n802) );
  XOR2_X1 U890 ( .A(KEYINPUT38), .B(n802), .Z(n803) );
  NOR2_X1 U891 ( .A1(n804), .A2(n803), .ZN(n806) );
  NAND2_X1 U892 ( .A1(n620), .A2(G129), .ZN(n805) );
  NAND2_X1 U893 ( .A1(n806), .A2(n805), .ZN(n880) );
  NAND2_X1 U894 ( .A1(G1996), .A2(n880), .ZN(n807) );
  NAND2_X1 U895 ( .A1(n808), .A2(n807), .ZN(n957) );
  NAND2_X1 U896 ( .A1(n957), .A2(n827), .ZN(n809) );
  XNOR2_X1 U897 ( .A(n809), .B(KEYINPUT91), .ZN(n818) );
  NOR2_X1 U898 ( .A1(n821), .A2(n818), .ZN(n810) );
  XOR2_X1 U899 ( .A(KEYINPUT92), .B(n810), .Z(n811) );
  XNOR2_X1 U900 ( .A(G1986), .B(G290), .ZN(n980) );
  NOR2_X1 U901 ( .A1(n811), .A2(n520), .ZN(n812) );
  NAND2_X1 U902 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U903 ( .A1(G1996), .A2(n880), .ZN(n950) );
  NOR2_X1 U904 ( .A1(n881), .A2(G1991), .ZN(n953) );
  NOR2_X1 U905 ( .A1(G1986), .A2(G290), .ZN(n815) );
  XNOR2_X1 U906 ( .A(KEYINPUT104), .B(n815), .ZN(n816) );
  NOR2_X1 U907 ( .A1(n953), .A2(n816), .ZN(n817) );
  NOR2_X1 U908 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U909 ( .A1(n950), .A2(n819), .ZN(n820) );
  XNOR2_X1 U910 ( .A(n820), .B(KEYINPUT39), .ZN(n823) );
  INV_X1 U911 ( .A(n821), .ZN(n822) );
  NAND2_X1 U912 ( .A1(n823), .A2(n822), .ZN(n825) );
  NAND2_X1 U913 ( .A1(n901), .A2(n824), .ZN(n946) );
  NAND2_X1 U914 ( .A1(n825), .A2(n946), .ZN(n826) );
  NAND2_X1 U915 ( .A1(n827), .A2(n826), .ZN(n828) );
  XOR2_X1 U916 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n829) );
  INV_X1 U917 ( .A(G301), .ZN(G171) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n830), .ZN(G217) );
  AND2_X1 U919 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U920 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U921 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U922 ( .A1(n833), .A2(n832), .ZN(G188) );
  XNOR2_X1 U923 ( .A(G120), .B(KEYINPUT107), .ZN(G236) );
  INV_X1 U925 ( .A(G108), .ZN(G238) );
  INV_X1 U926 ( .A(G96), .ZN(G221) );
  NOR2_X1 U927 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U928 ( .A(G325), .ZN(G261) );
  XOR2_X1 U929 ( .A(KEYINPUT43), .B(G2678), .Z(n837) );
  XNOR2_X1 U930 ( .A(KEYINPUT109), .B(KEYINPUT108), .ZN(n836) );
  XNOR2_X1 U931 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U932 ( .A(KEYINPUT42), .B(G2090), .Z(n839) );
  XNOR2_X1 U933 ( .A(G2067), .B(G2072), .ZN(n838) );
  XNOR2_X1 U934 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U935 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U936 ( .A(G2096), .B(G2100), .ZN(n842) );
  XNOR2_X1 U937 ( .A(n843), .B(n842), .ZN(n845) );
  XOR2_X1 U938 ( .A(G2084), .B(G2078), .Z(n844) );
  XNOR2_X1 U939 ( .A(n845), .B(n844), .ZN(G227) );
  XOR2_X1 U940 ( .A(G1981), .B(G1956), .Z(n847) );
  XNOR2_X1 U941 ( .A(G1966), .B(G1961), .ZN(n846) );
  XNOR2_X1 U942 ( .A(n847), .B(n846), .ZN(n857) );
  XOR2_X1 U943 ( .A(G2474), .B(KEYINPUT41), .Z(n849) );
  XNOR2_X1 U944 ( .A(G1991), .B(KEYINPUT111), .ZN(n848) );
  XNOR2_X1 U945 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U946 ( .A(G1976), .B(G1971), .Z(n851) );
  XNOR2_X1 U947 ( .A(G1996), .B(G1986), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U949 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U950 ( .A(KEYINPUT112), .B(KEYINPUT110), .ZN(n854) );
  XNOR2_X1 U951 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U952 ( .A(n857), .B(n856), .ZN(G229) );
  INV_X1 U953 ( .A(n858), .ZN(G319) );
  NAND2_X1 U954 ( .A1(G100), .A2(n891), .ZN(n859) );
  XNOR2_X1 U955 ( .A(n859), .B(KEYINPUT114), .ZN(n863) );
  XOR2_X1 U956 ( .A(KEYINPUT113), .B(KEYINPUT44), .Z(n861) );
  NAND2_X1 U957 ( .A1(G124), .A2(n620), .ZN(n860) );
  XNOR2_X1 U958 ( .A(n861), .B(n860), .ZN(n862) );
  NAND2_X1 U959 ( .A1(n863), .A2(n862), .ZN(n867) );
  NAND2_X1 U960 ( .A1(G112), .A2(n887), .ZN(n865) );
  NAND2_X1 U961 ( .A1(G136), .A2(n890), .ZN(n864) );
  NAND2_X1 U962 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U963 ( .A1(n867), .A2(n866), .ZN(G162) );
  XOR2_X1 U964 ( .A(KEYINPUT48), .B(KEYINPUT118), .Z(n869) );
  XNOR2_X1 U965 ( .A(KEYINPUT119), .B(KEYINPUT46), .ZN(n868) );
  XNOR2_X1 U966 ( .A(n869), .B(n868), .ZN(n886) );
  NAND2_X1 U967 ( .A1(G139), .A2(n890), .ZN(n871) );
  NAND2_X1 U968 ( .A1(G103), .A2(n891), .ZN(n870) );
  NAND2_X1 U969 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U970 ( .A(KEYINPUT116), .B(n872), .ZN(n878) );
  NAND2_X1 U971 ( .A1(G115), .A2(n887), .ZN(n874) );
  NAND2_X1 U972 ( .A1(G127), .A2(n620), .ZN(n873) );
  NAND2_X1 U973 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U974 ( .A(KEYINPUT47), .B(n875), .ZN(n876) );
  XNOR2_X1 U975 ( .A(KEYINPUT117), .B(n876), .ZN(n877) );
  NOR2_X1 U976 ( .A1(n878), .A2(n877), .ZN(n960) );
  XOR2_X1 U977 ( .A(n960), .B(G162), .Z(n879) );
  XNOR2_X1 U978 ( .A(n880), .B(n879), .ZN(n882) );
  XOR2_X1 U979 ( .A(n882), .B(n881), .Z(n884) );
  XNOR2_X1 U980 ( .A(G160), .B(G164), .ZN(n883) );
  XNOR2_X1 U981 ( .A(n884), .B(n883), .ZN(n885) );
  XNOR2_X1 U982 ( .A(n886), .B(n885), .ZN(n900) );
  NAND2_X1 U983 ( .A1(G118), .A2(n887), .ZN(n889) );
  NAND2_X1 U984 ( .A1(G130), .A2(n620), .ZN(n888) );
  NAND2_X1 U985 ( .A1(n889), .A2(n888), .ZN(n897) );
  NAND2_X1 U986 ( .A1(G142), .A2(n890), .ZN(n893) );
  NAND2_X1 U987 ( .A1(G106), .A2(n891), .ZN(n892) );
  NAND2_X1 U988 ( .A1(n893), .A2(n892), .ZN(n894) );
  XNOR2_X1 U989 ( .A(KEYINPUT115), .B(n894), .ZN(n895) );
  XNOR2_X1 U990 ( .A(KEYINPUT45), .B(n895), .ZN(n896) );
  NOR2_X1 U991 ( .A1(n897), .A2(n896), .ZN(n898) );
  XNOR2_X1 U992 ( .A(n954), .B(n898), .ZN(n899) );
  XNOR2_X1 U993 ( .A(n900), .B(n899), .ZN(n902) );
  XOR2_X1 U994 ( .A(n902), .B(n901), .Z(n903) );
  NOR2_X1 U995 ( .A1(G37), .A2(n903), .ZN(G395) );
  XNOR2_X1 U996 ( .A(G286), .B(n981), .ZN(n905) );
  XNOR2_X1 U997 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U998 ( .A(n906), .B(G171), .ZN(n907) );
  NOR2_X1 U999 ( .A1(G37), .A2(n907), .ZN(G397) );
  NOR2_X1 U1000 ( .A1(G227), .A2(G229), .ZN(n909) );
  XNOR2_X1 U1001 ( .A(KEYINPUT49), .B(KEYINPUT120), .ZN(n908) );
  XNOR2_X1 U1002 ( .A(n909), .B(n908), .ZN(n921) );
  XOR2_X1 U1003 ( .A(G2443), .B(G2451), .Z(n911) );
  XNOR2_X1 U1004 ( .A(G2446), .B(G2454), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1006 ( .A(n912), .B(G2427), .Z(n914) );
  XNOR2_X1 U1007 ( .A(G1348), .B(G1341), .ZN(n913) );
  XNOR2_X1 U1008 ( .A(n914), .B(n913), .ZN(n918) );
  XOR2_X1 U1009 ( .A(G2435), .B(KEYINPUT106), .Z(n916) );
  XNOR2_X1 U1010 ( .A(G2430), .B(G2438), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(n916), .B(n915), .ZN(n917) );
  XOR2_X1 U1012 ( .A(n918), .B(n917), .Z(n919) );
  NAND2_X1 U1013 ( .A1(G14), .A2(n919), .ZN(n924) );
  NAND2_X1 U1014 ( .A1(G319), .A2(n924), .ZN(n920) );
  NOR2_X1 U1015 ( .A1(n921), .A2(n920), .ZN(n923) );
  NOR2_X1 U1016 ( .A1(G395), .A2(G397), .ZN(n922) );
  NAND2_X1 U1017 ( .A1(n923), .A2(n922), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(G69), .ZN(G235) );
  INV_X1 U1020 ( .A(n924), .ZN(G401) );
  XNOR2_X1 U1021 ( .A(G2084), .B(G34), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(n925), .B(KEYINPUT54), .ZN(n942) );
  XNOR2_X1 U1023 ( .A(G2090), .B(G35), .ZN(n939) );
  XNOR2_X1 U1024 ( .A(G1996), .B(G32), .ZN(n927) );
  XNOR2_X1 U1025 ( .A(G33), .B(G2072), .ZN(n926) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n933) );
  XOR2_X1 U1027 ( .A(G2067), .B(G26), .Z(n928) );
  NAND2_X1 U1028 ( .A1(n928), .A2(G28), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(G25), .B(G1991), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(KEYINPUT122), .B(n929), .ZN(n930) );
  NOR2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n936) );
  XNOR2_X1 U1033 ( .A(G27), .B(n934), .ZN(n935) );
  NOR2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1035 ( .A(KEYINPUT53), .B(n937), .ZN(n938) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1037 ( .A(n940), .B(KEYINPUT123), .ZN(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1039 ( .A(KEYINPUT124), .B(n943), .ZN(n944) );
  NOR2_X1 U1040 ( .A1(G29), .A2(n944), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(n945), .B(KEYINPUT55), .ZN(n972) );
  INV_X1 U1042 ( .A(n946), .ZN(n948) );
  NOR2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n968) );
  XOR2_X1 U1044 ( .A(G2090), .B(G162), .Z(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1046 ( .A(KEYINPUT51), .B(n951), .Z(n959) );
  XOR2_X1 U1047 ( .A(G160), .B(G2084), .Z(n952) );
  NOR2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n955) );
  NAND2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(n966) );
  XNOR2_X1 U1052 ( .A(G2072), .B(n960), .ZN(n962) );
  XNOR2_X1 U1053 ( .A(G164), .B(G2078), .ZN(n961) );
  NAND2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1055 ( .A(KEYINPUT121), .B(n963), .Z(n964) );
  XNOR2_X1 U1056 ( .A(KEYINPUT50), .B(n964), .ZN(n965) );
  NOR2_X1 U1057 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1058 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1059 ( .A(KEYINPUT52), .B(n969), .ZN(n970) );
  NAND2_X1 U1060 ( .A1(G29), .A2(n970), .ZN(n971) );
  NAND2_X1 U1061 ( .A1(n972), .A2(n971), .ZN(n1023) );
  XOR2_X1 U1062 ( .A(G1956), .B(G299), .Z(n973) );
  NAND2_X1 U1063 ( .A1(n974), .A2(n973), .ZN(n976) );
  XNOR2_X1 U1064 ( .A(G1961), .B(G301), .ZN(n975) );
  NOR2_X1 U1065 ( .A1(n976), .A2(n975), .ZN(n978) );
  NAND2_X1 U1066 ( .A1(G1971), .A2(G303), .ZN(n977) );
  NAND2_X1 U1067 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1068 ( .A1(n980), .A2(n979), .ZN(n991) );
  XOR2_X1 U1069 ( .A(G1348), .B(n981), .Z(n982) );
  NAND2_X1 U1070 ( .A1(n983), .A2(n982), .ZN(n989) );
  XOR2_X1 U1071 ( .A(G1966), .B(G168), .Z(n984) );
  XNOR2_X1 U1072 ( .A(KEYINPUT125), .B(n984), .ZN(n985) );
  NAND2_X1 U1073 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1074 ( .A(KEYINPUT57), .B(n987), .Z(n988) );
  NOR2_X1 U1075 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1076 ( .A1(n991), .A2(n990), .ZN(n994) );
  XNOR2_X1 U1077 ( .A(G1341), .B(n992), .ZN(n993) );
  NOR2_X1 U1078 ( .A1(n994), .A2(n993), .ZN(n996) );
  XOR2_X1 U1079 ( .A(G16), .B(KEYINPUT56), .Z(n995) );
  NOR2_X1 U1080 ( .A1(n996), .A2(n995), .ZN(n1020) );
  XNOR2_X1 U1081 ( .A(G1971), .B(G22), .ZN(n998) );
  XNOR2_X1 U1082 ( .A(G23), .B(G1976), .ZN(n997) );
  NOR2_X1 U1083 ( .A1(n998), .A2(n997), .ZN(n1000) );
  XOR2_X1 U1084 ( .A(G1986), .B(G24), .Z(n999) );
  NAND2_X1 U1085 ( .A1(n1000), .A2(n999), .ZN(n1002) );
  XOR2_X1 U1086 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n1001) );
  XNOR2_X1 U1087 ( .A(n1002), .B(n1001), .ZN(n1006) );
  XNOR2_X1 U1088 ( .A(G1966), .B(G21), .ZN(n1004) );
  XNOR2_X1 U1089 ( .A(G5), .B(G1961), .ZN(n1003) );
  NOR2_X1 U1090 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1091 ( .A1(n1006), .A2(n1005), .ZN(n1016) );
  XOR2_X1 U1092 ( .A(G1348), .B(KEYINPUT59), .Z(n1007) );
  XNOR2_X1 U1093 ( .A(G4), .B(n1007), .ZN(n1009) );
  XNOR2_X1 U1094 ( .A(G20), .B(G1956), .ZN(n1008) );
  NOR2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1013) );
  XNOR2_X1 U1096 ( .A(G1341), .B(G19), .ZN(n1011) );
  XNOR2_X1 U1097 ( .A(G6), .B(G1981), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(KEYINPUT60), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1102 ( .A(KEYINPUT61), .B(n1017), .Z(n1018) );
  NOR2_X1 U1103 ( .A1(G16), .A2(n1018), .ZN(n1019) );
  NOR2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1105 ( .A(KEYINPUT127), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1106 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1107 ( .A1(n1024), .A2(G11), .ZN(n1025) );
  XOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1025), .Z(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

