//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 1 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 1 0 1 0 1 1 1 0 1 1 0 1 0 1 0 0 1 1 1 1 1 0 1 0 1 0 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(new_n188), .B(KEYINPUT78), .Z(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT1), .B1(new_n190), .B2(G146), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(G146), .ZN(new_n194));
  AOI22_X1  g008(.A1(new_n191), .A2(G128), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(KEYINPUT1), .ZN(new_n197));
  AND3_X1   g011(.A1(new_n197), .A2(new_n193), .A3(new_n194), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT10), .B1(new_n195), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G104), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT3), .B1(new_n200), .B2(G107), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n202));
  INV_X1    g016(.A(G107), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(G104), .ZN(new_n204));
  INV_X1    g018(.A(G101), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n200), .A2(G107), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n201), .A2(new_n204), .A3(new_n205), .A4(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n200), .A2(G107), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n203), .A2(G104), .ZN(new_n209));
  OAI21_X1  g023(.A(G101), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT81), .B1(new_n199), .B2(new_n211), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n207), .A2(new_n210), .ZN(new_n213));
  XNOR2_X1  g027(.A(G143), .B(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n197), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n196), .B1(new_n193), .B2(KEYINPUT1), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n215), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT81), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n213), .A2(new_n217), .A3(new_n218), .A4(KEYINPUT10), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n212), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT1), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n221), .B1(G143), .B2(new_n192), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT80), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n196), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n191), .A2(KEYINPUT80), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n214), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n213), .B1(new_n226), .B2(new_n198), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT10), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT11), .ZN(new_n230));
  INV_X1    g044(.A(G134), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(G137), .ZN(new_n232));
  INV_X1    g046(.A(G137), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(KEYINPUT11), .A3(G134), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n231), .A2(G137), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n232), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G131), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(KEYINPUT65), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n238), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n240), .A2(new_n232), .A3(new_n234), .A4(new_n235), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n201), .A2(new_n204), .A3(new_n206), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G101), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(KEYINPUT4), .A3(new_n207), .ZN(new_n246));
  AND2_X1   g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n193), .A2(new_n194), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT0), .B(G128), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n248), .B(KEYINPUT64), .C1(new_n214), .C2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n193), .A2(new_n194), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT64), .ZN(new_n252));
  INV_X1    g066(.A(new_n247), .ZN(new_n253));
  OR2_X1    g067(.A1(KEYINPUT0), .A2(G128), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n251), .A2(new_n252), .A3(new_n253), .A4(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n244), .A2(new_n257), .A3(G101), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n246), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n220), .A2(new_n229), .A3(new_n243), .A4(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(KEYINPUT82), .B1(new_n213), .B2(new_n217), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n195), .A2(new_n198), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT82), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(new_n263), .A3(new_n211), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n227), .A2(new_n261), .A3(new_n264), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n265), .A2(KEYINPUT12), .A3(new_n242), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT12), .B1(new_n265), .B2(new_n242), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n260), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(G110), .B(G140), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n269), .B(KEYINPUT79), .ZN(new_n270));
  INV_X1    g084(.A(G227), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n271), .A2(G953), .ZN(new_n272));
  XOR2_X1   g086(.A(new_n270), .B(new_n272), .Z(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n260), .A2(new_n273), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n220), .A2(new_n229), .A3(new_n259), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n242), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n268), .A2(new_n274), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(G469), .B1(new_n279), .B2(G902), .ZN(new_n280));
  INV_X1    g094(.A(G902), .ZN(new_n281));
  XNOR2_X1  g095(.A(KEYINPUT83), .B(G469), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n266), .A2(new_n267), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(new_n275), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n273), .B1(new_n278), .B2(new_n260), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n281), .B(new_n282), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n189), .B1(new_n280), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G475), .ZN(new_n288));
  XNOR2_X1  g102(.A(G113), .B(G122), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n289), .B(new_n200), .ZN(new_n290));
  INV_X1    g104(.A(G140), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(G125), .ZN(new_n292));
  INV_X1    g106(.A(G125), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G140), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT74), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n292), .A2(new_n294), .A3(new_n295), .A4(KEYINPUT16), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n292), .A2(new_n294), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT16), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n291), .A3(G125), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT74), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n192), .B(new_n296), .C1(new_n299), .C2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  OAI211_X1 g117(.A(KEYINPUT74), .B(new_n300), .C1(new_n297), .C2(new_n298), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n192), .B1(new_n304), .B2(new_n296), .ZN(new_n305));
  NOR2_X1   g119(.A1(G237), .A2(G953), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n306), .A2(G143), .A3(G214), .ZN(new_n307));
  AOI21_X1  g121(.A(G143), .B1(new_n306), .B2(G214), .ZN(new_n308));
  OAI21_X1  g122(.A(G131), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT17), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NOR3_X1   g125(.A1(new_n303), .A2(new_n305), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G237), .ZN(new_n313));
  INV_X1    g127(.A(G953), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n314), .A3(G214), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n190), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n306), .A2(G143), .A3(G214), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT89), .B1(new_n318), .B2(G131), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT89), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n316), .A2(new_n320), .A3(new_n237), .A4(new_n317), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n319), .A2(new_n310), .A3(new_n309), .A4(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT92), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n309), .A2(new_n321), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n325), .A2(KEYINPUT92), .A3(new_n310), .A4(new_n319), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n312), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(KEYINPUT18), .A2(G131), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n318), .B(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n293), .A2(G140), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n291), .A2(G125), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT88), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT88), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n292), .A2(new_n294), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n333), .A2(G146), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n292), .A2(new_n294), .A3(new_n192), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n330), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n290), .B1(new_n327), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT93), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n327), .A2(new_n290), .A3(new_n340), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(G902), .B1(new_n341), .B2(KEYINPUT93), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n288), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n344), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT90), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n292), .A2(new_n294), .A3(new_n334), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n334), .B1(new_n292), .B2(new_n294), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT19), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT19), .B1(new_n292), .B2(new_n294), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n349), .B1(new_n355), .B2(new_n192), .ZN(new_n356));
  AOI211_X1 g170(.A(KEYINPUT90), .B(G146), .C1(new_n352), .C2(new_n354), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n305), .B1(new_n325), .B2(new_n319), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n339), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT91), .B1(new_n360), .B2(new_n290), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n333), .A2(new_n335), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n353), .B1(new_n362), .B2(KEYINPUT19), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT90), .B1(new_n363), .B2(G146), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n355), .A2(new_n349), .A3(new_n192), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n359), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n340), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT91), .ZN(new_n368));
  INV_X1    g182(.A(new_n290), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n348), .B1(new_n361), .B2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(G475), .A2(G902), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT20), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n368), .B1(new_n367), .B2(new_n369), .ZN(new_n375));
  AOI211_X1 g189(.A(KEYINPUT91), .B(new_n290), .C1(new_n366), .C2(new_n340), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n344), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT20), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(new_n372), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n347), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT14), .ZN(new_n381));
  INV_X1    g195(.A(G116), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n381), .B1(new_n382), .B2(G122), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT96), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(G122), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G122), .ZN(new_n387));
  AOI21_X1  g201(.A(KEYINPUT14), .B1(new_n387), .B2(G116), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n387), .A2(G116), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT96), .B1(new_n385), .B2(KEYINPUT14), .ZN(new_n391));
  OAI211_X1 g205(.A(G107), .B(new_n386), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n382), .A2(G122), .ZN(new_n393));
  OR3_X1    g207(.A1(new_n389), .A2(new_n393), .A3(G107), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT94), .B1(new_n196), .B2(G143), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT94), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(new_n190), .A3(G128), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n196), .A2(G143), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n398), .A2(new_n231), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n231), .B1(new_n398), .B2(new_n399), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n392), .B(new_n394), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT97), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n398), .A2(new_n399), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G134), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n398), .A2(new_n231), .A3(new_n399), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n408), .A2(KEYINPUT97), .A3(new_n392), .A4(new_n394), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT13), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n398), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n399), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n398), .A2(new_n411), .ZN(new_n414));
  OAI21_X1  g228(.A(G134), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT95), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n398), .A2(new_n416), .A3(new_n231), .A4(new_n399), .ZN(new_n417));
  OAI21_X1  g231(.A(G107), .B1(new_n389), .B2(new_n393), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n394), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n407), .A2(KEYINPUT95), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n415), .A2(new_n417), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G217), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n187), .A2(new_n422), .A3(G953), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n410), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n423), .B1(new_n410), .B2(new_n421), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n281), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT98), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G478), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(KEYINPUT15), .ZN(new_n430));
  OAI211_X1 g244(.A(KEYINPUT98), .B(new_n281), .C1(new_n424), .C2(new_n425), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  OR2_X1    g246(.A1(new_n426), .A2(new_n430), .ZN(new_n433));
  AOI211_X1 g247(.A(new_n281), .B(new_n314), .C1(G234), .C2(G237), .ZN(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(G898), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n314), .A2(G952), .ZN(new_n437));
  INV_X1    g251(.A(G234), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n437), .B1(new_n438), .B2(new_n313), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n432), .A2(new_n433), .A3(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G214), .B1(G237), .B2(G902), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(G210), .B1(G237), .B2(G902), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n250), .A2(G125), .A3(new_n255), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n215), .B(new_n293), .C1(new_n214), .C2(new_n216), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT85), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT85), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT87), .ZN(new_n452));
  INV_X1    g266(.A(G224), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n452), .B1(new_n453), .B2(G953), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n314), .A2(KEYINPUT87), .A3(G224), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g270(.A(new_n456), .B(KEYINPUT86), .Z(new_n457));
  NAND3_X1  g271(.A1(new_n449), .A2(new_n451), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n457), .ZN(new_n459));
  INV_X1    g273(.A(new_n451), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n450), .B1(new_n446), .B2(new_n447), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(KEYINPUT2), .B(G113), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(G116), .B(G119), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n466), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n464), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n246), .A2(new_n470), .A3(new_n258), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n466), .A2(KEYINPUT5), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT84), .ZN(new_n473));
  INV_X1    g287(.A(G119), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(G116), .ZN(new_n475));
  OR2_X1    g289(.A1(new_n475), .A2(KEYINPUT5), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n472), .A2(new_n473), .A3(new_n476), .A4(G113), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n382), .A2(G119), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n475), .A2(new_n478), .A3(KEYINPUT5), .ZN(new_n479));
  OAI21_X1  g293(.A(G113), .B1(new_n475), .B2(KEYINPUT5), .ZN(new_n480));
  OAI21_X1  g294(.A(KEYINPUT84), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n213), .A2(new_n477), .A3(new_n481), .A4(new_n467), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n471), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(G110), .B(G122), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n471), .A2(new_n482), .A3(new_n484), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(KEYINPUT6), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT6), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n483), .A2(new_n489), .A3(new_n485), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n463), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT8), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n484), .B(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n467), .B1(new_n479), .B2(new_n480), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n493), .B1(new_n494), .B2(new_n213), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n477), .A2(new_n481), .A3(new_n467), .A4(new_n211), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n454), .A2(KEYINPUT7), .A3(new_n455), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n495), .A2(new_n496), .B1(new_n448), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n449), .A2(new_n451), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n487), .B(new_n498), .C1(new_n499), .C2(new_n497), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n281), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n445), .B1(new_n491), .B2(new_n501), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n500), .A2(new_n281), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n463), .A2(new_n488), .A3(new_n490), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(new_n444), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n443), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  AND4_X1   g320(.A1(new_n287), .A2(new_n380), .A3(new_n441), .A4(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT77), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT22), .B(G137), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n314), .A2(G221), .A3(G234), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n509), .B(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n196), .A2(G119), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n474), .A2(G128), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT24), .B(G110), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n474), .A2(G128), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n517), .B(new_n513), .C1(new_n518), .C2(KEYINPUT23), .ZN(new_n519));
  OR2_X1    g333(.A1(new_n519), .A2(KEYINPUT73), .ZN(new_n520));
  INV_X1    g334(.A(G110), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n521), .B1(new_n519), .B2(KEYINPUT73), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n516), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n303), .B2(new_n305), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n514), .A2(new_n515), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n525), .B1(new_n519), .B2(G110), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n304), .A2(new_n296), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n526), .B(new_n337), .C1(new_n527), .C2(new_n192), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT75), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT75), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n524), .A2(new_n528), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n511), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n529), .A2(new_n511), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n422), .B1(G234), .B2(new_n281), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(G902), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n508), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n536), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(KEYINPUT77), .A3(new_n538), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT76), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT25), .ZN(new_n544));
  AOI21_X1  g358(.A(G902), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n533), .B2(new_n535), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n543), .A2(new_n544), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n537), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n546), .A2(new_n547), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n540), .B(new_n542), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n232), .A2(new_n234), .A3(new_n237), .A4(new_n235), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n231), .A2(G137), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n233), .A2(G134), .ZN(new_n555));
  OAI21_X1  g369(.A(G131), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n262), .A2(new_n557), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n558), .A2(KEYINPUT66), .B1(new_n242), .B2(new_n256), .ZN(new_n559));
  INV_X1    g373(.A(new_n470), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT66), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n561), .B1(new_n262), .B2(new_n557), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n559), .A2(KEYINPUT67), .A3(new_n560), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n256), .A2(new_n242), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n217), .A2(KEYINPUT66), .A3(new_n553), .A4(new_n556), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n564), .A2(new_n562), .A3(new_n565), .A4(new_n560), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT67), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n564), .A2(new_n562), .A3(new_n565), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n470), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT69), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n570), .A2(KEYINPUT69), .A3(new_n470), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n569), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT28), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT28), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n217), .A2(new_n553), .A3(new_n556), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n564), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n577), .B1(new_n579), .B2(new_n470), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT70), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g396(.A(KEYINPUT70), .B(new_n577), .C1(new_n579), .C2(new_n470), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(KEYINPUT26), .B(G101), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n306), .A2(G210), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT29), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n576), .A2(new_n585), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n580), .A2(new_n591), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n563), .A2(new_n568), .B1(new_n470), .B2(new_n579), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n596), .B1(new_n597), .B2(new_n577), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n563), .A2(new_n568), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n570), .A2(KEYINPUT30), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT30), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n564), .A2(new_n601), .A3(new_n578), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n560), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n590), .B1(new_n599), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT29), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n598), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n594), .A2(new_n606), .A3(new_n281), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n607), .A2(KEYINPUT71), .A3(G472), .ZN(new_n608));
  AOI21_X1  g422(.A(KEYINPUT71), .B1(new_n607), .B2(G472), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT32), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n564), .A2(new_n601), .A3(new_n578), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(KEYINPUT30), .B2(new_n570), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n569), .B(new_n591), .C1(new_n613), .C2(new_n560), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT31), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n600), .A2(new_n602), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n617), .A2(new_n470), .B1(new_n563), .B2(new_n568), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n618), .A2(KEYINPUT31), .A3(new_n591), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n580), .B1(new_n597), .B2(new_n577), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n616), .A2(new_n619), .B1(new_n620), .B2(new_n590), .ZN(new_n621));
  INV_X1    g435(.A(G472), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n281), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n611), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT72), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n623), .A2(new_n611), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n625), .B1(new_n621), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n620), .A2(new_n590), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n614), .A2(new_n615), .ZN(new_n630));
  AOI21_X1  g444(.A(KEYINPUT31), .B1(new_n618), .B2(new_n591), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n632), .A2(KEYINPUT72), .A3(new_n626), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n624), .A2(new_n628), .A3(new_n633), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n507), .B(new_n552), .C1(new_n610), .C2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G101), .ZN(G3));
  NAND2_X1  g450(.A1(new_n280), .A2(new_n286), .ZN(new_n637));
  INV_X1    g451(.A(new_n189), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n551), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n622), .B1(new_n632), .B2(new_n281), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n621), .A2(new_n623), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n506), .A2(new_n440), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n640), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n348), .A2(new_n341), .A3(KEYINPUT93), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n341), .A2(KEYINPUT93), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n281), .ZN(new_n649));
  OAI21_X1  g463(.A(G475), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n377), .A2(new_n378), .A3(new_n372), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n378), .B1(new_n377), .B2(new_n372), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT33), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n654), .B1(new_n424), .B2(new_n425), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n429), .A2(G902), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n410), .A2(new_n421), .A3(new_n423), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT100), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n654), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n659), .B1(new_n658), .B2(new_n657), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n425), .B(KEYINPUT99), .ZN(new_n661));
  OAI211_X1 g475(.A(new_n655), .B(new_n656), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n428), .A2(new_n429), .A3(new_n431), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n653), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n646), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT34), .B(G104), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT101), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n666), .B(new_n668), .ZN(G6));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n670), .B1(new_n651), .B2(new_n652), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n374), .A2(KEYINPUT102), .A3(new_n379), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n347), .B1(new_n432), .B2(new_n433), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n646), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT35), .B(G107), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G9));
  NAND2_X1  g491(.A1(new_n530), .A2(new_n532), .ZN(new_n678));
  INV_X1    g492(.A(new_n511), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n679), .A2(KEYINPUT36), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n678), .B(new_n680), .ZN(new_n681));
  OAI22_X1  g495(.A1(new_n549), .A2(new_n550), .B1(new_n539), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n287), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n380), .A2(new_n441), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n684), .A2(new_n685), .A3(new_n506), .A4(new_n643), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT37), .B(G110), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G12));
  AND3_X1   g502(.A1(new_n624), .A2(new_n628), .A3(new_n633), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n605), .B1(new_n618), .B2(new_n591), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n579), .A2(new_n470), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n566), .A2(new_n567), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n566), .A2(new_n567), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n595), .B1(new_n694), .B2(KEYINPUT28), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n281), .B1(new_n690), .B2(new_n695), .ZN(new_n696));
  AOI211_X1 g510(.A(new_n592), .B(new_n584), .C1(new_n575), .C2(KEYINPUT28), .ZN(new_n697));
  OAI21_X1  g511(.A(G472), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT71), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n607), .A2(KEYINPUT71), .A3(G472), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n689), .A2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n439), .ZN(new_n704));
  INV_X1    g518(.A(G900), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n704), .B1(new_n434), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n674), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n703), .A2(new_n506), .A3(new_n684), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G128), .ZN(G30));
  XNOR2_X1  g523(.A(new_n706), .B(KEYINPUT39), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n639), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT40), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n281), .B1(new_n575), .B2(new_n591), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n618), .A2(new_n590), .ZN(new_n714));
  OAI21_X1  g528(.A(G472), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n624), .A2(new_n628), .A3(new_n633), .A4(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n432), .A2(new_n433), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n653), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n502), .A2(new_n505), .ZN(new_n719));
  XOR2_X1   g533(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NOR4_X1   g535(.A1(new_n718), .A2(new_n721), .A3(new_n443), .A4(new_n682), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n712), .A2(new_n716), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G143), .ZN(G45));
  INV_X1    g538(.A(new_n706), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n653), .A2(new_n664), .A3(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n703), .A2(new_n506), .A3(new_n684), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G146), .ZN(G48));
  OAI21_X1  g543(.A(new_n276), .B1(new_n266), .B2(new_n267), .ZN(new_n730));
  INV_X1    g544(.A(new_n285), .ZN(new_n731));
  AOI21_X1  g545(.A(G902), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(G469), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n286), .B(new_n188), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n665), .A2(new_n644), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n703), .A2(new_n552), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(KEYINPUT41), .B(G113), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G15));
  NOR2_X1   g553(.A1(new_n674), .A2(new_n644), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n703), .A2(new_n552), .A3(new_n735), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G116), .ZN(G18));
  NAND2_X1  g556(.A1(new_n719), .A2(new_n442), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n734), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n744), .A2(new_n380), .A3(new_n441), .A4(new_n682), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n745), .B1(new_n702), .B2(new_n689), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n474), .ZN(G21));
  NAND2_X1  g561(.A1(new_n576), .A2(new_n585), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n590), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n616), .A2(new_n619), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n623), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n551), .A2(new_n641), .A3(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n440), .A3(new_n735), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT104), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n743), .B1(new_n718), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n653), .A2(KEYINPUT104), .A3(new_n717), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(KEYINPUT105), .A3(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n717), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n754), .B1(new_n380), .B2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n756), .A3(new_n506), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT105), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n753), .B1(new_n757), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n387), .ZN(G24));
  NOR2_X1   g578(.A1(new_n641), .A2(new_n751), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n682), .ZN(new_n766));
  INV_X1    g580(.A(new_n744), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n766), .A2(new_n726), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(new_n293), .ZN(G27));
  NAND3_X1  g583(.A1(new_n502), .A2(new_n505), .A3(new_n442), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT106), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n502), .A2(new_n505), .A3(KEYINPUT106), .A4(new_n442), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n772), .A2(new_n637), .A3(new_n188), .A4(new_n773), .ZN(new_n774));
  AOI211_X1 g588(.A(new_n551), .B(new_n774), .C1(new_n689), .C2(new_n702), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n726), .A2(KEYINPUT42), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n726), .A2(new_n774), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT107), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n624), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n632), .A2(new_n626), .ZN(new_n780));
  OAI211_X1 g594(.A(KEYINPUT107), .B(new_n611), .C1(new_n621), .C2(new_n623), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n777), .B(new_n552), .C1(new_n610), .C2(new_n782), .ZN(new_n783));
  AOI22_X1  g597(.A1(new_n775), .A2(new_n776), .B1(new_n783), .B2(KEYINPUT42), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G131), .ZN(G33));
  INV_X1    g599(.A(new_n774), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n703), .A2(new_n552), .A3(new_n707), .A4(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G134), .ZN(G36));
  NAND2_X1  g602(.A1(new_n380), .A2(new_n664), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT43), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n789), .B(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT108), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n682), .B1(new_n641), .B2(new_n642), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OR3_X1    g608(.A1(new_n794), .A2(KEYINPUT109), .A3(KEYINPUT44), .ZN(new_n795));
  OAI21_X1  g609(.A(KEYINPUT109), .B1(new_n794), .B2(KEYINPUT44), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n279), .A2(KEYINPUT45), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n279), .A2(KEYINPUT45), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n797), .A2(G469), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(G469), .A2(G902), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT46), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n286), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n799), .A2(KEYINPUT46), .A3(new_n800), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n188), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n805), .A2(new_n710), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n772), .A2(new_n773), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n794), .B2(KEYINPUT44), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n795), .A2(new_n796), .A3(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(KEYINPUT110), .B(G137), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n811), .B(new_n812), .ZN(G39));
  XNOR2_X1  g627(.A(new_n805), .B(KEYINPUT47), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NOR4_X1   g629(.A1(new_n703), .A2(new_n552), .A3(new_n726), .A4(new_n807), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G140), .ZN(G42));
  INV_X1    g632(.A(new_n732), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n802), .B1(G469), .B2(new_n819), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n820), .B(KEYINPUT49), .Z(new_n821));
  NOR4_X1   g635(.A1(new_n821), .A2(new_n551), .A3(new_n189), .A4(new_n443), .ZN(new_n822));
  INV_X1    g636(.A(new_n716), .ZN(new_n823));
  INV_X1    g637(.A(new_n789), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n822), .A2(new_n823), .A3(new_n721), .A4(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n807), .A2(new_n734), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n823), .A2(new_n552), .A3(new_n704), .A4(new_n826), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n827), .A2(new_n653), .A3(new_n664), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n791), .A2(new_n704), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n826), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n766), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n829), .A2(new_n752), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n721), .A2(new_n443), .A3(new_n735), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT50), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n835), .A2(KEYINPUT114), .ZN(new_n836));
  AOI211_X1 g650(.A(new_n828), .B(new_n831), .C1(new_n834), .C2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n835), .A2(KEYINPUT114), .ZN(new_n838));
  OR2_X1    g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n837), .B1(new_n834), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n820), .A2(new_n189), .ZN(new_n841));
  AOI211_X1 g655(.A(new_n807), .B(new_n832), .C1(new_n814), .C2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  OR2_X1    g657(.A1(new_n843), .A2(KEYINPUT51), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(KEYINPUT51), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n552), .B1(new_n782), .B2(new_n610), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n830), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT48), .ZN(new_n848));
  OAI221_X1 g662(.A(new_n437), .B1(new_n665), .B2(new_n827), .C1(new_n832), .C2(new_n767), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n844), .A2(new_n845), .A3(new_n850), .ZN(new_n851));
  AOI211_X1 g665(.A(new_n743), .B(new_n683), .C1(new_n689), .C2(new_n702), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n768), .B1(new_n852), .B2(new_n707), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT52), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n637), .A2(new_n188), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n855), .A2(new_n682), .A3(new_n706), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n716), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT105), .B1(new_n755), .B2(new_n756), .ZN(new_n859));
  AND4_X1   g673(.A1(KEYINPUT105), .A2(new_n759), .A3(new_n756), .A4(new_n506), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n853), .A2(new_n854), .A3(new_n861), .A4(new_n728), .ZN(new_n862));
  INV_X1    g676(.A(new_n766), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n863), .A2(new_n727), .A3(new_n744), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n708), .A2(new_n728), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n857), .B1(new_n757), .B2(new_n762), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT52), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n650), .A2(new_n433), .A3(new_n432), .A4(new_n725), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n869), .A2(new_n672), .A3(new_n671), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT111), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT111), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n869), .A2(new_n872), .A3(new_n671), .A4(new_n672), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n871), .A2(new_n808), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT112), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n683), .B1(new_n689), .B2(new_n702), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT112), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n871), .A2(new_n877), .A3(new_n808), .A4(new_n873), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n875), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n863), .A2(new_n727), .A3(new_n786), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n787), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n784), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  AOI211_X1 g696(.A(new_n551), .B(new_n734), .C1(new_n689), .C2(new_n702), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n746), .B1(new_n883), .B2(new_n736), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n380), .A2(new_n717), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n665), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n886), .A2(new_n640), .A3(new_n643), .A4(new_n645), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n635), .A2(new_n686), .A3(new_n887), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n752), .A2(new_n440), .A3(new_n735), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n889), .B1(new_n859), .B2(new_n860), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n884), .A2(new_n888), .A3(new_n890), .A4(new_n741), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n882), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT53), .B1(new_n868), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n783), .A2(KEYINPUT42), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n703), .A2(new_n552), .A3(new_n786), .A4(new_n776), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n894), .A2(new_n895), .A3(new_n787), .A4(new_n880), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n703), .A2(new_n685), .A3(new_n682), .A4(new_n744), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n737), .A2(new_n741), .A3(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n899), .A2(new_n763), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n897), .A2(new_n900), .A3(new_n888), .A4(new_n879), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n862), .A2(new_n867), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT53), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n904), .B1(new_n853), .B2(new_n854), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n893), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT113), .B1(new_n899), .B2(new_n763), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT113), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n884), .A2(new_n910), .A3(new_n890), .A4(new_n741), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n878), .A2(new_n876), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n807), .B1(new_n870), .B2(KEYINPUT111), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n877), .B1(new_n914), .B2(new_n873), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n896), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n635), .A2(new_n686), .A3(new_n887), .A4(KEYINPUT53), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n708), .A2(new_n864), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n918), .B1(KEYINPUT52), .B2(new_n919), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n912), .A2(new_n868), .A3(new_n917), .A4(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n904), .B1(new_n901), .B2(new_n902), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n921), .A2(new_n922), .A3(new_n907), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n851), .A2(new_n908), .A3(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(G952), .A2(G953), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n825), .B1(new_n925), .B2(new_n926), .ZN(G75));
  INV_X1    g741(.A(KEYINPUT56), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n921), .A2(new_n922), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(G902), .ZN(new_n930));
  INV_X1    g744(.A(G210), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n488), .A2(new_n490), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(new_n463), .ZN(new_n934));
  XNOR2_X1  g748(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n934), .B(new_n935), .Z(new_n936));
  XNOR2_X1  g750(.A(new_n932), .B(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n314), .A2(G952), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT116), .Z(new_n939));
  AND2_X1   g753(.A1(new_n937), .A2(new_n939), .ZN(G51));
  INV_X1    g754(.A(KEYINPUT120), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n917), .A2(new_n920), .A3(new_n909), .A4(new_n911), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n942), .A2(new_n902), .ZN(new_n943));
  OAI21_X1  g757(.A(KEYINPUT54), .B1(new_n943), .B2(new_n893), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n944), .A2(KEYINPUT118), .A3(new_n923), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT118), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n929), .A2(new_n946), .A3(KEYINPUT54), .ZN(new_n947));
  XNOR2_X1  g761(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(new_n800), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n945), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT119), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n945), .A2(KEYINPUT119), .A3(new_n947), .A4(new_n949), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n284), .A2(new_n285), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n941), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n930), .A2(new_n799), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n955), .B1(new_n952), .B2(new_n953), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n957), .B1(new_n958), .B2(KEYINPUT120), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n938), .B1(new_n956), .B2(new_n959), .ZN(G54));
  INV_X1    g774(.A(KEYINPUT58), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n930), .A2(new_n961), .A3(new_n288), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n962), .A2(new_n377), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n962), .A2(new_n377), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n963), .A2(new_n964), .A3(new_n938), .ZN(G60));
  NAND2_X1  g779(.A1(G478), .A2(G902), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT59), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n908), .B2(new_n924), .ZN(new_n968));
  OR2_X1    g782(.A1(new_n660), .A2(new_n661), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n655), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n968), .A2(KEYINPUT121), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(KEYINPUT121), .B1(new_n968), .B2(new_n970), .ZN(new_n972));
  INV_X1    g786(.A(new_n970), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n945), .A2(new_n973), .A3(new_n947), .A4(new_n967), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n939), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n971), .A2(new_n972), .A3(new_n975), .ZN(G63));
  NAND2_X1  g790(.A1(G217), .A2(G902), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT60), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(new_n921), .B2(new_n922), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n939), .B1(new_n979), .B2(new_n541), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n681), .B(KEYINPUT122), .Z(new_n981));
  AOI21_X1  g795(.A(new_n980), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT61), .ZN(G66));
  OAI21_X1  g797(.A(G953), .B1(new_n435), .B2(new_n453), .ZN(new_n984));
  INV_X1    g798(.A(new_n891), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n984), .B1(new_n985), .B2(G953), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n933), .B1(G898), .B2(new_n314), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n986), .B(new_n987), .ZN(G69));
  INV_X1    g802(.A(new_n817), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n989), .A2(new_n865), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n846), .B1(new_n757), .B2(new_n762), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n806), .A2(new_n991), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n990), .A2(new_n784), .A3(new_n787), .A4(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n811), .A2(new_n314), .ZN(new_n994));
  OAI22_X1  g808(.A1(new_n993), .A2(new_n994), .B1(new_n271), .B2(new_n314), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n363), .B(KEYINPUT123), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n617), .B(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(G900), .B1(new_n997), .B2(G227), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(G953), .ZN(new_n1000));
  NOR3_X1   g814(.A1(new_n807), .A2(new_n639), .A3(new_n710), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n703), .A2(new_n552), .A3(new_n886), .A4(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n811), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(KEYINPUT124), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT124), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n811), .A2(new_n1005), .A3(new_n1002), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n853), .A2(new_n723), .A3(new_n728), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(KEYINPUT62), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n989), .A2(new_n1009), .ZN(new_n1010));
  AND2_X1   g824(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  OR2_X1    g825(.A1(new_n997), .A2(G953), .ZN(new_n1012));
  OAI211_X1 g826(.A(new_n998), .B(new_n1000), .C1(new_n1011), .C2(new_n1012), .ZN(G72));
  XOR2_X1   g827(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n1014));
  NOR2_X1   g828(.A1(new_n622), .A2(new_n281), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n811), .A2(new_n985), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1017), .B1(new_n993), .B2(new_n1018), .ZN(new_n1019));
  NOR3_X1   g833(.A1(new_n599), .A2(new_n603), .A3(new_n591), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n938), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1016), .B1(new_n604), .B2(new_n614), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1022), .B(KEYINPUT127), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1021), .B1(new_n906), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1007), .A2(new_n985), .A3(new_n1010), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1025), .A2(new_n1017), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1026), .A2(new_n714), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1027), .A2(KEYINPUT126), .ZN(new_n1028));
  INV_X1    g842(.A(KEYINPUT126), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1026), .A2(new_n1029), .A3(new_n714), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1024), .B1(new_n1028), .B2(new_n1030), .ZN(G57));
endmodule


