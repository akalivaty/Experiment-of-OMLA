//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(new_n188), .B(KEYINPUT82), .Z(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n193), .A2(new_n195), .A3(KEYINPUT0), .A4(G128), .ZN(new_n196));
  XNOR2_X1  g010(.A(G143), .B(G146), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT0), .B(G128), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n196), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT83), .B(G101), .ZN(new_n201));
  INV_X1    g015(.A(G104), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT3), .B1(new_n202), .B2(G107), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n204));
  INV_X1    g018(.A(G107), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(G104), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(G107), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n201), .A2(new_n203), .A3(new_n206), .A4(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n203), .A2(new_n206), .A3(new_n207), .ZN(new_n209));
  AOI22_X1  g023(.A1(new_n208), .A2(KEYINPUT4), .B1(G101), .B2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(KEYINPUT4), .A3(G101), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n200), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT84), .ZN(new_n214));
  XNOR2_X1  g028(.A(G104), .B(G107), .ZN(new_n215));
  INV_X1    g029(.A(G101), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n202), .A2(G107), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n205), .A2(G104), .ZN(new_n219));
  OAI211_X1 g033(.A(KEYINPUT84), .B(G101), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT1), .B1(new_n194), .B2(G146), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n194), .A2(G146), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n192), .A2(G143), .ZN(new_n224));
  OAI211_X1 g038(.A(G128), .B(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G128), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n193), .B(new_n195), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AND2_X1   g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n221), .A2(KEYINPUT10), .A3(new_n228), .A4(new_n208), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT10), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n217), .A2(new_n208), .A3(new_n220), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n225), .A2(new_n227), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT11), .ZN(new_n234));
  INV_X1    g048(.A(G134), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n234), .B1(new_n235), .B2(G137), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(G137), .ZN(new_n237));
  INV_X1    g051(.A(G137), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(KEYINPUT11), .A3(G134), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n236), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G131), .ZN(new_n241));
  INV_X1    g055(.A(G131), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n236), .A2(new_n239), .A3(new_n242), .A4(new_n237), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n241), .A2(KEYINPUT64), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT64), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n240), .A2(new_n245), .A3(G131), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n213), .A2(new_n229), .A3(new_n233), .A4(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT72), .B(G953), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G227), .ZN(new_n250));
  XOR2_X1   g064(.A(G110), .B(G140), .Z(new_n251));
  XOR2_X1   g065(.A(new_n250), .B(new_n251), .Z(new_n252));
  NAND2_X1  g066(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n244), .A2(new_n246), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n231), .A2(new_n232), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n231), .A2(new_n232), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n254), .B(KEYINPUT12), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT12), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n253), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n213), .A2(new_n229), .A3(new_n233), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n254), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n252), .B1(new_n263), .B2(new_n248), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n190), .B(new_n191), .C1(new_n261), .C2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(G469), .A2(G902), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n260), .A2(new_n257), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n252), .B1(new_n268), .B2(new_n248), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n253), .B1(new_n254), .B2(new_n262), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT85), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n253), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(new_n263), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT85), .ZN(new_n274));
  INV_X1    g088(.A(new_n248), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n275), .B1(new_n257), .B2(new_n260), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n273), .B(new_n274), .C1(new_n276), .C2(new_n252), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n271), .A2(G469), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n189), .B1(new_n267), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(G113), .B(G122), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n280), .B(new_n202), .ZN(new_n281));
  NAND2_X1  g095(.A1(KEYINPUT76), .A2(G125), .ZN(new_n282));
  INV_X1    g096(.A(G140), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(KEYINPUT76), .A2(G125), .A3(G140), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(KEYINPUT16), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n283), .A2(G125), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT16), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G146), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n284), .A2(KEYINPUT19), .A3(new_n285), .ZN(new_n292));
  INV_X1    g106(.A(G125), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G140), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT19), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n287), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n292), .A2(new_n296), .A3(new_n192), .ZN(new_n297));
  INV_X1    g111(.A(G953), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT72), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G953), .ZN(new_n301));
  INV_X1    g115(.A(G237), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n299), .A2(new_n301), .A3(G214), .A4(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n194), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n249), .A2(G143), .A3(G214), .A4(new_n302), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n305), .A3(new_n242), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n242), .B1(new_n304), .B2(new_n305), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n291), .B(new_n297), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n304), .A2(new_n305), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT18), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n311), .A2(new_n242), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n284), .A2(G146), .A3(new_n285), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n287), .A2(new_n294), .A3(new_n192), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n304), .B(new_n305), .C1(new_n311), .C2(new_n242), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n313), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n281), .B1(new_n309), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n286), .A2(new_n192), .A3(new_n289), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n291), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n321), .B1(KEYINPUT17), .B2(new_n308), .ZN(new_n322));
  INV_X1    g136(.A(new_n308), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT17), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(new_n324), .A3(new_n306), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n317), .A2(new_n316), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n322), .A2(new_n325), .B1(new_n326), .B2(new_n313), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n319), .B1(new_n327), .B2(new_n281), .ZN(new_n328));
  INV_X1    g142(.A(G475), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n191), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT20), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n319), .ZN(new_n332));
  NOR3_X1   g146(.A1(new_n307), .A2(KEYINPUT17), .A3(new_n308), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n291), .A2(new_n320), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n308), .A2(KEYINPUT17), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n281), .B(new_n318), .C1(new_n333), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT20), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n338), .A2(new_n339), .A3(new_n329), .A4(new_n191), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n331), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n337), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n322), .A2(new_n325), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n281), .B1(new_n343), .B2(new_n318), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n191), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT89), .ZN(new_n346));
  OAI21_X1  g160(.A(G475), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n318), .B1(new_n333), .B2(new_n336), .ZN(new_n348));
  INV_X1    g162(.A(new_n281), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(G902), .B1(new_n350), .B2(new_n337), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n351), .A2(KEYINPUT89), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n341), .B1(new_n347), .B2(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n226), .A2(G143), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT13), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n235), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n194), .A2(G128), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n226), .A2(G143), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(KEYINPUT13), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n357), .A2(new_n358), .A3(new_n235), .ZN(new_n360));
  AOI22_X1  g174(.A1(new_n356), .A2(new_n359), .B1(new_n360), .B2(KEYINPUT90), .ZN(new_n361));
  OR2_X1    g175(.A1(new_n360), .A2(KEYINPUT90), .ZN(new_n362));
  INV_X1    g176(.A(G116), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT68), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT68), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G116), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(new_n366), .A3(G122), .ZN(new_n367));
  OR2_X1    g181(.A1(new_n363), .A2(G122), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n367), .A2(new_n205), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n205), .B1(new_n367), .B2(new_n368), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n361), .B(new_n362), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n367), .A2(new_n205), .A3(new_n368), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n357), .A2(new_n358), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G134), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n360), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT14), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n367), .A2(new_n376), .A3(new_n368), .ZN(new_n377));
  OAI21_X1  g191(.A(G107), .B1(new_n367), .B2(new_n376), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n372), .B(new_n375), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n371), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G217), .ZN(new_n381));
  NOR3_X1   g195(.A1(new_n187), .A2(new_n381), .A3(G953), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n371), .A2(new_n379), .A3(new_n382), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(KEYINPUT91), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT91), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n380), .A2(new_n387), .A3(new_n383), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n191), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G478), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n390), .A2(KEYINPUT15), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n391), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n386), .A2(new_n191), .A3(new_n388), .A4(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n353), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G952), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n397), .A2(G953), .ZN(new_n398));
  INV_X1    g212(.A(G234), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n398), .B1(new_n399), .B2(new_n302), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  AOI211_X1 g215(.A(new_n191), .B(new_n249), .C1(G234), .C2(G237), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT21), .B(G898), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(G214), .B1(G237), .B2(G902), .ZN(new_n406));
  XOR2_X1   g220(.A(new_n406), .B(KEYINPUT86), .Z(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(G210), .B1(G237), .B2(G902), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(G110), .B(G122), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  OR2_X1    g226(.A1(KEYINPUT67), .A2(G119), .ZN(new_n413));
  NAND2_X1  g227(.A1(KEYINPUT67), .A2(G119), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(G116), .A3(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n364), .A2(new_n366), .A3(G119), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT69), .ZN(new_n418));
  NOR2_X1   g232(.A1(KEYINPUT2), .A2(G113), .ZN(new_n419));
  NAND2_X1  g233(.A1(KEYINPUT2), .A2(G113), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT66), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(KEYINPUT66), .A2(KEYINPUT2), .A3(G113), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n419), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT69), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n415), .A2(new_n416), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n418), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n424), .A2(new_n415), .A3(new_n416), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n208), .A2(KEYINPUT4), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n209), .A2(G101), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n428), .A2(new_n429), .B1(new_n432), .B2(new_n211), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n429), .A2(new_n208), .A3(new_n220), .A4(new_n217), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n415), .A2(new_n416), .A3(new_n426), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n426), .B1(new_n415), .B2(new_n416), .ZN(new_n436));
  OAI21_X1  g250(.A(KEYINPUT5), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(G113), .B1(new_n415), .B2(KEYINPUT5), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n434), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n412), .B1(new_n433), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n428), .A2(new_n429), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n432), .A2(new_n211), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n429), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n231), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT5), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(new_n418), .B2(new_n427), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n446), .B1(new_n448), .B2(new_n438), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n444), .A2(new_n449), .A3(new_n411), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n441), .A2(new_n450), .A3(KEYINPUT6), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n232), .A2(new_n293), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n452), .B1(new_n293), .B2(new_n200), .ZN(new_n453));
  XOR2_X1   g267(.A(KEYINPUT87), .B(G224), .Z(new_n454));
  NOR2_X1   g268(.A1(new_n454), .A2(G953), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n453), .B(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT6), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n457), .B(new_n412), .C1(new_n433), .C2(new_n440), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n451), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  XOR2_X1   g273(.A(new_n411), .B(KEYINPUT8), .Z(new_n460));
  NAND2_X1  g274(.A1(new_n437), .A2(new_n439), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n429), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n231), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n438), .A2(KEYINPUT88), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT88), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n465), .B(G113), .C1(new_n415), .C2(KEYINPUT5), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n464), .B(new_n466), .C1(new_n447), .C2(new_n417), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n446), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n460), .B1(new_n463), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(KEYINPUT7), .B1(new_n454), .B2(G953), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n453), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n470), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n452), .B(new_n472), .C1(new_n293), .C2(new_n200), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n450), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n191), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n410), .B1(new_n459), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n471), .A2(new_n473), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n433), .A2(new_n440), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n477), .B1(new_n478), .B2(new_n411), .ZN(new_n479));
  INV_X1    g293(.A(new_n460), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n461), .A2(new_n429), .B1(new_n208), .B2(new_n221), .ZN(new_n481));
  INV_X1    g295(.A(new_n468), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(G902), .B1(new_n479), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n451), .A2(new_n456), .A3(new_n458), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n485), .A3(new_n409), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n408), .B1(new_n476), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n279), .A2(new_n396), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT92), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n249), .A2(G210), .A3(new_n302), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT26), .B(G101), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n490), .B(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT73), .B(KEYINPUT27), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n492), .B(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n235), .A2(G137), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n238), .A2(G134), .ZN(new_n497));
  OAI21_X1  g311(.A(G131), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n225), .A2(new_n243), .A3(new_n498), .A4(new_n227), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT71), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n499), .B(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n244), .A2(new_n246), .A3(new_n200), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT70), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT70), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n244), .A2(new_n200), .A3(new_n504), .A4(new_n246), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n435), .A2(new_n436), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n445), .B1(new_n506), .B2(new_n425), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n501), .A2(new_n503), .A3(new_n505), .A4(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n499), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n510), .B1(new_n502), .B2(KEYINPUT65), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT65), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n244), .A2(new_n200), .A3(new_n512), .A4(new_n246), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n507), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT28), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n442), .A2(new_n510), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT28), .B1(new_n516), .B2(new_n502), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n495), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n508), .A2(new_n495), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT74), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n508), .A2(KEYINPUT74), .A3(new_n495), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n502), .A2(KEYINPUT65), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(new_n499), .A3(new_n513), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT30), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n501), .A2(new_n503), .A3(KEYINPUT30), .A4(new_n505), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n442), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(KEYINPUT31), .B1(new_n525), .B2(new_n531), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n508), .A2(KEYINPUT74), .A3(new_n495), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT74), .B1(new_n508), .B2(new_n495), .ZN(new_n534));
  OAI211_X1 g348(.A(KEYINPUT31), .B(new_n531), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n520), .B1(new_n532), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT75), .ZN(new_n538));
  NOR2_X1   g352(.A1(G472), .A2(G902), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT32), .A4(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT31), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n519), .B1(new_n543), .B2(new_n535), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n539), .A2(KEYINPUT32), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT75), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT32), .ZN(new_n547));
  INV_X1    g361(.A(new_n539), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n547), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n515), .A2(new_n518), .A3(new_n495), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n495), .B1(new_n531), .B2(new_n508), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n550), .A2(new_n551), .A3(KEYINPUT29), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n501), .A2(new_n503), .A3(new_n505), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n508), .B1(new_n554), .B2(new_n507), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n517), .B1(new_n555), .B2(KEYINPUT28), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n495), .A2(KEYINPUT29), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n191), .ZN(new_n559));
  OAI21_X1  g373(.A(G472), .B1(new_n552), .B2(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n540), .A2(new_n546), .A3(new_n549), .A4(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT78), .ZN(new_n562));
  AND2_X1   g376(.A1(KEYINPUT67), .A2(G119), .ZN(new_n563));
  NOR2_X1   g377(.A1(KEYINPUT67), .A2(G119), .ZN(new_n564));
  OAI21_X1  g378(.A(G128), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(G119), .A2(G128), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(KEYINPUT23), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(G110), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n226), .B1(new_n563), .B2(new_n564), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT23), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n568), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n413), .A2(new_n414), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n566), .B1(new_n574), .B2(G128), .ZN(new_n575));
  XNOR2_X1  g389(.A(KEYINPUT24), .B(G110), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n192), .B1(new_n286), .B2(new_n289), .ZN(new_n579));
  INV_X1    g393(.A(new_n315), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT77), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT77), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n578), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n569), .B1(new_n568), .B2(new_n572), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n575), .A2(new_n576), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n583), .A2(new_n585), .B1(new_n321), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n249), .A2(G221), .A3(G234), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT22), .B(G137), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n562), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n588), .A2(new_n321), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n578), .A2(new_n584), .A3(new_n581), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n584), .B1(new_n578), .B2(new_n581), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n592), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n597), .A2(KEYINPUT78), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(KEYINPUT79), .B1(new_n597), .B2(new_n598), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n583), .A2(new_n585), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT79), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n602), .A2(new_n603), .A3(new_n594), .A4(new_n592), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n600), .A2(new_n191), .A3(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n607), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n600), .A2(new_n191), .A3(new_n605), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n608), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n381), .B1(G234), .B2(new_n191), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(G902), .ZN(new_n614));
  XOR2_X1   g428(.A(new_n614), .B(KEYINPUT81), .Z(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n600), .A2(new_n605), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n612), .A2(new_n613), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT92), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n279), .A2(new_n396), .A3(new_n619), .A4(new_n487), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n489), .A2(new_n561), .A3(new_n618), .A4(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(new_n621), .B(new_n201), .Z(G3));
  OAI21_X1  g436(.A(G472), .B1(new_n544), .B2(G902), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n537), .A2(new_n539), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n626), .A2(new_n618), .A3(new_n279), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT93), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n476), .A2(KEYINPUT94), .A3(new_n486), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT94), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n484), .A2(new_n485), .A3(new_n630), .A4(new_n409), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n631), .A2(new_n406), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT33), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n386), .A2(new_n634), .A3(new_n388), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n390), .A2(G902), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n634), .B1(new_n380), .B2(new_n383), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n637), .A2(KEYINPUT95), .A3(new_n385), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(KEYINPUT95), .B1(new_n637), .B2(new_n385), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n635), .B(new_n636), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT96), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n640), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n638), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n645), .A2(KEYINPUT96), .A3(new_n635), .A4(new_n636), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n389), .A2(new_n390), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n643), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n353), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n633), .A2(new_n649), .A3(new_n404), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n628), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT34), .B(G104), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  NAND3_X1  g467(.A1(new_n629), .A2(new_n632), .A3(new_n405), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n341), .B(new_n395), .C1(new_n347), .C2(new_n352), .ZN(new_n655));
  OAI21_X1  g469(.A(KEYINPUT97), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n631), .A2(new_n406), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n484), .A2(new_n485), .A3(new_n409), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n409), .B1(new_n484), .B2(new_n485), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n657), .B1(new_n660), .B2(KEYINPUT94), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT97), .ZN(new_n662));
  INV_X1    g476(.A(new_n655), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n661), .A2(new_n662), .A3(new_n405), .A4(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n656), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n628), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT35), .B(G107), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  NAND2_X1  g482(.A1(new_n612), .A2(new_n613), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n598), .A2(KEYINPUT36), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n597), .B(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n616), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n489), .A2(new_n626), .A3(new_n620), .A4(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT37), .B(G110), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT98), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n674), .B(new_n676), .ZN(G12));
  INV_X1    g491(.A(G900), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n401), .B1(new_n402), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n655), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n661), .A2(new_n680), .A3(KEYINPUT99), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT99), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n329), .B1(new_n351), .B2(KEYINPUT89), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n345), .A2(new_n346), .ZN(new_n684));
  AOI22_X1  g498(.A1(new_n683), .A2(new_n684), .B1(new_n331), .B2(new_n340), .ZN(new_n685));
  INV_X1    g499(.A(new_n679), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n685), .A2(new_n395), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n682), .B1(new_n633), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n681), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n689), .A2(new_n561), .A3(new_n279), .A4(new_n673), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G128), .ZN(G30));
  AND2_X1   g505(.A1(new_n540), .A2(new_n546), .ZN(new_n692));
  INV_X1    g506(.A(new_n541), .ZN(new_n693));
  INV_X1    g507(.A(new_n495), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n693), .B1(new_n694), .B2(new_n555), .ZN(new_n695));
  OAI21_X1  g509(.A(G472), .B1(new_n695), .B2(G902), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n696), .A2(new_n549), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n673), .B1(new_n692), .B2(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(new_n679), .B(KEYINPUT39), .Z(new_n699));
  NAND2_X1  g513(.A1(new_n279), .A2(new_n699), .ZN(new_n700));
  OR2_X1    g514(.A1(new_n700), .A2(KEYINPUT40), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(KEYINPUT40), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT38), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n703), .B1(new_n658), .B2(new_n659), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n476), .A2(KEYINPUT38), .A3(new_n486), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n406), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n353), .A2(new_n395), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n698), .A2(new_n701), .A3(new_n702), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT100), .B(G143), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G45));
  NAND3_X1  g526(.A1(new_n648), .A2(new_n353), .A3(new_n686), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT101), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT101), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n648), .A2(new_n353), .A3(new_n715), .A4(new_n686), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n661), .A3(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n718), .A2(new_n561), .A3(new_n279), .A4(new_n673), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G146), .ZN(G48));
  INV_X1    g534(.A(KEYINPUT103), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n263), .A2(new_n248), .ZN(new_n722));
  INV_X1    g536(.A(new_n252), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n268), .A2(new_n272), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g538(.A(G469), .B1(new_n724), .B2(G902), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT102), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n725), .A2(new_n726), .A3(new_n265), .ZN(new_n727));
  OAI211_X1 g541(.A(KEYINPUT102), .B(G469), .C1(new_n724), .C2(G902), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n721), .B1(new_n729), .B2(new_n188), .ZN(new_n730));
  INV_X1    g544(.A(new_n188), .ZN(new_n731));
  AOI211_X1 g545(.A(KEYINPUT103), .B(new_n731), .C1(new_n727), .C2(new_n728), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n733), .A2(new_n561), .A3(new_n618), .A4(new_n650), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT41), .B(G113), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G15));
  NAND4_X1  g550(.A1(new_n665), .A2(new_n561), .A3(new_n618), .A4(new_n733), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G116), .ZN(G18));
  NAND2_X1  g552(.A1(new_n729), .A2(new_n188), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(new_n633), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n353), .A2(new_n395), .A3(new_n404), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n561), .A2(new_n740), .A3(new_n673), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G119), .ZN(G21));
  OAI22_X1  g557(.A1(new_n532), .A2(new_n536), .B1(new_n495), .B2(new_n556), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n539), .B(KEYINPUT104), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT105), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n623), .A2(new_n748), .ZN(new_n749));
  OAI211_X1 g563(.A(KEYINPUT105), .B(G472), .C1(new_n544), .C2(G902), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n747), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n654), .A2(new_n708), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n751), .A2(new_n733), .A3(new_n618), .A4(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G122), .ZN(G24));
  AND2_X1   g568(.A1(new_n714), .A2(new_n716), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n751), .A2(new_n755), .A3(new_n673), .A4(new_n740), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G125), .ZN(G27));
  NAND3_X1  g571(.A1(new_n476), .A2(new_n486), .A3(new_n406), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT107), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n476), .A2(KEYINPUT107), .A3(new_n486), .A4(new_n406), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n266), .B(KEYINPUT106), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n269), .A2(new_n270), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n763), .B1(new_n764), .B2(G469), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n731), .B1(new_n765), .B2(new_n265), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n760), .A2(new_n761), .A3(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n716), .A3(new_n714), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT42), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT108), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n537), .A2(new_n771), .A3(KEYINPUT32), .A4(new_n539), .ZN(new_n772));
  OAI21_X1  g586(.A(KEYINPUT108), .B1(new_n544), .B2(new_n545), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n549), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT109), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n772), .A2(new_n549), .A3(new_n773), .A4(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n775), .A2(new_n560), .A3(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n770), .A2(new_n778), .A3(new_n618), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n561), .A2(new_n767), .A3(new_n618), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n714), .A2(new_n716), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n769), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G131), .ZN(G33));
  NAND4_X1  g598(.A1(new_n561), .A2(new_n767), .A3(new_n618), .A4(new_n680), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G134), .ZN(G36));
  NAND2_X1  g600(.A1(new_n760), .A2(new_n761), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT112), .ZN(new_n788));
  AOI21_X1  g602(.A(KEYINPUT43), .B1(new_n648), .B2(new_n685), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n685), .A2(KEYINPUT111), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT111), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n353), .A2(new_n791), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n648), .A2(KEYINPUT43), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n789), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n673), .A2(new_n625), .ZN(new_n797));
  OAI21_X1  g611(.A(KEYINPUT44), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n789), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n790), .A2(new_n792), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n799), .B1(new_n800), .B2(new_n794), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT44), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n801), .A2(new_n802), .A3(new_n625), .A4(new_n673), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n788), .B1(new_n798), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n764), .A2(KEYINPUT45), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(G469), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT45), .B1(new_n271), .B2(new_n277), .ZN(new_n807));
  OAI211_X1 g621(.A(KEYINPUT46), .B(new_n762), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(KEYINPUT110), .A3(new_n265), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n806), .A2(new_n807), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(new_n763), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n809), .B1(KEYINPUT46), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT110), .B1(new_n808), .B2(new_n265), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n188), .B(new_n699), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n804), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G137), .ZN(G39));
  OAI21_X1  g631(.A(new_n188), .B1(new_n812), .B2(new_n813), .ZN(new_n818));
  OR2_X1    g632(.A1(KEYINPUT113), .A2(KEYINPUT47), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XOR2_X1   g634(.A(KEYINPUT113), .B(KEYINPUT47), .Z(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n188), .B(new_n822), .C1(new_n812), .C2(new_n813), .ZN(new_n823));
  NOR4_X1   g637(.A1(new_n781), .A2(new_n561), .A3(new_n618), .A4(new_n787), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n820), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT114), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n825), .B(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G140), .ZN(G42));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n561), .A2(new_n279), .A3(new_n673), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n681), .A2(new_n688), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n537), .A2(new_n191), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT105), .B1(new_n832), .B2(G472), .ZN(new_n833));
  INV_X1    g647(.A(new_n750), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n673), .B(new_n746), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n731), .B1(new_n727), .B2(new_n728), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n714), .A2(new_n661), .A3(new_n716), .A4(new_n836), .ZN(new_n837));
  OAI22_X1  g651(.A1(new_n830), .A2(new_n831), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n673), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n765), .A2(new_n265), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(new_n188), .A3(new_n686), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n841), .A2(new_n633), .A3(new_n708), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n540), .A2(new_n546), .A3(new_n696), .A4(new_n549), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n839), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n844), .B1(new_n830), .B2(new_n717), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT117), .B1(new_n838), .B2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(KEYINPUT116), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT116), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n849), .B1(new_n838), .B2(new_n845), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT52), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n719), .A2(new_n756), .A3(new_n690), .A4(new_n844), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n849), .B1(new_n852), .B2(KEYINPUT117), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n848), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n392), .A2(KEYINPUT115), .A3(new_n394), .ZN(new_n855));
  AOI21_X1  g669(.A(KEYINPUT115), .B1(new_n392), .B2(new_n394), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n686), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n857), .A2(new_n353), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n858), .A2(new_n760), .A3(new_n761), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n561), .A2(new_n859), .A3(new_n279), .A4(new_n673), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n860), .B(new_n785), .C1(new_n835), .C2(new_n768), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(new_n779), .B2(new_n782), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n737), .A2(new_n753), .A3(new_n734), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n279), .A2(new_n487), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n855), .A2(new_n856), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n649), .B1(new_n865), .B2(new_n353), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n626), .A2(new_n864), .A3(new_n618), .A4(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n621), .A2(new_n674), .A3(new_n742), .A4(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n862), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n829), .B1(new_n854), .B2(new_n870), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n561), .A2(new_n279), .A3(new_n673), .ZN(new_n872));
  AOI22_X1  g686(.A1(new_n872), .A2(new_n718), .B1(new_n698), .B2(new_n842), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n873), .A2(new_n847), .A3(new_n690), .A4(new_n756), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT52), .B1(new_n838), .B2(new_n845), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n862), .A2(new_n874), .A3(new_n869), .A4(new_n875), .ZN(new_n876));
  OR2_X1    g690(.A1(new_n876), .A2(new_n829), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n871), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(KEYINPUT54), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n862), .A2(new_n869), .A3(KEYINPUT53), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n846), .A2(KEYINPUT116), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n847), .B1(new_n852), .B2(new_n849), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n880), .A2(new_n883), .A3(new_n848), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT54), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n876), .A2(new_n829), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n884), .A2(KEYINPUT118), .A3(new_n885), .A4(new_n886), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n751), .A2(new_n618), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n796), .A2(new_n400), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n892), .A2(new_n740), .A3(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n843), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n787), .A2(new_n739), .A3(new_n400), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n895), .A2(new_n896), .A3(new_n618), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n894), .B(new_n398), .C1(new_n649), .C2(new_n897), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n778), .A2(new_n618), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n760), .A2(new_n761), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n901), .A2(new_n401), .A3(new_n836), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n900), .B1(new_n902), .B2(new_n796), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n896), .A2(new_n801), .A3(KEYINPUT120), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n899), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT48), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT48), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n899), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n898), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n835), .B1(new_n903), .B2(new_n904), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n648), .A2(new_n353), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n897), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n836), .A2(new_n706), .A3(new_n707), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT119), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n915), .B(new_n916), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n892), .A2(new_n917), .A3(KEYINPUT50), .A4(new_n893), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT50), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n751), .A2(new_n801), .A3(new_n618), .A4(new_n401), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n915), .B(KEYINPUT119), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n189), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n727), .B2(new_n728), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n925), .B1(new_n820), .B2(new_n823), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n920), .A2(new_n788), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n914), .B(new_n923), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT51), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n910), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT121), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n928), .A2(KEYINPUT121), .A3(new_n929), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n879), .A2(new_n889), .A3(new_n890), .A4(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n397), .A2(new_n298), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n706), .A2(new_n924), .A3(new_n407), .A4(new_n648), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n939), .A2(new_n800), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n729), .B(KEYINPUT49), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n940), .A2(new_n895), .A3(new_n618), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n938), .A2(new_n942), .ZN(G75));
  NAND2_X1  g757(.A1(new_n884), .A2(new_n886), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n944), .A2(G210), .A3(G902), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n451), .A2(new_n458), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(new_n456), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT55), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT122), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n949), .A2(KEYINPUT56), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n945), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n948), .B1(new_n945), .B2(new_n950), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n249), .A2(G952), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(G51));
  XOR2_X1   g768(.A(new_n762), .B(KEYINPUT57), .Z(new_n955));
  AND3_X1   g769(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n885), .B1(new_n884), .B2(new_n886), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n264), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n272), .A2(new_n268), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n944), .A2(G902), .A3(new_n810), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n953), .B1(new_n962), .B2(new_n963), .ZN(G54));
  NAND2_X1  g778(.A1(KEYINPUT58), .A2(G475), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n944), .A2(G902), .A3(new_n966), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n967), .A2(new_n328), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n967), .A2(new_n328), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n968), .A2(new_n969), .A3(new_n953), .ZN(G60));
  NAND2_X1  g784(.A1(G478), .A2(G902), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT59), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n645), .A2(new_n635), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n973), .B1(new_n956), .B2(new_n957), .ZN(new_n974));
  INV_X1    g788(.A(new_n953), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n876), .A2(new_n829), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n862), .A2(new_n869), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n883), .A2(new_n978), .A3(new_n848), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n977), .B1(new_n979), .B2(new_n829), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n890), .B1(new_n980), .B2(new_n885), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n887), .A2(new_n888), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n972), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n645), .A2(new_n635), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n976), .B1(new_n983), .B2(new_n984), .ZN(G63));
  INV_X1    g799(.A(KEYINPUT61), .ZN(new_n986));
  NAND2_X1  g800(.A1(G217), .A2(G902), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT123), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT60), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n944), .A2(new_n671), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n975), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n617), .B(KEYINPUT124), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n993), .B1(new_n944), .B2(new_n989), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n986), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n994), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n996), .A2(KEYINPUT61), .A3(new_n975), .A4(new_n990), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n995), .A2(new_n997), .ZN(G66));
  OAI21_X1  g812(.A(G953), .B1(new_n454), .B2(new_n403), .ZN(new_n999));
  INV_X1    g813(.A(new_n249), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n999), .B1(new_n869), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n946), .B1(G898), .B2(new_n249), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1001), .B(new_n1002), .ZN(G69));
  AOI21_X1  g817(.A(new_n249), .B1(G227), .B2(G900), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  AND2_X1   g819(.A1(new_n529), .A2(new_n530), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n292), .A2(new_n296), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1006), .B(new_n1007), .Z(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(new_n785), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1010), .B1(new_n804), .B2(new_n815), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n838), .B1(new_n872), .B2(new_n718), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n633), .A2(new_n708), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n815), .A2(new_n899), .A3(new_n1013), .ZN(new_n1014));
  AND4_X1   g828(.A1(new_n783), .A2(new_n1011), .A3(new_n1012), .A4(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(new_n827), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n249), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1000), .A2(new_n678), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1018), .B(KEYINPUT125), .Z(new_n1019));
  AOI21_X1  g833(.A(new_n1009), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n710), .A2(new_n690), .A3(new_n719), .A4(new_n756), .ZN(new_n1021));
  XOR2_X1   g835(.A(new_n1021), .B(KEYINPUT62), .Z(new_n1022));
  INV_X1    g836(.A(new_n700), .ZN(new_n1023));
  AND2_X1   g837(.A1(new_n1023), .A2(new_n866), .ZN(new_n1024));
  NAND4_X1  g838(.A1(new_n1024), .A2(new_n561), .A3(new_n618), .A4(new_n901), .ZN(new_n1025));
  AND2_X1   g839(.A1(new_n816), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1022), .A2(new_n827), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1008), .B1(new_n1027), .B2(new_n249), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1005), .B1(new_n1020), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1000), .B1(new_n1015), .B2(new_n827), .ZN(new_n1030));
  INV_X1    g844(.A(new_n1019), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1008), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AND2_X1   g846(.A1(new_n1027), .A2(new_n249), .ZN(new_n1033));
  OAI211_X1 g847(.A(new_n1032), .B(new_n1004), .C1(new_n1033), .C2(new_n1008), .ZN(new_n1034));
  AND2_X1   g848(.A1(new_n1029), .A2(new_n1034), .ZN(G72));
  NAND3_X1  g849(.A1(new_n1015), .A2(new_n827), .A3(new_n869), .ZN(new_n1036));
  XNOR2_X1  g850(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1037));
  NAND2_X1  g851(.A1(G472), .A2(G902), .ZN(new_n1038));
  XNOR2_X1  g852(.A(new_n1037), .B(new_n1038), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g854(.A1(new_n1040), .A2(new_n508), .A3(new_n694), .A4(new_n531), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n1039), .B1(new_n693), .B2(new_n551), .ZN(new_n1042));
  OAI211_X1 g856(.A(new_n1041), .B(new_n975), .C1(new_n980), .C2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g857(.A1(new_n1022), .A2(new_n827), .A3(new_n869), .A4(new_n1026), .ZN(new_n1044));
  AND3_X1   g858(.A1(new_n1044), .A2(KEYINPUT127), .A3(new_n1039), .ZN(new_n1045));
  AOI21_X1  g859(.A(KEYINPUT127), .B1(new_n1044), .B2(new_n1039), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n531), .A2(new_n508), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n1047), .A2(new_n495), .ZN(new_n1048));
  NOR3_X1   g862(.A1(new_n1045), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  NOR2_X1   g863(.A1(new_n1043), .A2(new_n1049), .ZN(G57));
endmodule


