//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n785, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045;
  XNOR2_X1  g000(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n202));
  INV_X1    g001(.A(G155gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G183gat), .B(G211gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G57gat), .B(G64gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(G71gat), .A2(G78gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(G71gat), .A2(G78gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT9), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n209), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n211), .B(new_n210), .C1(new_n208), .C2(new_n213), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT21), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G231gat), .A2(G233gat), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n219), .B(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G127gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n219), .B(new_n220), .ZN(new_n224));
  INV_X1    g023(.A(G127gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G15gat), .B(G22gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT16), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n227), .B1(new_n228), .B2(G1gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(G1gat), .B2(new_n227), .ZN(new_n230));
  INV_X1    g029(.A(G8gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n230), .B(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(new_n218), .B2(new_n217), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n223), .A2(new_n226), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n233), .B1(new_n223), .B2(new_n226), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n207), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n223), .A2(new_n226), .ZN(new_n238));
  INV_X1    g037(.A(new_n233), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(new_n234), .A3(new_n206), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  XOR2_X1   g041(.A(G190gat), .B(G218gat), .Z(new_n243));
  NAND2_X1  g042(.A1(G99gat), .A2(G106gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT8), .ZN(new_n245));
  NAND2_X1  g044(.A1(G85gat), .A2(G92gat), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT7), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G85gat), .ZN(new_n249));
  INV_X1    g048(.A(G92gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n245), .A2(new_n248), .A3(new_n251), .A4(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G99gat), .B(G106gat), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT87), .ZN(new_n257));
  AOI22_X1  g056(.A1(KEYINPUT8), .A2(new_n244), .B1(new_n249), .B2(new_n250), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n258), .A2(new_n254), .A3(new_n248), .A4(new_n252), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n256), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n253), .A2(KEYINPUT87), .A3(new_n255), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(KEYINPUT88), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT88), .B1(new_n260), .B2(new_n261), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G43gat), .B(G50gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT15), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT14), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n269), .B(KEYINPUT84), .C1(G29gat), .C2(G36gat), .ZN(new_n270));
  INV_X1    g069(.A(G29gat), .ZN(new_n271));
  INV_X1    g070(.A(G36gat), .ZN(new_n272));
  OAI221_X1 g071(.A(new_n270), .B1(new_n271), .B2(new_n272), .C1(new_n266), .C2(KEYINPUT15), .ZN(new_n273));
  OR3_X1    g072(.A1(KEYINPUT84), .A2(G29gat), .A3(G36gat), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT84), .B1(G29gat), .B2(G36gat), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(KEYINPUT14), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n268), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  XOR2_X1   g077(.A(G43gat), .B(G50gat), .Z(new_n279));
  INV_X1    g078(.A(KEYINPUT15), .ZN(new_n280));
  AOI22_X1  g079(.A1(new_n279), .A2(new_n280), .B1(G29gat), .B2(G36gat), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n281), .A2(new_n267), .A3(new_n276), .A4(new_n270), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT85), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT17), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT17), .ZN(new_n286));
  AOI211_X1 g085(.A(KEYINPUT85), .B(new_n286), .C1(new_n278), .C2(new_n282), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n265), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n283), .B1(new_n263), .B2(new_n264), .ZN(new_n290));
  AND2_X1   g089(.A1(G232gat), .A2(G233gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT41), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n243), .B1(new_n289), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n291), .A2(KEYINPUT41), .ZN(new_n295));
  XNOR2_X1  g094(.A(G134gat), .B(G162gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n293), .ZN(new_n298));
  INV_X1    g097(.A(new_n243), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n288), .A3(new_n299), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n294), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n297), .B1(new_n294), .B2(new_n300), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n242), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT89), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT89), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n242), .B(new_n305), .C1(new_n301), .C2(new_n302), .ZN(new_n306));
  XOR2_X1   g105(.A(G120gat), .B(G148gat), .Z(new_n307));
  XNOR2_X1  g106(.A(new_n307), .B(KEYINPUT92), .ZN(new_n308));
  XNOR2_X1  g107(.A(G176gat), .B(G204gat), .ZN(new_n309));
  XOR2_X1   g108(.A(new_n308), .B(new_n309), .Z(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n260), .A2(new_n217), .A3(new_n261), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT90), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT90), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n260), .A2(new_n217), .A3(new_n314), .A4(new_n261), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n217), .B1(new_n255), .B2(new_n253), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n313), .A2(new_n315), .B1(new_n259), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT10), .ZN(new_n318));
  AND3_X1   g117(.A1(new_n317), .A2(KEYINPUT91), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT91), .B1(new_n317), .B2(new_n318), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT10), .ZN(new_n321));
  OAI22_X1  g120(.A1(new_n319), .A2(new_n320), .B1(new_n265), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G230gat), .A2(G233gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n317), .A2(new_n323), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n311), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  AOI211_X1 g126(.A(new_n325), .B(new_n310), .C1(new_n322), .C2(new_n323), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n304), .A2(new_n306), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT93), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT93), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n304), .A2(new_n329), .A3(new_n332), .A4(new_n306), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G120gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G113gat), .ZN(new_n336));
  INV_X1    g135(.A(G113gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(G120gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n338), .A3(KEYINPUT71), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT71), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(new_n337), .A3(G120gat), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT1), .ZN(new_n343));
  INV_X1    g142(.A(G134gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(G127gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n225), .A2(G134gat), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n342), .A2(new_n343), .A3(new_n345), .A4(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n346), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT1), .B1(new_n336), .B2(new_n338), .ZN(new_n350));
  OAI22_X1  g149(.A1(new_n340), .A2(new_n347), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(G169gat), .A2(G176gat), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT26), .ZN(new_n354));
  NAND2_X1  g153(.A1(G169gat), .A2(G176gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n352), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n357));
  INV_X1    g156(.A(G183gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT27), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT27), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(G183gat), .ZN(new_n361));
  INV_X1    g160(.A(G190gat), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n359), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n356), .B(new_n357), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n364), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT70), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n356), .A2(new_n357), .ZN(new_n369));
  OR2_X1    g168(.A1(new_n363), .A2(new_n364), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT70), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n369), .A2(new_n370), .A3(new_n371), .A4(new_n366), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n362), .ZN(new_n374));
  NAND3_X1  g173(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(G183gat), .A2(G190gat), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT24), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(KEYINPUT64), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n378), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT64), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n376), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n352), .A2(KEYINPUT23), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT23), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n385), .A2(G169gat), .A3(G176gat), .ZN(new_n386));
  INV_X1    g185(.A(new_n355), .ZN(new_n387));
  NOR3_X1   g186(.A1(new_n384), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT25), .B1(new_n383), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT67), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT65), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n391), .B1(new_n386), .B2(new_n387), .ZN(new_n392));
  INV_X1    g191(.A(G169gat), .ZN(new_n393));
  INV_X1    g192(.A(G176gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(new_n394), .A3(KEYINPUT23), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n395), .A2(KEYINPUT65), .A3(new_n355), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT25), .B1(new_n352), .B2(KEYINPUT23), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n392), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n374), .A2(new_n375), .ZN(new_n400));
  NAND3_X1  g199(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT66), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT24), .B1(new_n377), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n400), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n390), .B1(new_n399), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT65), .B1(new_n395), .B2(new_n355), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n406), .A2(new_n397), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n403), .A2(new_n401), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n376), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n407), .A2(new_n409), .A3(KEYINPUT67), .A4(new_n396), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n389), .B1(new_n405), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n373), .B1(new_n411), .B2(KEYINPUT68), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT68), .ZN(new_n413));
  AOI211_X1 g212(.A(new_n413), .B(new_n389), .C1(new_n405), .C2(new_n410), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n351), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n389), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n395), .A2(KEYINPUT65), .A3(new_n355), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n417), .A2(new_n406), .A3(new_n397), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT67), .B1(new_n418), .B2(new_n409), .ZN(new_n419));
  NOR3_X1   g218(.A1(new_n399), .A2(new_n390), .A3(new_n404), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n416), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n413), .ZN(new_n422));
  INV_X1    g221(.A(new_n347), .ZN(new_n423));
  INV_X1    g222(.A(new_n350), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n423), .A2(new_n339), .B1(new_n424), .B2(new_n348), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n411), .A2(KEYINPUT68), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n422), .A2(new_n425), .A3(new_n426), .A4(new_n373), .ZN(new_n427));
  NAND2_X1  g226(.A1(G227gat), .A2(G233gat), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n415), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT34), .B1(new_n429), .B2(KEYINPUT73), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n429), .A2(KEYINPUT73), .A3(KEYINPUT34), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  XOR2_X1   g232(.A(G15gat), .B(G43gat), .Z(new_n434));
  XNOR2_X1  g233(.A(G71gat), .B(G99gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n428), .B1(new_n415), .B2(new_n427), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n436), .B1(new_n437), .B2(KEYINPUT33), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT32), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n415), .A2(new_n427), .ZN(new_n442));
  INV_X1    g241(.A(new_n428), .ZN(new_n443));
  AOI221_X4 g242(.A(new_n439), .B1(KEYINPUT33), .B2(new_n436), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n433), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(G211gat), .B(G218gat), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(G211gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT75), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT75), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(G211gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT22), .B1(new_n452), .B2(G218gat), .ZN(new_n453));
  OR2_X1    g252(.A1(KEYINPUT74), .A2(G197gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(KEYINPUT74), .A2(G197gat), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(G204gat), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(G204gat), .ZN(new_n457));
  AND2_X1   g256(.A1(KEYINPUT74), .A2(G197gat), .ZN(new_n458));
  NOR2_X1   g257(.A1(KEYINPUT74), .A2(G197gat), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n447), .B1(new_n453), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT76), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT22), .ZN(new_n464));
  XNOR2_X1  g263(.A(KEYINPUT75), .B(G211gat), .ZN(new_n465));
  INV_X1    g264(.A(G218gat), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n467), .A2(new_n446), .A3(new_n456), .A4(new_n460), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n462), .A2(new_n463), .A3(new_n468), .ZN(new_n469));
  OAI211_X1 g268(.A(KEYINPUT76), .B(new_n447), .C1(new_n453), .C2(new_n461), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AND2_X1   g270(.A1(G155gat), .A2(G162gat), .ZN(new_n472));
  NOR2_X1   g271(.A1(G155gat), .A2(G162gat), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(G141gat), .B(G148gat), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT2), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n476), .B1(G155gat), .B2(G162gat), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n474), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(G141gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(G148gat), .ZN(new_n480));
  INV_X1    g279(.A(G148gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(G141gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(G155gat), .B(G162gat), .ZN(new_n484));
  INV_X1    g283(.A(G162gat), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT2), .B1(new_n203), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT3), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n478), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT29), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n471), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n478), .A2(new_n487), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT29), .B1(new_n462), .B2(new_n468), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n493), .B1(new_n494), .B2(KEYINPUT3), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(G228gat), .A2(G233gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n478), .A2(new_n487), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n469), .A2(new_n490), .A3(new_n470), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n499), .B1(new_n500), .B2(new_n488), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n492), .A2(G228gat), .A3(G233gat), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(G22gat), .ZN(new_n504));
  INV_X1    g303(.A(G22gat), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n498), .B(new_n505), .C1(new_n501), .C2(new_n502), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n506), .A2(KEYINPUT82), .ZN(new_n508));
  XNOR2_X1  g307(.A(G78gat), .B(G106gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT31), .B(G50gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n507), .B1(new_n508), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT82), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n504), .A2(new_n506), .A3(new_n514), .A4(new_n511), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n429), .A2(KEYINPUT73), .A3(KEYINPUT34), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n517), .A2(new_n430), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n368), .A2(new_n372), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n519), .B1(new_n421), .B2(new_n413), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n425), .B1(new_n520), .B2(new_n426), .ZN(new_n521));
  NOR3_X1   g320(.A1(new_n412), .A2(new_n351), .A3(new_n414), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n443), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT32), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT33), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n524), .A2(new_n526), .A3(new_n436), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n438), .A2(new_n440), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n518), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n445), .A2(new_n516), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n490), .B1(new_n412), .B2(new_n414), .ZN(new_n531));
  NAND2_X1  g330(.A1(G226gat), .A2(G233gat), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n531), .A2(KEYINPUT77), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n369), .A2(new_n370), .A3(new_n366), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n421), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n532), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n531), .A2(new_n532), .B1(new_n537), .B2(KEYINPUT77), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n471), .B1(new_n533), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G8gat), .B(G36gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(G64gat), .B(G92gat), .ZN(new_n541));
  XOR2_X1   g340(.A(new_n540), .B(new_n541), .Z(new_n542));
  NAND3_X1  g341(.A1(new_n520), .A2(new_n536), .A3(new_n426), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n535), .A2(new_n490), .A3(new_n532), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n471), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n539), .A2(new_n542), .A3(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(KEYINPUT78), .B(KEYINPUT30), .Z(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT4), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n425), .A2(new_n499), .A3(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT4), .B1(new_n351), .B2(new_n493), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT80), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n493), .A2(KEYINPUT3), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n555), .A2(new_n351), .A3(new_n489), .ZN(new_n556));
  OAI211_X1 g355(.A(KEYINPUT80), .B(KEYINPUT4), .C1(new_n351), .C2(new_n493), .ZN(new_n557));
  NAND2_X1  g356(.A1(G225gat), .A2(G233gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT79), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n559), .A2(KEYINPUT5), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n554), .A2(new_n556), .A3(new_n557), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT81), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n556), .A2(new_n557), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT81), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n563), .A2(new_n564), .A3(new_n554), .A4(new_n560), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n551), .A2(new_n552), .ZN(new_n566));
  INV_X1    g365(.A(new_n559), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n566), .A2(new_n567), .A3(new_n556), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT5), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n425), .A2(new_n499), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n351), .A2(new_n493), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n569), .B1(new_n572), .B2(new_n559), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n562), .A2(new_n565), .B1(new_n568), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G1gat), .B(G29gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT0), .ZN(new_n576));
  XNOR2_X1  g375(.A(G57gat), .B(G85gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  AOI21_X1  g377(.A(KEYINPUT6), .B1(new_n574), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n565), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n568), .A2(new_n573), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n578), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n582), .A2(KEYINPUT6), .A3(new_n583), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n542), .ZN(new_n588));
  INV_X1    g387(.A(new_n471), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n531), .A2(new_n532), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n537), .A2(KEYINPUT77), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n531), .A2(KEYINPUT77), .A3(new_n532), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n589), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n588), .B1(new_n594), .B2(new_n545), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n539), .A2(KEYINPUT30), .A3(new_n542), .A4(new_n546), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n549), .A2(new_n587), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n530), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(KEYINPUT72), .B1(new_n441), .B2(new_n444), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT72), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n527), .A2(new_n600), .A3(new_n528), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n599), .A2(new_n601), .A3(new_n433), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n602), .A2(new_n516), .A3(new_n529), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n595), .A2(new_n596), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n604), .A2(KEYINPUT35), .A3(new_n587), .A4(new_n549), .ZN(new_n605));
  OAI22_X1  g404(.A1(new_n598), .A2(KEYINPUT35), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n567), .B1(new_n563), .B2(new_n554), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT39), .B1(new_n572), .B2(new_n559), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT39), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n583), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT40), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  AND3_X1   g411(.A1(new_n609), .A2(KEYINPUT40), .A3(new_n611), .ZN(new_n613));
  AOI211_X1 g412(.A(new_n612), .B(new_n613), .C1(new_n583), .C2(new_n582), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n595), .A2(new_n596), .ZN(new_n615));
  INV_X1    g414(.A(new_n548), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n422), .A2(new_n426), .A3(new_n373), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n536), .B1(new_n617), .B2(new_n490), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n537), .A2(KEYINPUT77), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n593), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n545), .B1(new_n620), .B2(new_n471), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n616), .B1(new_n621), .B2(new_n542), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n614), .B1(new_n615), .B2(new_n622), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n547), .A2(new_n586), .A3(new_n585), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n589), .B1(new_n533), .B2(new_n538), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT37), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n543), .A2(new_n544), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n626), .B1(new_n627), .B2(new_n471), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT38), .B1(new_n625), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n542), .B1(new_n539), .B2(new_n546), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n542), .A2(new_n626), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n624), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n542), .B1(new_n621), .B2(new_n626), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT37), .B1(new_n594), .B2(new_n545), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n516), .B(new_n623), .C1(new_n633), .C2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n602), .A2(KEYINPUT36), .A3(new_n529), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT36), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n518), .A2(new_n527), .A3(new_n528), .ZN(new_n641));
  AOI22_X1  g440(.A1(new_n527), .A2(new_n528), .B1(new_n432), .B2(new_n431), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n516), .ZN(new_n644));
  AOI22_X1  g443(.A1(new_n639), .A2(new_n643), .B1(new_n644), .B2(new_n597), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n606), .B1(new_n638), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n232), .B1(new_n285), .B2(new_n287), .ZN(new_n647));
  NAND2_X1  g446(.A1(G229gat), .A2(G233gat), .ZN(new_n648));
  INV_X1    g447(.A(new_n232), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n283), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n647), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT18), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n647), .A2(KEYINPUT18), .A3(new_n648), .A4(new_n650), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n232), .B(new_n283), .Z(new_n655));
  XOR2_X1   g454(.A(new_n648), .B(KEYINPUT13), .Z(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n653), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(G113gat), .B(G141gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G197gat), .ZN(new_n660));
  XOR2_X1   g459(.A(KEYINPUT11), .B(G169gat), .Z(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n662), .B(KEYINPUT12), .Z(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  AND3_X1   g463(.A1(new_n658), .A2(KEYINPUT83), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n664), .B1(new_n658), .B2(KEYINPUT83), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT86), .B1(new_n646), .B2(new_n668), .ZN(new_n669));
  OR2_X1    g468(.A1(new_n530), .A2(new_n597), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT35), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n516), .A2(new_n529), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n527), .A2(new_n528), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n518), .B1(new_n673), .B2(KEYINPUT72), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n672), .B1(new_n601), .B2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n597), .A2(new_n671), .ZN(new_n676));
  AOI22_X1  g475(.A1(new_n670), .A2(new_n671), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n599), .A2(new_n601), .A3(new_n433), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n529), .A2(KEYINPUT36), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n643), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n597), .A2(new_n644), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n638), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT86), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n683), .A2(new_n684), .A3(new_n667), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n334), .B1(new_n669), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n587), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(G1gat), .ZN(G1324gat));
  INV_X1    g488(.A(KEYINPUT94), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n604), .A2(new_n549), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n231), .B1(new_n686), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n334), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n684), .B1(new_n683), .B2(new_n667), .ZN(new_n694));
  AOI211_X1 g493(.A(KEYINPUT86), .B(new_n668), .C1(new_n677), .C2(new_n682), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n691), .B(new_n693), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT16), .B(G8gat), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(KEYINPUT42), .B1(new_n692), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n669), .A2(new_n685), .ZN(new_n700));
  INV_X1    g499(.A(new_n697), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n700), .A2(new_n691), .A3(new_n693), .A4(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT42), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n690), .B1(new_n699), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n696), .A2(G8gat), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n703), .B1(new_n706), .B2(new_n702), .ZN(new_n707));
  INV_X1    g506(.A(new_n691), .ZN(new_n708));
  AOI211_X1 g507(.A(new_n708), .B(new_n334), .C1(new_n669), .C2(new_n685), .ZN(new_n709));
  AOI21_X1  g508(.A(KEYINPUT42), .B1(new_n709), .B2(new_n701), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n707), .A2(new_n710), .A3(KEYINPUT94), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n705), .A2(new_n711), .ZN(G1325gat));
  INV_X1    g511(.A(new_n680), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n686), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n445), .A2(new_n529), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(G15gat), .ZN(new_n716));
  AOI22_X1  g515(.A1(new_n714), .A2(G15gat), .B1(new_n686), .B2(new_n716), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(KEYINPUT95), .Z(G1326gat));
  NAND2_X1  g517(.A1(new_n686), .A2(new_n644), .ZN(new_n719));
  OR2_X1    g518(.A1(new_n719), .A2(KEYINPUT96), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(KEYINPUT96), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT43), .B(G22gat), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n720), .A2(new_n721), .A3(new_n723), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(G1327gat));
  INV_X1    g526(.A(new_n242), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n329), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n301), .A2(new_n302), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n700), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n733), .A2(new_n271), .A3(new_n687), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT45), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(new_n646), .B2(new_n731), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n683), .A2(KEYINPUT44), .A3(new_n730), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n729), .A2(new_n668), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(G29gat), .B1(new_n742), .B2(new_n587), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n734), .A2(new_n735), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n736), .A2(new_n743), .A3(new_n744), .ZN(G1328gat));
  NAND3_X1  g544(.A1(new_n733), .A2(new_n272), .A3(new_n691), .ZN(new_n746));
  OR2_X1    g545(.A1(new_n746), .A2(KEYINPUT46), .ZN(new_n747));
  OAI21_X1  g546(.A(G36gat), .B1(new_n742), .B2(new_n708), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(KEYINPUT46), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(G1329gat));
  OAI21_X1  g549(.A(G43gat), .B1(new_n742), .B2(new_n680), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n715), .A2(G43gat), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n733), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT97), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT47), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n751), .B(new_n753), .C1(new_n755), .C2(KEYINPUT47), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(G1330gat));
  NAND3_X1  g558(.A1(new_n700), .A2(new_n644), .A3(new_n732), .ZN(new_n760));
  INV_X1    g559(.A(G50gat), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n644), .A2(G50gat), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n742), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(KEYINPUT98), .B(KEYINPUT48), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(G1331gat));
  INV_X1    g565(.A(new_n329), .ZN(new_n767));
  AND4_X1   g566(.A1(new_n668), .A2(new_n767), .A3(new_n304), .A4(new_n306), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n683), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n687), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g570(.A(new_n708), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(new_n775));
  XOR2_X1   g574(.A(KEYINPUT99), .B(KEYINPUT100), .Z(new_n776));
  XNOR2_X1  g575(.A(new_n775), .B(new_n776), .ZN(G1333gat));
  NAND3_X1  g576(.A1(new_n769), .A2(G71gat), .A3(new_n713), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT101), .ZN(new_n779));
  INV_X1    g578(.A(G71gat), .ZN(new_n780));
  INV_X1    g579(.A(new_n769), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n780), .B1(new_n781), .B2(new_n715), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n644), .ZN(new_n785));
  XOR2_X1   g584(.A(KEYINPUT102), .B(G78gat), .Z(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(G1335gat));
  NOR2_X1   g586(.A1(new_n667), .A2(new_n242), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n683), .A2(new_n730), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n789), .B(new_n790), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n791), .A2(new_n767), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n792), .A2(new_n249), .A3(new_n687), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n788), .A2(new_n767), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT103), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n740), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(G85gat), .B1(new_n796), .B2(new_n587), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n793), .A2(new_n797), .ZN(G1336gat));
  NAND3_X1  g597(.A1(new_n791), .A2(new_n691), .A3(new_n767), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n250), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(KEYINPUT104), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n708), .A2(new_n250), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n738), .A2(new_n739), .A3(new_n795), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n801), .A2(KEYINPUT104), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n800), .A2(new_n803), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n803), .B1(new_n800), .B2(new_n807), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n808), .A2(new_n809), .ZN(G1337gat));
  NOR2_X1   g609(.A1(new_n715), .A2(G99gat), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n792), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(G99gat), .B1(new_n796), .B2(new_n680), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(G1338gat));
  NOR2_X1   g613(.A1(new_n516), .A2(G106gat), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n789), .A2(new_n790), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n789), .A2(new_n790), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n767), .B(new_n815), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT106), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n738), .A2(new_n644), .A3(new_n739), .A4(new_n795), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT105), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n821), .A2(new_n822), .A3(G106gat), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n818), .A2(new_n819), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT53), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n821), .A2(G106gat), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n822), .A2(KEYINPUT53), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n827), .B(new_n828), .C1(new_n818), .C2(KEYINPUT53), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n826), .A2(new_n829), .ZN(G1339gat));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n265), .A2(new_n321), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT91), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n313), .A2(new_n315), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n316), .A2(new_n259), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n833), .B1(new_n836), .B2(KEYINPUT10), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n317), .A2(KEYINPUT91), .A3(new_n318), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n832), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n323), .ZN(new_n840));
  OAI21_X1  g639(.A(KEYINPUT54), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n322), .A2(new_n323), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n322), .A2(new_n844), .A3(new_n323), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n310), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n831), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n839), .A2(new_n840), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n324), .A2(new_n848), .A3(KEYINPUT54), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n849), .A2(KEYINPUT55), .A3(new_n310), .A4(new_n845), .ZN(new_n850));
  INV_X1    g649(.A(new_n328), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n847), .A2(new_n667), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n648), .B1(new_n647), .B2(new_n650), .ZN(new_n853));
  OAI22_X1  g652(.A1(new_n853), .A2(KEYINPUT107), .B1(new_n655), .B2(new_n656), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n853), .A2(KEYINPUT107), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n662), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI221_X1 g655(.A(new_n856), .B1(new_n658), .B2(new_n663), .C1(new_n327), .C2(new_n328), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n852), .A2(KEYINPUT108), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT108), .B1(new_n852), .B2(new_n857), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n858), .A2(new_n859), .A3(new_n730), .ZN(new_n860));
  INV_X1    g659(.A(new_n847), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n850), .A2(new_n851), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n730), .B(new_n856), .C1(new_n658), .C2(new_n663), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n728), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n330), .A2(new_n667), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(new_n687), .A3(new_n675), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n869), .A2(new_n691), .ZN(new_n870));
  AOI21_X1  g669(.A(G113gat), .B1(new_n870), .B2(new_n667), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n852), .A2(new_n857), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT108), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n852), .A2(new_n857), .A3(KEYINPUT108), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n731), .A3(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n864), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n242), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(new_n866), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(new_n530), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n691), .A2(new_n587), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n882), .A2(new_n337), .A3(new_n668), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n871), .A2(new_n883), .ZN(G1340gat));
  AOI21_X1  g683(.A(G120gat), .B1(new_n870), .B2(new_n767), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n882), .A2(new_n335), .A3(new_n329), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n885), .A2(new_n886), .ZN(G1341gat));
  NAND4_X1  g686(.A1(new_n880), .A2(G127gat), .A3(new_n242), .A4(new_n881), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT109), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n888), .B(new_n889), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n869), .A2(new_n691), .A3(new_n728), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT110), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(G127gat), .B1(new_n891), .B2(new_n892), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n890), .B1(new_n893), .B2(new_n894), .ZN(G1342gat));
  NAND2_X1  g694(.A1(new_n708), .A2(new_n730), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT111), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n869), .A2(G134gat), .A3(new_n897), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT56), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n880), .A2(new_n730), .A3(new_n881), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT112), .B1(new_n900), .B2(G134gat), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n900), .A2(KEYINPUT112), .A3(G134gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(G1343gat));
  NAND2_X1  g702(.A1(new_n680), .A2(new_n881), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT57), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n905), .B1(new_n879), .B2(new_n516), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n516), .A2(new_n905), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n730), .B1(new_n852), .B2(new_n857), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n728), .B1(new_n909), .B2(new_n864), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n908), .B1(new_n910), .B2(new_n867), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n904), .B1(new_n906), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n479), .B1(new_n913), .B2(new_n667), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT113), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n713), .A2(new_n516), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n868), .A2(new_n687), .A3(new_n708), .A4(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n668), .A2(G141gat), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n915), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n687), .B(new_n916), .C1(new_n878), .C2(new_n866), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n921), .A2(new_n691), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(KEYINPUT113), .A3(new_n918), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(KEYINPUT58), .B1(new_n914), .B2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(new_n904), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT57), .B1(new_n868), .B2(new_n644), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n926), .B1(new_n927), .B2(new_n911), .ZN(new_n928));
  OAI21_X1  g727(.A(G141gat), .B1(new_n928), .B2(new_n668), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n922), .A2(new_n918), .ZN(new_n930));
  XNOR2_X1  g729(.A(KEYINPUT114), .B(KEYINPUT58), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n925), .A2(new_n932), .ZN(G1344gat));
  NAND3_X1  g732(.A1(new_n922), .A2(new_n481), .A3(new_n767), .ZN(new_n934));
  AOI211_X1 g733(.A(KEYINPUT59), .B(new_n481), .C1(new_n913), .C2(new_n767), .ZN(new_n935));
  XNOR2_X1  g734(.A(KEYINPUT115), .B(KEYINPUT59), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n331), .A2(new_n668), .A3(new_n333), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(KEYINPUT116), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT116), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n331), .A2(new_n939), .A3(new_n668), .A4(new_n333), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n910), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n644), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(new_n905), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n907), .B1(new_n878), .B2(new_n866), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(new_n767), .A3(new_n926), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n936), .B1(new_n946), .B2(G148gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n934), .B1(new_n935), .B2(new_n947), .ZN(G1345gat));
  OAI21_X1  g747(.A(G155gat), .B1(new_n928), .B2(new_n728), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n922), .A2(new_n203), .A3(new_n242), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1346gat));
  OAI21_X1  g750(.A(G162gat), .B1(new_n928), .B2(new_n731), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n897), .A2(G162gat), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n952), .B1(new_n921), .B2(new_n953), .ZN(G1347gat));
  NOR2_X1   g753(.A1(new_n603), .A2(new_n708), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n868), .A2(new_n587), .A3(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n957), .A2(new_n393), .A3(new_n667), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n691), .A2(new_n587), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n880), .A2(new_n667), .A3(new_n960), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n961), .A2(KEYINPUT117), .A3(G169gat), .ZN(new_n962));
  AOI21_X1  g761(.A(KEYINPUT117), .B1(new_n961), .B2(G169gat), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n958), .B1(new_n962), .B2(new_n963), .ZN(G1348gat));
  NAND2_X1  g763(.A1(new_n880), .A2(new_n960), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n767), .A2(G176gat), .ZN(new_n966));
  OAI21_X1  g765(.A(KEYINPUT118), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n394), .B1(new_n956), .B2(new_n329), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n965), .A2(KEYINPUT118), .A3(new_n966), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n969), .A2(new_n970), .ZN(G1349gat));
  NOR2_X1   g770(.A1(KEYINPUT119), .A2(KEYINPUT60), .ZN(new_n972));
  AND2_X1   g771(.A1(KEYINPUT119), .A2(KEYINPUT60), .ZN(new_n973));
  AND2_X1   g772(.A1(new_n359), .A2(new_n361), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n957), .A2(new_n974), .A3(new_n242), .ZN(new_n975));
  INV_X1    g774(.A(new_n530), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n868), .A2(new_n976), .A3(new_n242), .A4(new_n960), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(G183gat), .ZN(new_n978));
  AOI211_X1 g777(.A(new_n972), .B(new_n973), .C1(new_n975), .C2(new_n978), .ZN(new_n979));
  AND4_X1   g778(.A1(KEYINPUT119), .A2(new_n975), .A3(KEYINPUT60), .A4(new_n978), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n979), .A2(new_n980), .ZN(G1350gat));
  NOR3_X1   g780(.A1(new_n956), .A2(G190gat), .A3(new_n731), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n982), .B(KEYINPUT120), .ZN(new_n983));
  OAI21_X1  g782(.A(G190gat), .B1(new_n965), .B2(new_n731), .ZN(new_n984));
  AND2_X1   g783(.A1(new_n984), .A2(KEYINPUT61), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n984), .A2(KEYINPUT61), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n983), .B1(new_n985), .B2(new_n986), .ZN(G1351gat));
  NAND3_X1  g786(.A1(new_n680), .A2(new_n644), .A3(new_n691), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n988), .A2(KEYINPUT121), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT121), .ZN(new_n990));
  NAND4_X1  g789(.A1(new_n680), .A2(new_n990), .A3(new_n644), .A4(new_n691), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND4_X1  g791(.A1(new_n868), .A2(KEYINPUT122), .A3(new_n587), .A4(new_n992), .ZN(new_n993));
  OAI211_X1 g792(.A(new_n587), .B(new_n992), .C1(new_n878), .C2(new_n866), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT122), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g796(.A(G197gat), .B1(new_n997), .B2(new_n667), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n960), .A2(new_n680), .ZN(new_n999));
  AOI21_X1  g798(.A(new_n908), .B1(new_n865), .B2(new_n867), .ZN(new_n1000));
  AOI21_X1  g799(.A(KEYINPUT57), .B1(new_n941), .B2(new_n644), .ZN(new_n1001));
  OAI21_X1  g800(.A(KEYINPUT123), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g801(.A(KEYINPUT123), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n943), .A2(new_n944), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g803(.A(new_n999), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  AND2_X1   g804(.A1(new_n667), .A2(G197gat), .ZN(new_n1006));
  AOI21_X1  g805(.A(new_n998), .B1(new_n1005), .B2(new_n1006), .ZN(G1352gat));
  INV_X1    g806(.A(new_n994), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT62), .ZN(new_n1009));
  NOR2_X1   g808(.A1(new_n1009), .A2(KEYINPUT124), .ZN(new_n1010));
  NOR2_X1   g809(.A1(new_n329), .A2(G204gat), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n1008), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g811(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n1013));
  INV_X1    g812(.A(new_n1011), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n1013), .B1(new_n994), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g815(.A(new_n999), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1017), .A2(new_n767), .ZN(new_n1018));
  AOI21_X1  g817(.A(new_n1018), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1019));
  OAI21_X1  g818(.A(new_n1016), .B1(new_n1019), .B2(new_n457), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1020), .A2(KEYINPUT125), .ZN(new_n1021));
  INV_X1    g820(.A(KEYINPUT125), .ZN(new_n1022));
  OAI211_X1 g821(.A(new_n1022), .B(new_n1016), .C1(new_n1019), .C2(new_n457), .ZN(new_n1023));
  NAND2_X1  g822(.A1(new_n1021), .A2(new_n1023), .ZN(G1353gat));
  NAND3_X1  g823(.A1(new_n997), .A2(new_n465), .A3(new_n242), .ZN(new_n1025));
  NAND2_X1  g824(.A1(new_n1017), .A2(new_n242), .ZN(new_n1026));
  AOI21_X1  g825(.A(new_n1026), .B1(new_n943), .B2(new_n944), .ZN(new_n1027));
  INV_X1    g826(.A(KEYINPUT126), .ZN(new_n1028));
  AOI21_X1  g827(.A(new_n448), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g828(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1030));
  OAI21_X1  g829(.A(KEYINPUT126), .B1(new_n1030), .B2(new_n1026), .ZN(new_n1031));
  AND3_X1   g830(.A1(new_n1029), .A2(new_n1031), .A3(KEYINPUT63), .ZN(new_n1032));
  AOI21_X1  g831(.A(KEYINPUT63), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1033));
  OAI21_X1  g832(.A(new_n1025), .B1(new_n1032), .B2(new_n1033), .ZN(G1354gat));
  INV_X1    g833(.A(KEYINPUT127), .ZN(new_n1035));
  NOR2_X1   g834(.A1(new_n731), .A2(new_n466), .ZN(new_n1036));
  INV_X1    g835(.A(new_n1036), .ZN(new_n1037));
  AOI211_X1 g836(.A(new_n999), .B(new_n1037), .C1(new_n1002), .C2(new_n1004), .ZN(new_n1038));
  AOI21_X1  g837(.A(G218gat), .B1(new_n997), .B2(new_n730), .ZN(new_n1039));
  OAI21_X1  g838(.A(new_n1035), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g839(.A(new_n1004), .ZN(new_n1041));
  AOI21_X1  g840(.A(new_n1003), .B1(new_n943), .B2(new_n944), .ZN(new_n1042));
  OAI211_X1 g841(.A(new_n1017), .B(new_n1036), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g842(.A(new_n731), .B1(new_n993), .B2(new_n996), .ZN(new_n1044));
  OAI211_X1 g843(.A(new_n1043), .B(KEYINPUT127), .C1(G218gat), .C2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g844(.A1(new_n1040), .A2(new_n1045), .ZN(G1355gat));
endmodule


