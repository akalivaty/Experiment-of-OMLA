//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 1 0 0 1 1 0 0 0 0 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n552, new_n553, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n566, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n604,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1168;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(new_n454));
  OR2_X1    g029(.A1(new_n452), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT68), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G101), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n463), .A2(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n467), .A2(new_n470), .ZN(G160));
  NAND2_X1  g046(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n477), .B(new_n478), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n481));
  OR2_X1    g056(.A1(new_n481), .A2(KEYINPUT70), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(KEYINPUT70), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n475), .A2(new_n464), .ZN(new_n484));
  AOI22_X1  g059(.A1(new_n482), .A2(new_n483), .B1(G124), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  OR2_X1    g062(.A1(new_n464), .A2(G114), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AOI22_X1  g065(.A1(new_n484), .A2(G126), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n472), .A2(new_n474), .A3(G138), .A4(new_n464), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n463), .A2(new_n494), .A3(G138), .A4(new_n464), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  INV_X1    g073(.A(G651), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT6), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G651), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n500), .A2(new_n502), .A3(G50), .A4(G543), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n505), .A2(new_n507), .A3(new_n500), .A4(new_n502), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT71), .B(G88), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n503), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT72), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n512));
  OAI211_X1 g087(.A(new_n512), .B(new_n503), .C1(new_n508), .C2(new_n509), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT5), .B(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G62), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n499), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(G166));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  INV_X1    g098(.A(G89), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n524), .B2(new_n508), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT73), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n500), .A2(new_n502), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n504), .ZN(new_n528));
  AND2_X1   g103(.A1(G63), .A2(G651), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n528), .A2(G51), .B1(new_n515), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n531), .B(new_n532), .ZN(G168));
  AND2_X1   g108(.A1(new_n500), .A2(new_n502), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n535), .A2(new_n536), .B1(new_n537), .B2(new_n508), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n499), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n538), .A2(new_n540), .ZN(G171));
  INV_X1    g116(.A(G43), .ZN(new_n542));
  INV_X1    g117(.A(G81), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n535), .A2(new_n542), .B1(new_n543), .B2(new_n508), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n499), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(new_n528), .A2(G53), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT9), .ZN(new_n556));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n505), .A2(new_n507), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n508), .ZN(new_n561));
  AOI22_X1  g136(.A1(G651), .A2(new_n560), .B1(new_n561), .B2(G91), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n556), .A2(new_n562), .ZN(G299));
  INV_X1    g138(.A(G171), .ZN(G301));
  XNOR2_X1  g139(.A(new_n531), .B(KEYINPUT74), .ZN(G286));
  INV_X1    g140(.A(KEYINPUT75), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n566), .B1(new_n514), .B2(new_n519), .ZN(new_n567));
  AOI211_X1 g142(.A(KEYINPUT75), .B(new_n518), .C1(new_n511), .C2(new_n513), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n567), .A2(new_n568), .ZN(G303));
  NAND2_X1  g144(.A1(new_n561), .A2(G87), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n528), .A2(G49), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(KEYINPUT76), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(G288));
  NAND3_X1  g153(.A1(new_n534), .A2(G86), .A3(new_n515), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n500), .A2(new_n502), .A3(G48), .A4(G543), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n515), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(new_n499), .ZN(G305));
  XNOR2_X1  g157(.A(KEYINPUT77), .B(G47), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n561), .A2(G85), .B1(new_n528), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n499), .B2(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(G301), .A2(G868), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n561), .A2(KEYINPUT10), .A3(G92), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT10), .ZN(new_n589));
  INV_X1    g164(.A(G92), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n508), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n588), .A2(new_n591), .B1(G54), .B2(new_n528), .ZN(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n558), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n499), .B1(new_n595), .B2(KEYINPUT78), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n596), .B1(KEYINPUT78), .B2(new_n595), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n587), .B1(new_n599), .B2(G868), .ZN(G284));
  OAI21_X1  g175(.A(new_n587), .B1(new_n599), .B2(G868), .ZN(G321));
  MUX2_X1   g176(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g177(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n599), .B1(new_n604), .B2(G860), .ZN(G148));
  NAND2_X1  g180(.A1(new_n599), .A2(new_n604), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G868), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g184(.A1(new_n463), .A2(new_n461), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT12), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(KEYINPUT13), .Z(new_n612));
  OR2_X1    g187(.A1(new_n612), .A2(G2100), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n476), .A2(G135), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n484), .A2(G123), .ZN(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n616));
  INV_X1    g191(.A(G111), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n616), .A2(KEYINPUT79), .B1(new_n617), .B2(G2105), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(KEYINPUT79), .B2(new_n616), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n614), .A2(new_n615), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(G2096), .Z(new_n621));
  NAND2_X1  g196(.A1(new_n612), .A2(G2100), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n613), .A2(new_n621), .A3(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2435), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT81), .B(G2438), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n624), .B(new_n625), .Z(new_n626));
  XNOR2_X1  g201(.A(G2427), .B(G2430), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n624), .B(new_n625), .ZN(new_n629));
  INV_X1    g204(.A(new_n627), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n628), .A2(KEYINPUT14), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n632), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(G14), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n641), .B1(new_n638), .B2(new_n639), .ZN(new_n642));
  AND2_X1   g217(.A1(new_n640), .A2(new_n642), .ZN(G401));
  XOR2_X1   g218(.A(G2072), .B(G2078), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT82), .ZN(new_n645));
  XOR2_X1   g220(.A(G2067), .B(G2678), .Z(new_n646));
  XNOR2_X1  g221(.A(G2084), .B(G2090), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT18), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT17), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n646), .B2(new_n647), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n645), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n648), .B1(new_n645), .B2(new_n652), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n650), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2096), .B(G2100), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT83), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n655), .B(new_n657), .ZN(G227));
  XNOR2_X1  g233(.A(G1981), .B(G1986), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1971), .B(G1976), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1956), .B(G2474), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1961), .B(G1966), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n662), .A2(KEYINPUT20), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n663), .B(new_n664), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n666), .B(new_n667), .C1(new_n662), .C2(new_n668), .ZN(new_n669));
  AOI21_X1  g244(.A(KEYINPUT20), .B1(new_n662), .B2(new_n665), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(G1991), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n669), .A2(G1991), .A3(new_n670), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(G1996), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n675), .A2(G1996), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n659), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n678), .ZN(new_n680));
  INV_X1    g255(.A(new_n659), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n680), .A2(new_n681), .A3(new_n676), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n679), .A2(new_n682), .A3(new_n684), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(G229));
  XNOR2_X1  g263(.A(KEYINPUT92), .B(KEYINPUT93), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT25), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n461), .A2(G103), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n690), .B(new_n691), .Z(new_n692));
  NAND2_X1  g267(.A1(new_n476), .A2(G139), .ZN(new_n693));
  AOI22_X1  g268(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n692), .B(new_n693), .C1(new_n464), .C2(new_n694), .ZN(new_n695));
  MUX2_X1   g270(.A(G33), .B(new_n695), .S(G29), .Z(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(G2072), .Z(new_n697));
  NOR2_X1   g272(.A1(G29), .A2(G32), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n484), .A2(G129), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n476), .A2(G141), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n461), .A2(G105), .ZN(new_n701));
  NAND3_X1  g276(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT26), .Z(new_n703));
  NAND4_X1  g278(.A1(new_n699), .A2(new_n700), .A3(new_n701), .A4(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n698), .B1(new_n705), .B2(G29), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT27), .B(G1996), .Z(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT31), .B(G11), .ZN(new_n709));
  INV_X1    g284(.A(G28), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n710), .A2(KEYINPUT30), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT30), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(G28), .ZN(new_n714));
  OAI221_X1 g289(.A(new_n709), .B1(new_n711), .B2(new_n714), .C1(new_n620), .C2(new_n712), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n708), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G1961), .ZN(new_n717));
  NAND2_X1  g292(.A1(G171), .A2(G16), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G5), .B2(G16), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n697), .B(new_n716), .C1(new_n717), .C2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n712), .A2(G35), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G162), .B2(new_n712), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT29), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n723), .A2(G2090), .ZN(new_n724));
  NOR2_X1   g299(.A1(G4), .A2(G16), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n599), .B2(G16), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G1348), .ZN(new_n727));
  AND2_X1   g302(.A1(KEYINPUT87), .A2(G16), .ZN(new_n728));
  NOR2_X1   g303(.A1(KEYINPUT87), .A2(G16), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n548), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G19), .B2(new_n731), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n733), .A2(G1341), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(G1341), .ZN(new_n735));
  INV_X1    g310(.A(G2078), .ZN(new_n736));
  NOR2_X1   g311(.A1(G164), .A2(new_n712), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G27), .B2(new_n712), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n734), .A2(new_n735), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n736), .B2(new_n738), .ZN(new_n740));
  NOR4_X1   g315(.A1(new_n720), .A2(new_n724), .A3(new_n727), .A4(new_n740), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n719), .A2(new_n717), .B1(new_n706), .B2(new_n707), .ZN(new_n742));
  INV_X1    g317(.A(G34), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n743), .A2(KEYINPUT24), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(KEYINPUT24), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n712), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G160), .B2(new_n712), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT94), .Z(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n742), .B1(new_n749), .B2(G2084), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n750), .A2(KEYINPUT95), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n750), .A2(KEYINPUT95), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n712), .A2(G26), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT28), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n484), .A2(G128), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n476), .A2(G140), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n464), .A2(G116), .ZN(new_n757));
  OAI21_X1  g332(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n755), .B(new_n756), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G29), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n760), .A2(KEYINPUT90), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n760), .A2(KEYINPUT90), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n754), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT91), .B(G2067), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  INV_X1    g341(.A(G2084), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n765), .B(new_n766), .C1(new_n767), .C2(new_n748), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n751), .A2(new_n752), .A3(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G16), .A2(G21), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G168), .B2(G16), .ZN(new_n771));
  INV_X1    g346(.A(G1966), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n723), .A2(G2090), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n731), .A2(G20), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT23), .Z(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G299), .B2(G16), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1956), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT96), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n741), .A2(new_n769), .A3(new_n773), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n731), .A2(G22), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G166), .B2(new_n731), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n783), .A2(G1971), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(G1971), .ZN(new_n785));
  MUX2_X1   g360(.A(G6), .B(G305), .S(G16), .Z(new_n786));
  XOR2_X1   g361(.A(KEYINPUT32), .B(G1981), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(G16), .A2(G23), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n574), .B2(G16), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT33), .B(G1976), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n784), .A2(new_n785), .A3(new_n788), .A4(new_n792), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT89), .Z(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT88), .B(KEYINPUT34), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  MUX2_X1   g372(.A(G24), .B(G290), .S(new_n730), .Z(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(G1986), .Z(new_n799));
  NOR2_X1   g374(.A1(G25), .A2(G29), .ZN(new_n800));
  AOI22_X1  g375(.A1(G119), .A2(new_n484), .B1(new_n476), .B2(G131), .ZN(new_n801));
  OAI21_X1  g376(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n802));
  INV_X1    g377(.A(G107), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(G2105), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT85), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT86), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n800), .B1(new_n807), .B2(G29), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT35), .B(G1991), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n808), .B(new_n810), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n796), .A2(new_n797), .A3(new_n799), .A4(new_n811), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n812), .A2(KEYINPUT36), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(KEYINPUT36), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n781), .B1(new_n813), .B2(new_n814), .ZN(G311));
  XNOR2_X1  g390(.A(new_n812), .B(KEYINPUT36), .ZN(new_n816));
  AND3_X1   g391(.A1(new_n741), .A2(new_n773), .A3(new_n780), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n816), .A2(new_n769), .A3(new_n817), .ZN(G150));
  NOR2_X1   g393(.A1(new_n598), .A2(new_n604), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT97), .B(G55), .ZN(new_n822));
  INV_X1    g397(.A(G93), .ZN(new_n823));
  OAI22_X1  g398(.A1(new_n535), .A2(new_n822), .B1(new_n823), .B2(new_n508), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(new_n499), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n547), .B(new_n827), .Z(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(G860), .B1(new_n821), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n829), .B2(new_n821), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n827), .A2(G860), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT37), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(G145));
  XNOR2_X1  g409(.A(new_n620), .B(KEYINPUT98), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(new_n806), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n486), .B(G160), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n836), .B(new_n837), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n704), .B(new_n611), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n836), .B(new_n837), .ZN(new_n841));
  INV_X1    g416(.A(new_n839), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n496), .A2(KEYINPUT99), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT99), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n493), .A2(new_n495), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n845), .A2(new_n491), .A3(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n759), .ZN(new_n849));
  AOI22_X1  g424(.A1(G130), .A2(new_n484), .B1(new_n476), .B2(G142), .ZN(new_n850));
  OAI21_X1  g425(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n851));
  INV_X1    g426(.A(G118), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n851), .A2(KEYINPUT100), .B1(new_n852), .B2(G2105), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(KEYINPUT100), .B2(new_n851), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n849), .B(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n695), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n844), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(G37), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n840), .A2(new_n857), .A3(new_n843), .ZN(new_n861));
  AND4_X1   g436(.A1(KEYINPUT101), .A2(new_n859), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(G37), .B1(new_n844), .B2(new_n858), .ZN(new_n863));
  AOI21_X1  g438(.A(KEYINPUT101), .B1(new_n863), .B2(new_n861), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT40), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(G395));
  INV_X1    g442(.A(new_n827), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n868), .A2(G868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n828), .B(new_n606), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n599), .B(G299), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(KEYINPUT41), .B2(new_n873), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n874), .B1(new_n871), .B2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n520), .B(new_n573), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n515), .A2(G61), .ZN(new_n880));
  NAND2_X1  g455(.A1(G73), .A2(G543), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n499), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(G86), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n580), .B1(new_n508), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(G290), .B(new_n885), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n879), .B(new_n886), .Z(new_n887));
  XNOR2_X1  g462(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n878), .B(new_n889), .Z(new_n890));
  INV_X1    g465(.A(G868), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n870), .B1(new_n890), .B2(new_n891), .ZN(G295));
  INV_X1    g467(.A(KEYINPUT104), .ZN(new_n893));
  XNOR2_X1  g468(.A(G295), .B(new_n893), .ZN(G331));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n895));
  NAND2_X1  g470(.A1(G286), .A2(G301), .ZN(new_n896));
  NAND2_X1  g471(.A1(G168), .A2(G171), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n828), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n896), .A2(new_n897), .A3(new_n829), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n873), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n872), .A2(KEYINPUT41), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n903), .B1(new_n872), .B2(new_n875), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n899), .A2(new_n904), .A3(new_n900), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n901), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n905), .A2(new_n902), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n887), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n899), .A2(new_n900), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n872), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n877), .A2(new_n899), .A3(new_n900), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(new_n887), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n860), .ZN(new_n913));
  NOR3_X1   g488(.A1(new_n908), .A2(new_n913), .A3(KEYINPUT43), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n912), .A2(new_n860), .ZN(new_n916));
  INV_X1    g491(.A(new_n887), .ZN(new_n917));
  INV_X1    g492(.A(new_n911), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n917), .B1(new_n918), .B2(new_n901), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n915), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n895), .B1(new_n914), .B2(new_n920), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n916), .A2(KEYINPUT106), .A3(new_n915), .A4(new_n919), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT43), .B1(new_n908), .B2(new_n913), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n919), .A2(new_n912), .A3(new_n915), .A4(new_n860), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n922), .A2(new_n923), .A3(new_n926), .A4(KEYINPUT44), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n921), .A2(new_n927), .ZN(G397));
  NAND2_X1  g503(.A1(new_n488), .A2(new_n490), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n463), .A2(G2105), .ZN(new_n930));
  INV_X1    g505(.A(G126), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n932), .B1(new_n496), .B2(KEYINPUT99), .ZN(new_n933));
  AOI21_X1  g508(.A(G1384), .B1(new_n933), .B2(new_n847), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n468), .A2(new_n469), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(G2105), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n476), .A2(G137), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n936), .A2(new_n937), .A3(G40), .A4(new_n462), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n934), .A2(KEYINPUT45), .A3(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n759), .B(G2067), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n704), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XOR2_X1   g518(.A(new_n943), .B(KEYINPUT126), .Z(new_n944));
  INV_X1    g519(.A(G1996), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n939), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(KEYINPUT46), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT47), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n939), .A2(new_n945), .A3(new_n705), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n950), .A2(new_n951), .ZN(new_n953));
  OAI221_X1 g528(.A(new_n941), .B1(new_n945), .B2(new_n942), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT108), .ZN(new_n955));
  OR2_X1    g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n955), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n806), .B(new_n809), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n939), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n956), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(G290), .A2(G1986), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n939), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g537(.A(new_n962), .B(KEYINPUT48), .Z(new_n963));
  OAI21_X1  g538(.A(new_n949), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n956), .A2(new_n810), .A3(new_n807), .A4(new_n957), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(G2067), .B2(new_n759), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n964), .B1(new_n939), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT113), .ZN(new_n968));
  XNOR2_X1  g543(.A(KEYINPUT112), .B(G1981), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n968), .B1(G305), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n969), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n885), .A2(KEYINPUT113), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(G305), .A2(G1981), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT49), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G8), .ZN(new_n978));
  INV_X1    g553(.A(G40), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n467), .A2(new_n470), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n978), .B1(new_n934), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n973), .A2(KEYINPUT49), .A3(new_n974), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n977), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G1976), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT52), .B1(G288), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n574), .A2(G1976), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n985), .A2(new_n981), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1384), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n848), .A2(new_n988), .A3(new_n980), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n989), .A2(G8), .A3(new_n986), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n990), .A2(new_n991), .A3(KEYINPUT52), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n991), .B1(new_n990), .B2(KEYINPUT52), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n983), .B(new_n987), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G1971), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n996));
  AOI211_X1 g571(.A(new_n996), .B(G1384), .C1(new_n933), .C2(new_n847), .ZN(new_n997));
  AOI21_X1  g572(.A(G1384), .B1(new_n491), .B2(new_n496), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n980), .B1(new_n998), .B2(KEYINPUT45), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n995), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT50), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n938), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G2090), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n1002), .B(new_n1003), .C1(new_n934), .C2(new_n1001), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n978), .B1(new_n1000), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(G8), .B1(new_n567), .B2(new_n568), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI211_X1 g583(.A(KEYINPUT55), .B(G8), .C1(new_n567), .C2(new_n568), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1005), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n994), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n848), .A2(new_n1001), .A3(new_n988), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT109), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n848), .A2(KEYINPUT109), .A3(new_n1001), .A4(new_n988), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n980), .B1(new_n998), .B2(new_n1001), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1015), .A2(new_n1003), .A3(new_n1016), .A4(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT110), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1017), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1021), .A2(new_n1022), .A3(new_n1003), .A4(new_n1016), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1020), .A2(new_n1023), .A3(new_n1000), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1024), .A2(G8), .A3(new_n1010), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n980), .B1(new_n934), .B2(KEYINPUT45), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n988), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT117), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n998), .A2(new_n1029), .A3(KEYINPUT45), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n772), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1021), .A2(new_n767), .A3(new_n1016), .ZN(new_n1033));
  AOI211_X1 g608(.A(new_n978), .B(G286), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1012), .A2(new_n1025), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT63), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT118), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1035), .A2(new_n1039), .A3(new_n1036), .ZN(new_n1040));
  XNOR2_X1  g615(.A(new_n994), .B(KEYINPUT114), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1034), .A2(KEYINPUT63), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1024), .A2(G8), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1043), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1041), .A2(new_n1042), .A3(new_n1025), .A4(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1038), .A2(new_n1040), .A3(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n575), .A2(new_n984), .A3(new_n577), .ZN(new_n1047));
  XOR2_X1   g622(.A(new_n1047), .B(KEYINPUT115), .Z(new_n1048));
  AOI22_X1  g623(.A1(new_n1048), .A2(new_n983), .B1(new_n970), .B2(new_n972), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1049), .A2(KEYINPUT116), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1049), .A2(KEYINPUT116), .ZN(new_n1051));
  INV_X1    g626(.A(new_n981), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1025), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1053), .B1(new_n1054), .B2(new_n1041), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1046), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1033), .A2(new_n1032), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1057), .B(G8), .C1(new_n1058), .C2(G286), .ZN(new_n1059));
  NOR2_X1   g634(.A1(G168), .A2(new_n978), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n978), .B1(new_n1033), .B2(new_n1032), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n1063), .A2(new_n1060), .A3(new_n1057), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT125), .ZN(new_n1065));
  OAI22_X1  g640(.A1(new_n1062), .A2(new_n1064), .B1(new_n1065), .B2(KEYINPUT62), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(KEYINPUT62), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n1026), .A2(new_n1069), .A3(G2078), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1070), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n934), .A2(KEYINPUT45), .ZN(new_n1072));
  INV_X1    g647(.A(new_n999), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1072), .A2(new_n1073), .A3(new_n736), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n1069), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1071), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(G1961), .B1(new_n1021), .B2(new_n1016), .ZN(new_n1077));
  OAI21_X1  g652(.A(G171), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1065), .B(KEYINPUT62), .C1(new_n1062), .C2(new_n1064), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1068), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1070), .A2(new_n1072), .B1(new_n1069), .B2(new_n1074), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1021), .A2(new_n1016), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1083), .A2(KEYINPUT123), .A3(new_n717), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1077), .A2(KEYINPUT123), .ZN(new_n1085));
  OAI211_X1 g660(.A(G301), .B(new_n1082), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT54), .B1(new_n1078), .B2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1082), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT124), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(KEYINPUT124), .B(new_n1082), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1092), .A2(G171), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1095), .B1(new_n1096), .B2(G301), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1089), .A2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT56), .B(G2072), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1072), .A2(new_n1073), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n848), .A2(new_n988), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT50), .ZN(new_n1104));
  AOI21_X1  g679(.A(G1956), .B1(new_n1104), .B2(new_n1002), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1107), .A2(KEYINPUT119), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(KEYINPUT119), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT9), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n555), .B(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n562), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1108), .B(new_n1109), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n556), .A2(KEYINPUT119), .A3(new_n1107), .A4(new_n562), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1106), .A2(KEYINPUT120), .A3(new_n1116), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1104), .A2(new_n1002), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1116), .B(new_n1101), .C1(new_n1118), .C2(G1956), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT120), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(G1348), .ZN(new_n1123));
  INV_X1    g698(.A(G2067), .ZN(new_n1124));
  INV_X1    g699(.A(new_n989), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1083), .A2(new_n1123), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  OR2_X1    g701(.A1(new_n1126), .A2(new_n598), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1115), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1122), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1083), .A2(new_n1123), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1125), .A2(new_n1124), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1130), .A2(KEYINPUT60), .A3(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1132), .A2(KEYINPUT122), .A3(new_n599), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1126), .A2(KEYINPUT60), .A3(new_n598), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(KEYINPUT122), .B1(new_n1132), .B2(new_n599), .ZN(new_n1136));
  OAI22_X1  g711(.A1(new_n1135), .A2(new_n1136), .B1(KEYINPUT60), .B2(new_n1126), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1128), .A2(new_n1119), .A3(KEYINPUT61), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1072), .A2(new_n945), .A3(new_n1073), .ZN(new_n1139));
  XNOR2_X1  g714(.A(KEYINPUT58), .B(G1341), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1139), .B1(new_n1125), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n548), .ZN(new_n1142));
  NOR2_X1   g717(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  XOR2_X1   g719(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1145));
  NAND3_X1  g720(.A1(new_n1141), .A2(new_n548), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1138), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT61), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1117), .A2(new_n1121), .A3(new_n1128), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1129), .B1(new_n1137), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1081), .B1(new_n1099), .B2(new_n1151), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1012), .A2(new_n1025), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1056), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  AND2_X1   g729(.A1(G290), .A2(G1986), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n939), .B1(new_n961), .B2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n956), .A2(new_n1156), .A3(new_n957), .A4(new_n959), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n967), .B1(new_n1154), .B2(new_n1157), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g733(.A1(new_n914), .A2(new_n920), .ZN(new_n1160));
  AOI211_X1 g734(.A(new_n458), .B(G227), .C1(new_n640), .C2(new_n642), .ZN(new_n1161));
  NAND3_X1  g735(.A1(new_n1161), .A2(new_n686), .A3(new_n687), .ZN(new_n1162));
  NAND2_X1  g736(.A1(new_n1162), .A2(KEYINPUT127), .ZN(new_n1163));
  INV_X1    g737(.A(KEYINPUT127), .ZN(new_n1164));
  NAND4_X1  g738(.A1(new_n1161), .A2(new_n686), .A3(new_n1164), .A4(new_n687), .ZN(new_n1165));
  OAI211_X1 g739(.A(new_n1163), .B(new_n1165), .C1(new_n862), .C2(new_n864), .ZN(new_n1166));
  NOR2_X1   g740(.A1(new_n1160), .A2(new_n1166), .ZN(G308));
  AND2_X1   g741(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1168));
  OAI221_X1 g742(.A(new_n1168), .B1(new_n864), .B2(new_n862), .C1(new_n920), .C2(new_n914), .ZN(G225));
endmodule


