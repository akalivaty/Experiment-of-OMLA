

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584;

  NOR2_X1 U322 ( .A1(n533), .A2(n463), .ZN(n413) );
  XNOR2_X1 U323 ( .A(n360), .B(n359), .ZN(n361) );
  INV_X1 U324 ( .A(n406), .ZN(n359) );
  XNOR2_X1 U325 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U326 ( .A(n446), .B(KEYINPUT123), .ZN(n581) );
  XNOR2_X1 U327 ( .A(n368), .B(n367), .ZN(n577) );
  XOR2_X1 U328 ( .A(G134GAT), .B(G106GAT), .Z(n290) );
  XNOR2_X1 U329 ( .A(n460), .B(KEYINPUT90), .ZN(n461) );
  NOR2_X1 U330 ( .A1(n562), .A2(n387), .ZN(n388) );
  INV_X1 U331 ( .A(KEYINPUT54), .ZN(n412) );
  XNOR2_X1 U332 ( .A(n373), .B(n290), .ZN(n378) );
  NOR2_X1 U333 ( .A1(n475), .A2(n474), .ZN(n476) );
  XNOR2_X1 U334 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U335 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U336 ( .A(n430), .B(n429), .ZN(n466) );
  INV_X1 U337 ( .A(G204GAT), .ZN(n447) );
  NOR2_X1 U338 ( .A1(n464), .A2(n453), .ZN(n569) );
  XNOR2_X1 U339 ( .A(n495), .B(KEYINPUT38), .ZN(n504) );
  XNOR2_X1 U340 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U341 ( .A(n450), .B(n449), .ZN(G1353GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n292) );
  NAND2_X1 U343 ( .A1(G230GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U344 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U345 ( .A(n293), .B(KEYINPUT32), .Z(n302) );
  INV_X1 U346 ( .A(KEYINPUT71), .ZN(n294) );
  NAND2_X1 U347 ( .A1(KEYINPUT13), .A2(n294), .ZN(n297) );
  INV_X1 U348 ( .A(KEYINPUT13), .ZN(n295) );
  NAND2_X1 U349 ( .A1(n295), .A2(KEYINPUT71), .ZN(n296) );
  NAND2_X1 U350 ( .A1(n297), .A2(n296), .ZN(n299) );
  XNOR2_X1 U351 ( .A(G71GAT), .B(G57GAT), .ZN(n298) );
  XNOR2_X1 U352 ( .A(n299), .B(n298), .ZN(n355) );
  XNOR2_X1 U353 ( .A(G176GAT), .B(G92GAT), .ZN(n300) );
  XNOR2_X1 U354 ( .A(n300), .B(G64GAT), .ZN(n404) );
  XNOR2_X1 U355 ( .A(n355), .B(n404), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U357 ( .A(KEYINPUT72), .B(KEYINPUT75), .Z(n304) );
  XNOR2_X1 U358 ( .A(G120GAT), .B(G204GAT), .ZN(n303) );
  XNOR2_X1 U359 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U360 ( .A(n306), .B(n305), .Z(n311) );
  XOR2_X1 U361 ( .A(G78GAT), .B(G148GAT), .Z(n308) );
  XNOR2_X1 U362 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n307) );
  XNOR2_X1 U363 ( .A(n308), .B(n307), .ZN(n427) );
  XNOR2_X1 U364 ( .A(G99GAT), .B(G85GAT), .ZN(n309) );
  XNOR2_X1 U365 ( .A(n309), .B(KEYINPUT74), .ZN(n374) );
  XNOR2_X1 U366 ( .A(n427), .B(n374), .ZN(n310) );
  XNOR2_X1 U367 ( .A(n311), .B(n310), .ZN(n458) );
  XOR2_X1 U368 ( .A(KEYINPUT89), .B(KEYINPUT4), .Z(n313) );
  XNOR2_X1 U369 ( .A(KEYINPUT87), .B(KEYINPUT5), .ZN(n312) );
  XNOR2_X1 U370 ( .A(n313), .B(n312), .ZN(n318) );
  XNOR2_X1 U371 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n314) );
  XNOR2_X1 U372 ( .A(n314), .B(KEYINPUT2), .ZN(n425) );
  XOR2_X1 U373 ( .A(n425), .B(G1GAT), .Z(n316) );
  NAND2_X1 U374 ( .A1(G225GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U375 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U376 ( .A(n318), .B(n317), .ZN(n333) );
  XOR2_X1 U377 ( .A(KEYINPUT85), .B(KEYINPUT6), .Z(n320) );
  XNOR2_X1 U378 ( .A(G127GAT), .B(G155GAT), .ZN(n319) );
  XNOR2_X1 U379 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U380 ( .A(KEYINPUT86), .B(KEYINPUT88), .Z(n322) );
  XNOR2_X1 U381 ( .A(KEYINPUT1), .B(G57GAT), .ZN(n321) );
  XNOR2_X1 U382 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U383 ( .A(n324), .B(n323), .Z(n331) );
  XOR2_X1 U384 ( .A(G120GAT), .B(KEYINPUT0), .Z(n326) );
  XNOR2_X1 U385 ( .A(G113GAT), .B(G134GAT), .ZN(n325) );
  XNOR2_X1 U386 ( .A(n326), .B(n325), .ZN(n438) );
  XOR2_X1 U387 ( .A(G85GAT), .B(G162GAT), .Z(n328) );
  XNOR2_X1 U388 ( .A(G29GAT), .B(G148GAT), .ZN(n327) );
  XNOR2_X1 U389 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U390 ( .A(n438), .B(n329), .ZN(n330) );
  XNOR2_X1 U391 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U392 ( .A(n333), .B(n332), .ZN(n521) );
  XOR2_X1 U393 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n335) );
  XNOR2_X1 U394 ( .A(G43GAT), .B(G29GAT), .ZN(n334) );
  XNOR2_X1 U395 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U396 ( .A(KEYINPUT69), .B(n336), .ZN(n382) );
  XOR2_X1 U397 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n338) );
  XNOR2_X1 U398 ( .A(G8GAT), .B(KEYINPUT68), .ZN(n337) );
  XNOR2_X1 U399 ( .A(n338), .B(n337), .ZN(n351) );
  XOR2_X1 U400 ( .A(G141GAT), .B(G197GAT), .Z(n340) );
  XNOR2_X1 U401 ( .A(G36GAT), .B(G50GAT), .ZN(n339) );
  XNOR2_X1 U402 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U403 ( .A(G15GAT), .B(G113GAT), .Z(n342) );
  XNOR2_X1 U404 ( .A(G169GAT), .B(G22GAT), .ZN(n341) );
  XNOR2_X1 U405 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U406 ( .A(n344), .B(n343), .Z(n349) );
  XOR2_X1 U407 ( .A(G1GAT), .B(KEYINPUT70), .Z(n364) );
  XOR2_X1 U408 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n346) );
  NAND2_X1 U409 ( .A1(G229GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U410 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U411 ( .A(n364), .B(n347), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U413 ( .A(n351), .B(n350), .Z(n352) );
  XNOR2_X1 U414 ( .A(n382), .B(n352), .ZN(n572) );
  INV_X1 U415 ( .A(n572), .ZN(n562) );
  XOR2_X1 U416 ( .A(KEYINPUT79), .B(KEYINPUT12), .Z(n354) );
  XNOR2_X1 U417 ( .A(KEYINPUT14), .B(KEYINPUT78), .ZN(n353) );
  XNOR2_X1 U418 ( .A(n354), .B(n353), .ZN(n368) );
  XNOR2_X1 U419 ( .A(n355), .B(KEYINPUT15), .ZN(n357) );
  AND2_X1 U420 ( .A1(G231GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U421 ( .A(n357), .B(n356), .ZN(n362) );
  XOR2_X1 U422 ( .A(G15GAT), .B(G127GAT), .Z(n442) );
  XOR2_X1 U423 ( .A(G22GAT), .B(G155GAT), .Z(n419) );
  XNOR2_X1 U424 ( .A(n442), .B(n419), .ZN(n360) );
  XNOR2_X1 U425 ( .A(G8GAT), .B(G183GAT), .ZN(n358) );
  XNOR2_X1 U426 ( .A(n358), .B(G211GAT), .ZN(n406) );
  XNOR2_X1 U427 ( .A(n363), .B(G64GAT), .ZN(n366) );
  XOR2_X1 U428 ( .A(n364), .B(G78GAT), .Z(n365) );
  XNOR2_X1 U429 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U430 ( .A(KEYINPUT11), .B(KEYINPUT65), .Z(n370) );
  XNOR2_X1 U431 ( .A(G92GAT), .B(KEYINPUT10), .ZN(n369) );
  XOR2_X1 U432 ( .A(n370), .B(n369), .Z(n380) );
  XOR2_X1 U433 ( .A(G36GAT), .B(G190GAT), .Z(n405) );
  XOR2_X1 U434 ( .A(KEYINPUT9), .B(n405), .Z(n372) );
  XOR2_X1 U435 ( .A(G50GAT), .B(G162GAT), .Z(n418) );
  XNOR2_X1 U436 ( .A(G218GAT), .B(n418), .ZN(n371) );
  XNOR2_X1 U437 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U438 ( .A(n374), .B(KEYINPUT77), .ZN(n376) );
  AND2_X1 U439 ( .A1(G232GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U440 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U441 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n382), .B(n381), .ZN(n392) );
  XNOR2_X1 U443 ( .A(n392), .B(KEYINPUT36), .ZN(n582) );
  NOR2_X1 U444 ( .A1(n577), .A2(n582), .ZN(n384) );
  XNOR2_X1 U445 ( .A(KEYINPUT45), .B(KEYINPUT112), .ZN(n383) );
  XNOR2_X1 U446 ( .A(n384), .B(n383), .ZN(n385) );
  NAND2_X1 U447 ( .A1(n385), .A2(n458), .ZN(n386) );
  XOR2_X1 U448 ( .A(KEYINPUT113), .B(n386), .Z(n387) );
  XNOR2_X1 U449 ( .A(n388), .B(KEYINPUT114), .ZN(n397) );
  XOR2_X1 U450 ( .A(KEYINPUT111), .B(KEYINPUT47), .Z(n395) );
  XOR2_X1 U451 ( .A(KEYINPUT110), .B(n577), .Z(n565) );
  XOR2_X1 U452 ( .A(n458), .B(KEYINPUT64), .Z(n389) );
  XNOR2_X1 U453 ( .A(KEYINPUT41), .B(n389), .ZN(n553) );
  NOR2_X1 U454 ( .A1(n572), .A2(n553), .ZN(n390) );
  XNOR2_X1 U455 ( .A(n390), .B(KEYINPUT46), .ZN(n391) );
  NOR2_X1 U456 ( .A1(n565), .A2(n391), .ZN(n393) );
  BUF_X1 U457 ( .A(n392), .Z(n560) );
  NAND2_X1 U458 ( .A1(n393), .A2(n560), .ZN(n394) );
  XNOR2_X1 U459 ( .A(n395), .B(n394), .ZN(n396) );
  NOR2_X1 U460 ( .A1(n397), .A2(n396), .ZN(n398) );
  XNOR2_X1 U461 ( .A(KEYINPUT48), .B(n398), .ZN(n533) );
  XOR2_X1 U462 ( .A(KEYINPUT21), .B(G218GAT), .Z(n400) );
  XNOR2_X1 U463 ( .A(KEYINPUT82), .B(G204GAT), .ZN(n399) );
  XNOR2_X1 U464 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U465 ( .A(G197GAT), .B(n401), .Z(n428) );
  XOR2_X1 U466 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n403) );
  XNOR2_X1 U467 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n402) );
  XNOR2_X1 U468 ( .A(n403), .B(n402), .ZN(n437) );
  XNOR2_X1 U469 ( .A(n437), .B(n404), .ZN(n410) );
  XOR2_X1 U470 ( .A(n406), .B(n405), .Z(n408) );
  NAND2_X1 U471 ( .A1(G226GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U472 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U473 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U474 ( .A(n428), .B(n411), .ZN(n463) );
  NOR2_X1 U475 ( .A1(n521), .A2(n414), .ZN(n451) );
  XOR2_X1 U476 ( .A(G211GAT), .B(KEYINPUT83), .Z(n416) );
  XNOR2_X1 U477 ( .A(KEYINPUT22), .B(KEYINPUT84), .ZN(n415) );
  XNOR2_X1 U478 ( .A(n416), .B(n415), .ZN(n422) );
  XOR2_X1 U479 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n417) );
  XNOR2_X1 U480 ( .A(n418), .B(n417), .ZN(n420) );
  XNOR2_X1 U481 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U482 ( .A(n422), .B(n421), .Z(n424) );
  NAND2_X1 U483 ( .A1(G228GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U484 ( .A(n424), .B(n423), .ZN(n426) );
  XOR2_X1 U485 ( .A(n426), .B(n425), .Z(n430) );
  XNOR2_X1 U486 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U487 ( .A(KEYINPUT20), .B(KEYINPUT81), .Z(n432) );
  XNOR2_X1 U488 ( .A(G71GAT), .B(G183GAT), .ZN(n431) );
  XNOR2_X1 U489 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U490 ( .A(G176GAT), .B(G99GAT), .Z(n434) );
  XNOR2_X1 U491 ( .A(G43GAT), .B(G190GAT), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U493 ( .A(n436), .B(n435), .Z(n440) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U496 ( .A(n442), .B(n441), .Z(n444) );
  NAND2_X1 U497 ( .A1(G227GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n464) );
  INV_X1 U499 ( .A(n464), .ZN(n535) );
  NOR2_X1 U500 ( .A1(n466), .A2(n535), .ZN(n445) );
  XNOR2_X1 U501 ( .A(KEYINPUT26), .B(n445), .ZN(n549) );
  AND2_X1 U502 ( .A1(n451), .A2(n549), .ZN(n446) );
  NOR2_X1 U503 ( .A1(n458), .A2(n581), .ZN(n450) );
  XNOR2_X1 U504 ( .A(KEYINPUT125), .B(KEYINPUT61), .ZN(n448) );
  AND2_X1 U505 ( .A1(n466), .A2(n451), .ZN(n452) );
  XNOR2_X1 U506 ( .A(KEYINPUT55), .B(n452), .ZN(n453) );
  INV_X1 U507 ( .A(n553), .ZN(n539) );
  NAND2_X1 U508 ( .A1(n569), .A2(n539), .ZN(n457) );
  XOR2_X1 U509 ( .A(G176GAT), .B(KEYINPUT121), .Z(n455) );
  XOR2_X1 U510 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n454) );
  XNOR2_X1 U511 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U512 ( .A(n457), .B(n456), .ZN(G1349GAT) );
  XNOR2_X1 U513 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n482) );
  NAND2_X1 U514 ( .A1(n562), .A2(n458), .ZN(n459) );
  XNOR2_X1 U515 ( .A(n459), .B(KEYINPUT76), .ZN(n494) );
  XOR2_X2 U516 ( .A(n466), .B(KEYINPUT28), .Z(n537) );
  INV_X1 U517 ( .A(n463), .ZN(n524) );
  XNOR2_X1 U518 ( .A(KEYINPUT27), .B(n524), .ZN(n470) );
  NAND2_X1 U519 ( .A1(n521), .A2(n470), .ZN(n532) );
  NOR2_X1 U520 ( .A1(n537), .A2(n532), .ZN(n460) );
  NAND2_X1 U521 ( .A1(n461), .A2(n464), .ZN(n462) );
  XNOR2_X1 U522 ( .A(n462), .B(KEYINPUT91), .ZN(n475) );
  XOR2_X1 U523 ( .A(KEYINPUT25), .B(KEYINPUT93), .Z(n469) );
  NOR2_X1 U524 ( .A1(n464), .A2(n463), .ZN(n465) );
  XOR2_X1 U525 ( .A(KEYINPUT92), .B(n465), .Z(n467) );
  NAND2_X1 U526 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n469), .B(n468), .ZN(n472) );
  AND2_X1 U528 ( .A1(n549), .A2(n470), .ZN(n471) );
  NOR2_X1 U529 ( .A1(n472), .A2(n471), .ZN(n473) );
  NOR2_X1 U530 ( .A1(n521), .A2(n473), .ZN(n474) );
  XOR2_X1 U531 ( .A(KEYINPUT94), .B(n476), .Z(n490) );
  XOR2_X1 U532 ( .A(KEYINPUT16), .B(KEYINPUT80), .Z(n478) );
  INV_X1 U533 ( .A(n560), .ZN(n568) );
  OR2_X1 U534 ( .A1(n577), .A2(n568), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n478), .B(n477), .ZN(n479) );
  NAND2_X1 U536 ( .A1(n490), .A2(n479), .ZN(n508) );
  NOR2_X1 U537 ( .A1(n494), .A2(n508), .ZN(n480) );
  XOR2_X1 U538 ( .A(KEYINPUT95), .B(n480), .Z(n487) );
  NAND2_X1 U539 ( .A1(n521), .A2(n487), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n482), .B(n481), .ZN(G1324GAT) );
  NAND2_X1 U541 ( .A1(n487), .A2(n524), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n483), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT35), .B(KEYINPUT96), .Z(n485) );
  NAND2_X1 U544 ( .A1(n487), .A2(n535), .ZN(n484) );
  XNOR2_X1 U545 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U546 ( .A(G15GAT), .B(n486), .ZN(G1326GAT) );
  XOR2_X1 U547 ( .A(G22GAT), .B(KEYINPUT97), .Z(n489) );
  NAND2_X1 U548 ( .A1(n487), .A2(n537), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(G1327GAT) );
  AND2_X1 U550 ( .A1(n490), .A2(n577), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n491), .B(KEYINPUT99), .ZN(n492) );
  NOR2_X1 U552 ( .A1(n492), .A2(n582), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n493), .B(KEYINPUT37), .ZN(n520) );
  NOR2_X1 U554 ( .A1(n520), .A2(n494), .ZN(n495) );
  NAND2_X1 U555 ( .A1(n521), .A2(n504), .ZN(n497) );
  XOR2_X1 U556 ( .A(KEYINPUT98), .B(KEYINPUT39), .Z(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U558 ( .A(G29GAT), .B(n498), .ZN(G1328GAT) );
  XNOR2_X1 U559 ( .A(G36GAT), .B(KEYINPUT100), .ZN(n500) );
  NAND2_X1 U560 ( .A1(n524), .A2(n504), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(G1329GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT40), .B(KEYINPUT101), .Z(n502) );
  NAND2_X1 U563 ( .A1(n504), .A2(n535), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n506) );
  NAND2_X1 U567 ( .A1(n537), .A2(n504), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U569 ( .A(n507), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n511) );
  NAND2_X1 U571 ( .A1(n572), .A2(n539), .ZN(n519) );
  NOR2_X1 U572 ( .A1(n508), .A2(n519), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n509), .B(KEYINPUT104), .ZN(n514) );
  NAND2_X1 U574 ( .A1(n521), .A2(n514), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(G1332GAT) );
  NAND2_X1 U576 ( .A1(n514), .A2(n524), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U578 ( .A1(n514), .A2(n535), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n513), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n516) );
  NAND2_X1 U581 ( .A1(n537), .A2(n514), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(n518) );
  XOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT105), .Z(n517) );
  XNOR2_X1 U584 ( .A(n518), .B(n517), .ZN(G1335GAT) );
  XOR2_X1 U585 ( .A(G85GAT), .B(KEYINPUT107), .Z(n523) );
  NOR2_X1 U586 ( .A1(n520), .A2(n519), .ZN(n529) );
  NAND2_X1 U587 ( .A1(n529), .A2(n521), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n523), .B(n522), .ZN(G1336GAT) );
  NAND2_X1 U589 ( .A1(n529), .A2(n524), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n525), .B(KEYINPUT108), .ZN(n526) );
  XNOR2_X1 U591 ( .A(G92GAT), .B(n526), .ZN(G1337GAT) );
  XOR2_X1 U592 ( .A(G99GAT), .B(KEYINPUT109), .Z(n528) );
  NAND2_X1 U593 ( .A1(n529), .A2(n535), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n528), .B(n527), .ZN(G1338GAT) );
  NAND2_X1 U595 ( .A1(n529), .A2(n537), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n530), .B(KEYINPUT44), .ZN(n531) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  NOR2_X1 U598 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U599 ( .A(KEYINPUT115), .B(n534), .Z(n550) );
  NAND2_X1 U600 ( .A1(n550), .A2(n535), .ZN(n536) );
  NOR2_X1 U601 ( .A1(n537), .A2(n536), .ZN(n546) );
  NAND2_X1 U602 ( .A1(n546), .A2(n562), .ZN(n538) );
  XNOR2_X1 U603 ( .A(G113GAT), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n541) );
  NAND2_X1 U605 ( .A1(n546), .A2(n539), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U607 ( .A(G120GAT), .B(n542), .ZN(G1341GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n544) );
  NAND2_X1 U609 ( .A1(n546), .A2(n565), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n545), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U613 ( .A1(n546), .A2(n568), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  NAND2_X1 U615 ( .A1(n550), .A2(n549), .ZN(n559) );
  NOR2_X1 U616 ( .A1(n572), .A2(n559), .ZN(n551) );
  XOR2_X1 U617 ( .A(G141GAT), .B(n551), .Z(n552) );
  XNOR2_X1 U618 ( .A(KEYINPUT118), .B(n552), .ZN(G1344GAT) );
  NOR2_X1 U619 ( .A1(n559), .A2(n553), .ZN(n557) );
  XOR2_X1 U620 ( .A(KEYINPUT52), .B(KEYINPUT119), .Z(n555) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  NOR2_X1 U624 ( .A1(n577), .A2(n559), .ZN(n558) );
  XOR2_X1 U625 ( .A(G155GAT), .B(n558), .Z(G1346GAT) );
  NOR2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U627 ( .A(G162GAT), .B(n561), .Z(G1347GAT) );
  NAND2_X1 U628 ( .A1(n562), .A2(n569), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(KEYINPUT120), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G169GAT), .B(n564), .ZN(G1348GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n569), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(KEYINPUT122), .ZN(n567) );
  XNOR2_X1 U633 ( .A(G183GAT), .B(n567), .ZN(G1350GAT) );
  XNOR2_X1 U634 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n571) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1351GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n581), .ZN(n576) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(KEYINPUT60), .ZN(n574) );
  XNOR2_X1 U640 ( .A(KEYINPUT124), .B(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n581), .ZN(n578) );
  XOR2_X1 U643 ( .A(G211GAT), .B(n578), .Z(G1354GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n580) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n584) );
  NOR2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U648 ( .A(n584), .B(n583), .Z(G1355GAT) );
endmodule

