//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 0 1 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n805, new_n806,
    new_n807, new_n809, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n987, new_n988, new_n989, new_n991,
    new_n992, new_n993, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1022, new_n1023, new_n1024, new_n1025;
  INV_X1    g000(.A(G22gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G15gat), .ZN(new_n203));
  INV_X1    g002(.A(G15gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G22gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G1gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G8gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(KEYINPUT16), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n203), .A2(new_n205), .A3(new_n210), .ZN(new_n211));
  AND4_X1   g010(.A1(KEYINPUT94), .A2(new_n208), .A3(new_n209), .A4(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT94), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n213), .B1(new_n206), .B2(new_n207), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n209), .B1(new_n214), .B2(new_n211), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT21), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n218));
  INV_X1    g017(.A(G57gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G64gat), .ZN(new_n220));
  INV_X1    g019(.A(G64gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G57gat), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n218), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(G71gat), .A2(G78gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G71gat), .A2(G78gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(KEYINPUT96), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT96), .ZN(new_n228));
  INV_X1    g027(.A(new_n226), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n228), .B1(new_n229), .B2(new_n224), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n223), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n225), .A2(new_n226), .ZN(new_n232));
  XNOR2_X1  g031(.A(G57gat), .B(G64gat), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n232), .B(new_n228), .C1(new_n233), .C2(new_n218), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n216), .B1(new_n217), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G231gat), .ZN(new_n238));
  INV_X1    g037(.A(G233gat), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n235), .B(new_n217), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n238), .A2(new_n239), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n231), .A2(new_n234), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n241), .B1(new_n242), .B2(KEYINPUT21), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G127gat), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n244), .A2(G127gat), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n237), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n247), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n249), .A2(new_n236), .A3(new_n245), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(KEYINPUT97), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(G155gat), .ZN(new_n253));
  XOR2_X1   g052(.A(G183gat), .B(G211gat), .Z(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n248), .A2(new_n250), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n255), .B1(new_n248), .B2(new_n250), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(G43gat), .A2(G50gat), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NOR2_X1   g059(.A1(G43gat), .A2(G50gat), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT15), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G43gat), .ZN(new_n263));
  INV_X1    g062(.A(G50gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT15), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(new_n266), .A3(new_n259), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT14), .ZN(new_n268));
  INV_X1    g067(.A(G29gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n271));
  AOI21_X1  g070(.A(G36gat), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n269), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n262), .B(new_n267), .C1(new_n272), .C2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G36gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n271), .ZN(new_n277));
  NOR2_X1   g076(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n265), .A2(new_n259), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n279), .A2(new_n280), .A3(KEYINPUT15), .A4(new_n273), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT17), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n275), .A2(KEYINPUT17), .A3(new_n281), .ZN(new_n285));
  NAND2_X1  g084(.A1(G85gat), .A2(G92gat), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT7), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(KEYINPUT98), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G99gat), .A2(G106gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT8), .ZN(new_n290));
  INV_X1    g089(.A(G85gat), .ZN(new_n291));
  INV_X1    g090(.A(G92gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n288), .A2(new_n290), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n289), .ZN(new_n295));
  NOR2_X1   g094(.A1(G99gat), .A2(G106gat), .ZN(new_n296));
  OAI21_X1  g095(.A(KEYINPUT99), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OR2_X1    g096(.A1(G99gat), .A2(G106gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT99), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n299), .A3(new_n289), .ZN(new_n300));
  INV_X1    g099(.A(new_n286), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT98), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT7), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n287), .A2(KEYINPUT98), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n301), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n294), .A2(new_n297), .A3(new_n300), .A4(new_n305), .ZN(new_n306));
  AND3_X1   g105(.A1(new_n301), .A2(new_n303), .A3(new_n304), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n288), .A2(new_n290), .A3(new_n293), .ZN(new_n308));
  NOR3_X1   g107(.A1(new_n295), .A2(new_n296), .A3(KEYINPUT99), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n299), .B1(new_n298), .B2(new_n289), .ZN(new_n310));
  OAI22_X1  g109(.A1(new_n307), .A2(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n284), .A2(new_n285), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n282), .A2(new_n306), .A3(new_n311), .ZN(new_n314));
  NAND3_X1  g113(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n315));
  AND3_X1   g114(.A1(new_n314), .A2(KEYINPUT100), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT100), .B1(new_n314), .B2(new_n315), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n313), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  XOR2_X1   g117(.A(G190gat), .B(G218gat), .Z(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G134gat), .B(G162gat), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n321), .B(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n324), .A2(KEYINPUT101), .ZN(new_n325));
  INV_X1    g124(.A(new_n319), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n313), .B(new_n326), .C1(new_n316), .C2(new_n317), .ZN(new_n327));
  AND3_X1   g126(.A1(new_n320), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n323), .B(KEYINPUT101), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n330), .B1(new_n320), .B2(new_n327), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n312), .A2(new_n235), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT10), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n242), .A2(new_n306), .A3(new_n311), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n242), .A2(new_n306), .A3(new_n311), .A4(KEYINPUT10), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G230gat), .A2(G233gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n334), .A2(new_n336), .ZN(new_n342));
  INV_X1    g141(.A(new_n340), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G120gat), .B(G148gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(G176gat), .B(G204gat), .ZN(new_n346));
  XOR2_X1   g145(.A(new_n345), .B(new_n346), .Z(new_n347));
  NAND3_X1  g146(.A1(new_n341), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n347), .B1(new_n341), .B2(new_n344), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n258), .A2(new_n333), .A3(new_n351), .ZN(new_n352));
  XOR2_X1   g151(.A(KEYINPUT68), .B(G127gat), .Z(new_n353));
  INV_X1    g152(.A(G134gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(G120gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n356), .A2(G113gat), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(G113gat), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT1), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(G127gat), .A2(G134gat), .ZN(new_n361));
  NOR3_X1   g160(.A1(new_n355), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n356), .A2(KEYINPUT69), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT69), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(G120gat), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n364), .A2(new_n366), .A3(G113gat), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT70), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n367), .A2(new_n368), .A3(new_n358), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n368), .B1(new_n367), .B2(new_n358), .ZN(new_n370));
  AND2_X1   g169(.A1(G127gat), .A2(G134gat), .ZN(new_n371));
  AND2_X1   g170(.A1(KEYINPUT71), .A2(KEYINPUT1), .ZN(new_n372));
  NOR2_X1   g171(.A1(KEYINPUT71), .A2(KEYINPUT1), .ZN(new_n373));
  OAI22_X1  g172(.A1(new_n361), .A2(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NOR4_X1   g173(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT72), .A4(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT72), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n367), .A2(new_n358), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n374), .B1(new_n377), .B2(KEYINPUT70), .ZN(new_n378));
  XNOR2_X1  g177(.A(KEYINPUT69), .B(G120gat), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n357), .B1(new_n379), .B2(G113gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(new_n368), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n376), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n363), .B1(new_n375), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(G169gat), .A2(G176gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT23), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT23), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n386), .B1(G169gat), .B2(G176gat), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n385), .B1(new_n387), .B2(new_n384), .ZN(new_n388));
  NAND2_X1  g187(.A1(G183gat), .A2(G190gat), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n390));
  AND2_X1   g189(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n389), .A2(new_n390), .B1(new_n391), .B2(G190gat), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT25), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n388), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n390), .A2(new_n389), .ZN(new_n395));
  NAND3_X1  g194(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT66), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n395), .A2(KEYINPUT66), .A3(new_n396), .ZN(new_n400));
  NOR3_X1   g199(.A1(new_n386), .A2(G169gat), .A3(G176gat), .ZN(new_n401));
  INV_X1    g200(.A(new_n384), .ZN(new_n402));
  INV_X1    g201(.A(G169gat), .ZN(new_n403));
  INV_X1    g202(.A(G176gat), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT23), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n401), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n399), .A2(new_n400), .A3(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT65), .B(KEYINPUT25), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n394), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT26), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n384), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n411), .B(new_n412), .C1(new_n403), .C2(new_n404), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n389), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT27), .B(G183gat), .ZN(new_n415));
  INV_X1    g214(.A(G190gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT67), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n418), .A2(KEYINPUT28), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n415), .B(new_n416), .C1(new_n418), .C2(KEYINPUT28), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n414), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n409), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n383), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n420), .A2(new_n421), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n425), .A2(new_n389), .A3(new_n413), .ZN(new_n426));
  INV_X1    g225(.A(new_n408), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT66), .B1(new_n395), .B2(new_n396), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n428), .A2(new_n388), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n427), .B1(new_n429), .B2(new_n400), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n426), .B1(new_n430), .B2(new_n394), .ZN(new_n431));
  INV_X1    g230(.A(new_n374), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n432), .B1(new_n380), .B2(new_n368), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT72), .B1(new_n433), .B2(new_n369), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n378), .A2(new_n376), .A3(new_n381), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n431), .A2(new_n436), .A3(new_n363), .ZN(new_n437));
  NAND2_X1  g236(.A1(G227gat), .A2(G233gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(KEYINPUT64), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n424), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT33), .ZN(new_n441));
  XNOR2_X1  g240(.A(G15gat), .B(G43gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(G71gat), .B(G99gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n440), .B(KEYINPUT32), .C1(new_n441), .C2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n444), .B1(new_n440), .B2(new_n441), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n440), .A2(KEYINPUT73), .A3(KEYINPUT32), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT73), .B1(new_n440), .B2(KEYINPUT32), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n445), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT75), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n449), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n453), .A2(new_n447), .A3(new_n446), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n454), .A2(KEYINPUT75), .A3(new_n445), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n424), .A2(new_n437), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n457), .A2(KEYINPUT34), .A3(new_n439), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n456), .A2(KEYINPUT74), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT74), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n460), .B1(new_n424), .B2(new_n437), .ZN(new_n461));
  INV_X1    g260(.A(new_n438), .ZN(new_n462));
  OR3_X1    g261(.A1(new_n459), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n458), .B1(new_n463), .B2(KEYINPUT34), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n452), .A2(new_n455), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n458), .ZN(new_n466));
  NOR3_X1   g265(.A1(new_n459), .A2(new_n461), .A3(new_n462), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT34), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n469), .A2(KEYINPUT75), .A3(new_n445), .A4(new_n454), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n465), .A2(new_n470), .A3(KEYINPUT36), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT36), .B1(new_n465), .B2(new_n470), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AND2_X1   g272(.A1(G155gat), .A2(G162gat), .ZN(new_n474));
  NOR2_X1   g273(.A1(G155gat), .A2(G162gat), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(G141gat), .B(G148gat), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT2), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n478), .B1(G155gat), .B2(G162gat), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n476), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(G141gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(G148gat), .ZN(new_n482));
  INV_X1    g281(.A(G148gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(G141gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G155gat), .B(G162gat), .ZN(new_n486));
  INV_X1    g285(.A(G155gat), .ZN(new_n487));
  INV_X1    g286(.A(G162gat), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT2), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n485), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n480), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n363), .B(new_n492), .C1(new_n375), .C2(new_n382), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT3), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n480), .A2(new_n490), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT79), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT79), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n480), .A2(new_n490), .A3(new_n499), .A4(new_n496), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n498), .A2(new_n500), .B1(KEYINPUT3), .B2(new_n491), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n383), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(G225gat), .A2(G233gat), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n436), .A2(KEYINPUT4), .A3(new_n363), .A4(new_n492), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n495), .A2(new_n502), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT80), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n493), .A2(new_n494), .B1(new_n383), .B2(new_n501), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT80), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n507), .A2(new_n508), .A3(new_n503), .A4(new_n504), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n503), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n492), .B1(new_n436), .B2(new_n363), .ZN(new_n512));
  AOI211_X1 g311(.A(new_n362), .B(new_n491), .C1(new_n434), .C2(new_n435), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT6), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  XOR2_X1   g319(.A(G1gat), .B(G29gat), .Z(new_n521));
  XNOR2_X1  g320(.A(G57gat), .B(G85gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n521), .B(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n523), .B(new_n524), .Z(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n517), .A2(new_n518), .A3(new_n520), .A4(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(KEYINPUT6), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n518), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n515), .B1(new_n506), .B2(new_n509), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n528), .B(new_n529), .C1(new_n530), .C2(new_n519), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G211gat), .A2(G218gat), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT22), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(G197gat), .A2(G204gat), .ZN(new_n536));
  AND2_X1   g335(.A1(G197gat), .A2(G204gat), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  XOR2_X1   g337(.A(G211gat), .B(G218gat), .Z(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G211gat), .B(G218gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(G197gat), .B(G204gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(new_n542), .A3(new_n535), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(G226gat), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n546), .A2(new_n239), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n547), .A2(KEYINPUT29), .ZN(new_n548));
  INV_X1    g347(.A(new_n394), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n395), .A2(KEYINPUT66), .A3(new_n396), .ZN(new_n550));
  NOR3_X1   g349(.A1(new_n550), .A2(new_n428), .A3(new_n388), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n549), .B1(new_n551), .B2(new_n427), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n548), .B1(new_n552), .B2(new_n426), .ZN(new_n553));
  NOR3_X1   g352(.A1(new_n409), .A2(new_n422), .A3(new_n547), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n545), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT76), .ZN(new_n556));
  INV_X1    g355(.A(new_n548), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n557), .B1(new_n409), .B2(new_n422), .ZN(new_n558));
  INV_X1    g357(.A(new_n547), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n426), .B(new_n559), .C1(new_n430), .C2(new_n394), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n558), .A2(new_n544), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n555), .A2(new_n556), .A3(new_n561), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n558), .A2(new_n544), .A3(new_n560), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n544), .B1(new_n558), .B2(new_n560), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n563), .B1(new_n564), .B2(KEYINPUT76), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G8gat), .B(G36gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(G64gat), .B(G92gat), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n567), .B(new_n568), .Z(new_n569));
  NAND4_X1  g368(.A1(new_n566), .A2(KEYINPUT77), .A3(KEYINPUT30), .A4(new_n569), .ZN(new_n570));
  NOR3_X1   g369(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT76), .ZN(new_n571));
  NOR4_X1   g370(.A1(new_n553), .A2(new_n554), .A3(new_n556), .A4(new_n545), .ZN(new_n572));
  OAI211_X1 g371(.A(KEYINPUT30), .B(new_n569), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT77), .ZN(new_n574));
  INV_X1    g373(.A(new_n569), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n562), .A2(new_n565), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n573), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(KEYINPUT78), .B(KEYINPUT30), .Z(new_n578));
  AOI21_X1  g377(.A(new_n578), .B1(new_n566), .B2(new_n569), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n570), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n532), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT82), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT88), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n498), .A2(new_n500), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT29), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n544), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT3), .B1(new_n544), .B2(new_n585), .ZN(new_n587));
  OAI211_X1 g386(.A(G228gat), .B(G233gat), .C1(new_n587), .C2(new_n492), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT85), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G228gat), .A2(G233gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n538), .A2(new_n539), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n541), .B1(new_n535), .B2(new_n542), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n585), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(new_n496), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n590), .B1(new_n594), .B2(new_n491), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT85), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT29), .B1(new_n498), .B2(new_n500), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n595), .B(new_n596), .C1(new_n544), .C2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n589), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT87), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT29), .B1(new_n540), .B2(new_n543), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n496), .B1(new_n601), .B2(KEYINPUT84), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(KEYINPUT84), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n492), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n590), .B1(new_n605), .B2(new_n586), .ZN(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT86), .B(G22gat), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n599), .A2(new_n600), .A3(new_n606), .A4(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G78gat), .B(G106gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(KEYINPUT31), .B(G50gat), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n609), .B(new_n610), .Z(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n604), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n491), .B1(new_n613), .B2(new_n602), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n614), .B1(new_n544), .B2(new_n597), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n589), .A2(new_n598), .B1(new_n615), .B2(new_n590), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n608), .B(new_n612), .C1(new_n202), .C2(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n600), .B1(new_n616), .B2(new_n607), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n583), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n599), .A2(new_n606), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n611), .B1(new_n620), .B2(G22gat), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n599), .A2(new_n606), .A3(new_n607), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT87), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n621), .A2(new_n623), .A3(KEYINPUT88), .A4(new_n608), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n616), .B(new_n607), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n611), .B(KEYINPUT83), .Z(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT82), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n532), .A2(new_n580), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n582), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n473), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT93), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT91), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n555), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n564), .A2(KEYINPUT91), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n561), .A2(KEYINPUT90), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT90), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n558), .A2(new_n560), .A3(new_n639), .A4(new_n544), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n636), .A2(new_n637), .A3(new_n638), .A4(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT38), .B1(new_n641), .B2(KEYINPUT37), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT37), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n569), .B1(new_n566), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT92), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n566), .A2(new_n569), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT92), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n642), .A2(new_n644), .A3(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n646), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n634), .B1(new_n650), .B2(new_n532), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n649), .A2(new_n647), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n527), .A2(new_n531), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n652), .A2(new_n653), .A3(KEYINPUT93), .A4(new_n646), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n644), .B1(new_n643), .B2(new_n566), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(KEYINPUT38), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n651), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT89), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n526), .B1(new_n530), .B2(new_n519), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT39), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n512), .A2(new_n513), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n660), .B1(new_n661), .B2(new_n503), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n495), .A2(new_n504), .A3(new_n502), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(new_n511), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n526), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT40), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n663), .A2(new_n660), .A3(new_n511), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n666), .B1(new_n665), .B2(new_n667), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n659), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n658), .B1(new_n671), .B2(new_n580), .ZN(new_n672));
  INV_X1    g471(.A(new_n570), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n573), .A2(new_n574), .A3(new_n576), .ZN(new_n674));
  INV_X1    g473(.A(new_n579), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n662), .A2(new_n664), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n677), .A2(new_n525), .A3(new_n667), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(KEYINPUT40), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(new_n668), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n676), .A2(KEYINPUT89), .A3(new_n659), .A4(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n629), .B1(new_n672), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n657), .A2(new_n682), .ZN(new_n683));
  AOI22_X1  g482(.A1(new_n470), .A2(new_n465), .B1(new_n625), .B2(new_n628), .ZN(new_n684));
  AND3_X1   g483(.A1(new_n532), .A2(new_n580), .A3(new_n630), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n630), .B1(new_n532), .B2(new_n580), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(KEYINPUT35), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n581), .A2(KEYINPUT35), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n684), .ZN(new_n690));
  AOI22_X1  g489(.A1(new_n633), .A2(new_n683), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n216), .A2(new_n284), .A3(new_n285), .ZN(new_n692));
  NAND2_X1  g491(.A1(G229gat), .A2(G233gat), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n214), .A2(new_n211), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(G8gat), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n214), .A2(new_n209), .A3(new_n211), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n282), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n692), .A2(new_n693), .A3(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT18), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n692), .A2(new_n698), .A3(KEYINPUT18), .A4(new_n693), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n693), .B(KEYINPUT13), .Z(new_n703));
  AND2_X1   g502(.A1(new_n697), .A2(new_n282), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n697), .A2(new_n282), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n701), .A2(new_n702), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(G113gat), .B(G141gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(G197gat), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT11), .B(G169gat), .Z(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT12), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n707), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n701), .A2(new_n712), .A3(new_n702), .A4(new_n706), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT95), .B1(new_n691), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT95), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n473), .A2(new_n632), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n720), .B1(new_n657), .B2(new_n682), .ZN(new_n721));
  AOI22_X1  g520(.A1(new_n687), .A2(KEYINPUT35), .B1(new_n684), .B2(new_n689), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n719), .B(new_n716), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n352), .B1(new_n718), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n653), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g525(.A1(new_n718), .A2(new_n723), .ZN(new_n727));
  INV_X1    g526(.A(new_n352), .ZN(new_n728));
  XOR2_X1   g527(.A(KEYINPUT16), .B(G8gat), .Z(new_n729));
  NAND4_X1  g528(.A1(new_n727), .A2(new_n676), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT42), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT103), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  AOI211_X1 g531(.A(new_n580), .B(new_n352), .C1(new_n718), .C2(new_n723), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT103), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n733), .A2(new_n734), .A3(KEYINPUT42), .A4(new_n729), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n727), .A2(new_n728), .ZN(new_n737));
  OAI21_X1  g536(.A(G8gat), .B1(new_n737), .B2(new_n580), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT102), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n739), .B1(new_n730), .B2(new_n731), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n730), .A2(new_n739), .A3(new_n731), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n736), .B(new_n738), .C1(new_n740), .C2(new_n741), .ZN(G1325gat));
  OAI21_X1  g541(.A(G15gat), .B1(new_n737), .B2(new_n473), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n465), .A2(new_n470), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n724), .A2(new_n204), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(G1326gat));
  INV_X1    g545(.A(KEYINPUT104), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n625), .A2(new_n628), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n737), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n724), .A2(KEYINPUT104), .A3(new_n629), .ZN(new_n750));
  XNOR2_X1  g549(.A(KEYINPUT43), .B(G22gat), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n751), .B1(new_n749), .B2(new_n750), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n752), .A2(new_n753), .ZN(G1327gat));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n755), .B1(new_n691), .B2(new_n333), .ZN(new_n756));
  OAI211_X1 g555(.A(KEYINPUT44), .B(new_n332), .C1(new_n721), .C2(new_n722), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n258), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n351), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(new_n717), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(G29gat), .B1(new_n762), .B2(new_n532), .ZN(new_n763));
  AOI211_X1 g562(.A(new_n333), .B(new_n760), .C1(new_n718), .C2(new_n723), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n532), .A2(G29gat), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n765), .B1(new_n764), .B2(new_n766), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n763), .B1(new_n767), .B2(new_n768), .ZN(G1328gat));
  NAND3_X1  g568(.A1(new_n764), .A2(new_n276), .A3(new_n676), .ZN(new_n770));
  OR2_X1    g569(.A1(new_n770), .A2(KEYINPUT46), .ZN(new_n771));
  OAI21_X1  g570(.A(G36gat), .B1(new_n762), .B2(new_n580), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(KEYINPUT46), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(G1329gat));
  NAND3_X1  g573(.A1(new_n764), .A2(new_n263), .A3(new_n744), .ZN(new_n775));
  INV_X1    g574(.A(new_n473), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n756), .A2(new_n757), .A3(new_n776), .A4(new_n761), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G43gat), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT47), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n775), .A2(KEYINPUT47), .A3(new_n778), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(G1330gat));
  NAND2_X1  g582(.A1(new_n629), .A2(new_n264), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT105), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n764), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n756), .A2(new_n757), .A3(new_n629), .A4(new_n761), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G50gat), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT48), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n786), .A2(KEYINPUT48), .A3(new_n788), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(G1331gat));
  INV_X1    g592(.A(new_n351), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n258), .A2(new_n333), .A3(new_n717), .A4(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n691), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n653), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g597(.A1(new_n691), .A2(new_n580), .A3(new_n795), .ZN(new_n799));
  NOR2_X1   g598(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n800));
  AND2_X1   g599(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n802), .B1(new_n799), .B2(new_n800), .ZN(G1333gat));
  NAND3_X1  g602(.A1(new_n796), .A2(G71gat), .A3(new_n776), .ZN(new_n804));
  XOR2_X1   g603(.A(new_n744), .B(KEYINPUT106), .Z(new_n805));
  AND2_X1   g604(.A1(new_n796), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n806), .B2(G71gat), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g607(.A1(new_n796), .A2(new_n629), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g609(.A1(new_n258), .A2(new_n716), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n812), .A2(new_n351), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n758), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(G85gat), .B1(new_n814), .B2(new_n532), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n633), .A2(new_n683), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n688), .A2(new_n690), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n333), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT51), .B1(new_n818), .B2(new_n811), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n819), .A2(KEYINPUT107), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n811), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT51), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n818), .A2(KEYINPUT51), .A3(new_n811), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n820), .B1(new_n825), .B2(KEYINPUT107), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n653), .A2(new_n291), .A3(new_n794), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n815), .B1(new_n826), .B2(new_n827), .ZN(G1336gat));
  XOR2_X1   g627(.A(KEYINPUT109), .B(KEYINPUT52), .Z(new_n829));
  NAND4_X1  g628(.A1(new_n756), .A2(new_n757), .A3(new_n676), .A4(new_n813), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n829), .B1(new_n830), .B2(G92gat), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n676), .A2(new_n292), .A3(new_n794), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n831), .B1(new_n826), .B2(new_n832), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n830), .A2(KEYINPUT108), .A3(G92gat), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT108), .B1(new_n830), .B2(G92gat), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n832), .B1(new_n823), .B2(new_n824), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n833), .B1(new_n837), .B2(new_n838), .ZN(G1337gat));
  XOR2_X1   g638(.A(KEYINPUT110), .B(G99gat), .Z(new_n840));
  OAI21_X1  g639(.A(new_n840), .B1(new_n814), .B2(new_n473), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n351), .A2(new_n840), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n744), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(KEYINPUT111), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n841), .B1(new_n826), .B2(new_n844), .ZN(G1338gat));
  NAND4_X1  g644(.A1(new_n756), .A2(new_n757), .A3(new_n629), .A4(new_n813), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT53), .B1(new_n846), .B2(G106gat), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n748), .A2(G106gat), .A3(new_n351), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n847), .B1(new_n826), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT112), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n846), .A2(G106gat), .ZN(new_n852));
  NOR4_X1   g651(.A1(new_n691), .A2(new_n822), .A3(new_n333), .A4(new_n812), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n848), .B1(new_n819), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n851), .B1(new_n855), .B2(KEYINPUT53), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n857));
  AOI211_X1 g656(.A(KEYINPUT112), .B(new_n857), .C1(new_n852), .C2(new_n854), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n850), .B1(new_n856), .B2(new_n858), .ZN(G1339gat));
  NOR2_X1   g658(.A1(new_n352), .A2(new_n716), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT55), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n337), .A2(new_n338), .A3(new_n343), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n343), .B1(new_n337), .B2(new_n338), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n339), .A2(new_n864), .A3(new_n340), .ZN(new_n866));
  INV_X1    g665(.A(new_n347), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n861), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n337), .A2(new_n338), .A3(new_n343), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n341), .A2(KEYINPUT54), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n347), .B1(new_n863), .B2(new_n864), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(KEYINPUT55), .A3(new_n872), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n716), .A2(new_n869), .A3(new_n348), .A4(new_n873), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n704), .A2(new_n705), .A3(new_n703), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n693), .B1(new_n692), .B2(new_n698), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n711), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n715), .B(new_n877), .C1(new_n349), .C2(new_n350), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n333), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n869), .A2(new_n348), .A3(new_n873), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n314), .A2(new_n315), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT100), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n314), .A2(KEYINPUT100), .A3(new_n315), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n326), .B1(new_n886), .B2(new_n313), .ZN(new_n887));
  INV_X1    g686(.A(new_n327), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n329), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n320), .A2(new_n325), .A3(new_n327), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n889), .A2(new_n715), .A3(new_n890), .A4(new_n877), .ZN(new_n891));
  OAI21_X1  g690(.A(KEYINPUT113), .B1(new_n881), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n715), .A2(new_n877), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n328), .A2(new_n893), .A3(new_n331), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT113), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n873), .A2(new_n348), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n894), .A2(new_n895), .A3(new_n896), .A4(new_n869), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n880), .A2(new_n892), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n860), .B1(new_n898), .B2(new_n759), .ZN(new_n899));
  INV_X1    g698(.A(new_n684), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n653), .A2(new_n580), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n716), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(G113gat), .ZN(G1340gat));
  INV_X1    g703(.A(new_n902), .ZN(new_n905));
  OAI21_X1  g704(.A(G120gat), .B1(new_n905), .B2(new_n351), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n794), .A2(new_n379), .ZN(new_n907));
  XOR2_X1   g706(.A(new_n907), .B(KEYINPUT114), .Z(new_n908));
  OAI21_X1  g707(.A(new_n906), .B1(new_n905), .B2(new_n908), .ZN(G1341gat));
  NAND2_X1  g708(.A1(new_n902), .A2(new_n258), .ZN(new_n910));
  XOR2_X1   g709(.A(new_n910), .B(new_n353), .Z(G1342gat));
  NOR2_X1   g710(.A1(new_n905), .A2(new_n333), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n354), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n913), .A2(KEYINPUT56), .ZN(new_n914));
  XOR2_X1   g713(.A(new_n914), .B(KEYINPUT115), .Z(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(KEYINPUT56), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n915), .B(new_n916), .C1(new_n354), .C2(new_n912), .ZN(G1343gat));
  INV_X1    g716(.A(KEYINPUT58), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n776), .A2(new_n901), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n897), .A2(new_n892), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n332), .B1(new_n874), .B2(new_n878), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n759), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n860), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n748), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n919), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n716), .A2(new_n481), .ZN(new_n926));
  XOR2_X1   g725(.A(new_n926), .B(KEYINPUT118), .Z(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(KEYINPUT116), .B1(new_n924), .B2(KEYINPUT57), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT116), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT57), .ZN(new_n931));
  OAI211_X1 g730(.A(new_n930), .B(new_n931), .C1(new_n899), .C2(new_n748), .ZN(new_n932));
  AOI22_X1  g731(.A1(new_n929), .A2(new_n932), .B1(KEYINPUT57), .B2(new_n924), .ZN(new_n933));
  INV_X1    g732(.A(new_n919), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n933), .A2(new_n717), .A3(new_n934), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n918), .B(new_n928), .C1(new_n935), .C2(new_n481), .ZN(new_n936));
  INV_X1    g735(.A(new_n928), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n929), .A2(new_n932), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n939), .A2(KEYINPUT57), .A3(new_n629), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n941), .A2(KEYINPUT117), .A3(new_n919), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT117), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n943), .B1(new_n933), .B2(new_n934), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n942), .A2(new_n944), .A3(new_n716), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n937), .B1(new_n945), .B2(G141gat), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n936), .B1(new_n946), .B2(new_n918), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT119), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI211_X1 g748(.A(KEYINPUT119), .B(new_n936), .C1(new_n946), .C2(new_n918), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1344gat));
  NAND3_X1  g750(.A1(new_n925), .A2(new_n483), .A3(new_n794), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n483), .A2(KEYINPUT59), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n942), .A2(new_n944), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n953), .B1(new_n954), .B2(new_n351), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT120), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n894), .A2(new_n869), .A3(new_n896), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n258), .B1(new_n880), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n629), .B1(new_n959), .B2(new_n860), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(new_n931), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n961), .A2(new_n940), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n962), .A2(new_n934), .A3(new_n351), .ZN(new_n963));
  OAI21_X1  g762(.A(KEYINPUT59), .B1(new_n963), .B2(new_n483), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n957), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n955), .A2(new_n956), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n952), .B1(new_n965), .B2(new_n966), .ZN(G1345gat));
  OAI21_X1  g766(.A(G155gat), .B1(new_n954), .B2(new_n759), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n925), .A2(new_n487), .A3(new_n258), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(G1346gat));
  NOR3_X1   g769(.A1(new_n954), .A2(new_n488), .A3(new_n333), .ZN(new_n971));
  AOI21_X1  g770(.A(G162gat), .B1(new_n925), .B2(new_n332), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n971), .A2(new_n972), .ZN(G1347gat));
  NOR3_X1   g772(.A1(new_n629), .A2(new_n653), .A3(new_n580), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n805), .A2(new_n939), .A3(new_n974), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n975), .A2(new_n403), .A3(new_n717), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n939), .A2(new_n532), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n977), .B(KEYINPUT121), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n900), .A2(new_n580), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g779(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(new_n716), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n976), .B1(new_n982), .B2(new_n403), .ZN(G1348gat));
  OAI21_X1  g782(.A(G176gat), .B1(new_n975), .B2(new_n351), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n794), .A2(new_n404), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n984), .B1(new_n980), .B2(new_n985), .ZN(G1349gat));
  OAI21_X1  g785(.A(G183gat), .B1(new_n975), .B2(new_n759), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n258), .A2(new_n415), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n987), .B1(new_n980), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g788(.A(new_n989), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g789(.A1(new_n981), .A2(new_n416), .A3(new_n332), .ZN(new_n991));
  OAI21_X1  g790(.A(G190gat), .B1(new_n975), .B2(new_n333), .ZN(new_n992));
  XNOR2_X1  g791(.A(new_n992), .B(KEYINPUT61), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n991), .A2(new_n993), .ZN(G1351gat));
  NOR3_X1   g793(.A1(new_n776), .A2(new_n748), .A3(new_n580), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n995), .ZN(new_n996));
  INV_X1    g795(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g796(.A(G197gat), .B1(new_n997), .B2(new_n716), .ZN(new_n998));
  XNOR2_X1  g797(.A(new_n962), .B(KEYINPUT122), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n473), .A2(new_n532), .A3(new_n676), .ZN(new_n1000));
  INV_X1    g799(.A(G197gat), .ZN(new_n1001));
  NOR3_X1   g800(.A1(new_n1000), .A2(new_n1001), .A3(new_n717), .ZN(new_n1002));
  AOI21_X1  g801(.A(new_n998), .B1(new_n999), .B2(new_n1002), .ZN(G1352gat));
  NOR3_X1   g802(.A1(new_n996), .A2(G204gat), .A3(new_n351), .ZN(new_n1004));
  XNOR2_X1  g803(.A(new_n1004), .B(KEYINPUT62), .ZN(new_n1005));
  NOR2_X1   g804(.A1(new_n1000), .A2(new_n351), .ZN(new_n1006));
  AND2_X1   g805(.A1(new_n999), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g806(.A(KEYINPUT123), .ZN(new_n1008));
  AND2_X1   g807(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g808(.A(G204gat), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1010));
  OAI21_X1  g809(.A(new_n1005), .B1(new_n1009), .B2(new_n1010), .ZN(G1353gat));
  NOR3_X1   g810(.A1(new_n962), .A2(new_n759), .A3(new_n1000), .ZN(new_n1012));
  INV_X1    g811(.A(G211gat), .ZN(new_n1013));
  NOR2_X1   g812(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g813(.A1(KEYINPUT124), .A2(KEYINPUT63), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n997), .A2(new_n1013), .A3(new_n258), .ZN(new_n1017));
  XOR2_X1   g816(.A(KEYINPUT124), .B(KEYINPUT63), .Z(new_n1018));
  OAI21_X1  g817(.A(new_n1018), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1019));
  NAND3_X1  g818(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g819(.A(new_n1020), .B(KEYINPUT125), .ZN(G1354gat));
  AOI21_X1  g820(.A(G218gat), .B1(new_n997), .B2(new_n332), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n332), .A2(G218gat), .ZN(new_n1023));
  XOR2_X1   g822(.A(new_n1023), .B(KEYINPUT126), .Z(new_n1024));
  NOR2_X1   g823(.A1(new_n1000), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g824(.A(new_n1022), .B1(new_n999), .B2(new_n1025), .ZN(G1355gat));
endmodule


