//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004;
  INV_X1    g000(.A(KEYINPUT5), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT67), .ZN(new_n203));
  INV_X1    g002(.A(G113gat), .ZN(new_n204));
  AND2_X1   g003(.A1(new_n204), .A2(G120gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(G120gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G113gat), .B(G120gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT67), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n207), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(KEYINPUT66), .B(G127gat), .Z(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G134gat), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n211), .B(new_n213), .C1(G127gat), .C2(G134gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(G127gat), .B(G134gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n216));
  XOR2_X1   g015(.A(KEYINPUT68), .B(G120gat), .Z(new_n217));
  NOR2_X1   g016(.A1(new_n217), .A2(new_n204), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n215), .B(new_n216), .C1(new_n218), .C2(new_n205), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(G141gat), .B(G148gat), .Z(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT77), .ZN(new_n222));
  XNOR2_X1  g021(.A(G141gat), .B(G148gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT77), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT2), .ZN(new_n227));
  INV_X1    g026(.A(G155gat), .ZN(new_n228));
  INV_X1    g027(.A(G162gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  AOI22_X1  g029(.A1(new_n222), .A2(new_n225), .B1(new_n226), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT78), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n228), .A2(new_n229), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(new_n226), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n234), .B1(new_n221), .B2(new_n227), .ZN(new_n235));
  NOR3_X1   g034(.A1(new_n231), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n230), .A2(new_n226), .ZN(new_n237));
  INV_X1    g036(.A(new_n225), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n223), .A2(new_n224), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n235), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT78), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n220), .B1(new_n236), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n222), .A2(new_n225), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n235), .B1(new_n244), .B2(new_n237), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n214), .A2(new_n245), .A3(new_n219), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G225gat), .A2(G233gat), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n202), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n246), .A2(KEYINPUT80), .A3(KEYINPUT4), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT79), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT3), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n252), .B1(new_n245), .B2(new_n253), .ZN(new_n254));
  NOR4_X1   g053(.A1(new_n231), .A2(KEYINPUT79), .A3(KEYINPUT3), .A4(new_n235), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n220), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n245), .A2(KEYINPUT78), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n232), .B1(new_n231), .B2(new_n235), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n253), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n251), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n246), .A2(KEYINPUT4), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n214), .A2(new_n245), .A3(new_n262), .A4(new_n219), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT80), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n248), .B1(new_n261), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n250), .B1(new_n260), .B2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n268));
  XNOR2_X1  g067(.A(G1gat), .B(G29gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G57gat), .B(G85gat), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n270), .B(new_n271), .Z(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n259), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n240), .A2(new_n253), .A3(new_n241), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT79), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n245), .A2(new_n252), .A3(new_n253), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n276), .A2(new_n277), .B1(new_n214), .B2(new_n219), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n246), .A2(KEYINPUT4), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(new_n263), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n279), .A2(new_n202), .A3(new_n248), .A4(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n267), .A2(new_n273), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT82), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n267), .A2(new_n282), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(new_n272), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n267), .A2(new_n282), .A3(KEYINPUT82), .A4(new_n273), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n285), .A2(new_n287), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n273), .B1(new_n267), .B2(new_n282), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT6), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT26), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT65), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n295), .A2(new_n296), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT65), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n300), .B(new_n294), .C1(new_n295), .C2(new_n296), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n298), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT27), .B(G183gat), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT28), .B1(new_n304), .B2(G190gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(G183gat), .A2(G190gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT28), .ZN(new_n307));
  INV_X1    g106(.A(G190gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n303), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n302), .A2(new_n305), .A3(new_n306), .A4(new_n309), .ZN(new_n310));
  OR2_X1    g109(.A1(new_n295), .A2(KEYINPUT23), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n295), .A2(KEYINPUT23), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n311), .A2(new_n294), .A3(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT25), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT24), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n306), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317));
  OR2_X1    g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n319), .B(KEYINPUT64), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n313), .B(new_n314), .C1(new_n318), .C2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n311), .A2(new_n294), .A3(new_n312), .ZN(new_n322));
  NOR3_X1   g121(.A1(new_n316), .A2(new_n319), .A3(new_n317), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT25), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n310), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT29), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G226gat), .A2(G233gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n325), .A2(KEYINPUT71), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT71), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n310), .A2(new_n321), .A3(new_n331), .A4(new_n324), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n328), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT73), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT73), .ZN(new_n336));
  AOI211_X1 g135(.A(new_n336), .B(new_n328), .C1(new_n330), .C2(new_n332), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n329), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT70), .B(G197gat), .ZN(new_n339));
  INV_X1    g138(.A(G204gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G211gat), .ZN(new_n342));
  INV_X1    g141(.A(G218gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n341), .B1(KEYINPUT22), .B2(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(G211gat), .B(G218gat), .Z(new_n346));
  XNOR2_X1  g145(.A(new_n345), .B(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n338), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n326), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n328), .ZN(new_n350));
  INV_X1    g149(.A(new_n346), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n345), .B(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n325), .A2(new_n334), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(KEYINPUT72), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n350), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G64gat), .B(G92gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n356), .B(KEYINPUT76), .ZN(new_n357));
  XOR2_X1   g156(.A(G8gat), .B(G36gat), .Z(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n348), .A2(new_n355), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT30), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n361), .B1(new_n348), .B2(new_n355), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI211_X1 g164(.A(KEYINPUT30), .B(new_n361), .C1(new_n348), .C2(new_n355), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n293), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT83), .ZN(new_n368));
  INV_X1    g167(.A(new_n364), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(KEYINPUT30), .A3(new_n362), .ZN(new_n370));
  INV_X1    g169(.A(new_n366), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT83), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(new_n373), .A3(new_n293), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n368), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT85), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n276), .A2(new_n277), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT84), .B1(new_n377), .B2(new_n326), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT84), .ZN(new_n379));
  AOI211_X1 g178(.A(new_n379), .B(KEYINPUT29), .C1(new_n276), .C2(new_n277), .ZN(new_n380));
  NOR3_X1   g179(.A1(new_n378), .A2(new_n380), .A3(new_n347), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT3), .B1(new_n347), .B2(new_n326), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n257), .A2(new_n258), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  OAI211_X1 g183(.A(G228gat), .B(G233gat), .C1(new_n382), .C2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n376), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n378), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n377), .A2(KEYINPUT84), .A3(new_n326), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n352), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(G228gat), .A2(G233gat), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n253), .B1(new_n352), .B2(KEYINPUT29), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n390), .B1(new_n391), .B2(new_n383), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n389), .A2(KEYINPUT85), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n386), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n245), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n377), .A2(new_n326), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n352), .ZN(new_n398));
  AOI22_X1  g197(.A1(new_n396), .A2(new_n398), .B1(G228gat), .B2(G233gat), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n394), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(G106gat), .ZN(new_n402));
  INV_X1    g201(.A(G106gat), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n394), .A2(new_n403), .A3(new_n400), .ZN(new_n404));
  XNOR2_X1  g203(.A(G22gat), .B(G78gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT31), .B(G50gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n402), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n407), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n403), .B1(new_n394), .B2(new_n400), .ZN(new_n410));
  AOI211_X1 g209(.A(G106gat), .B(new_n399), .C1(new_n386), .C2(new_n393), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n361), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n348), .A2(new_n355), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT37), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n418), .B1(new_n417), .B2(new_n416), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT38), .ZN(new_n420));
  OR2_X1    g219(.A1(new_n291), .A2(KEYINPUT87), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n291), .A2(KEYINPUT87), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n285), .A2(new_n288), .A3(new_n289), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n423), .A2(new_n424), .B1(KEYINPUT6), .B2(new_n291), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT38), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n350), .A2(new_n354), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n347), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n428), .B(KEYINPUT37), .C1(new_n347), .C2(new_n338), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n418), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n420), .A2(new_n425), .A3(new_n369), .A4(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n365), .A2(new_n366), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n279), .A2(new_n281), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n249), .ZN(new_n434));
  OR2_X1    g233(.A1(new_n434), .A2(KEYINPUT39), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n434), .B(KEYINPUT39), .C1(new_n249), .C2(new_n247), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n436), .A3(new_n273), .ZN(new_n437));
  NOR2_X1   g236(.A1(KEYINPUT86), .A2(KEYINPUT40), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n435), .A2(new_n436), .A3(new_n273), .A4(new_n438), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n440), .A2(new_n441), .B1(new_n421), .B2(new_n422), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n432), .A2(new_n442), .B1(new_n408), .B2(new_n412), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n375), .A2(new_n414), .B1(new_n431), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n325), .B(new_n220), .ZN(new_n445));
  AND2_X1   g244(.A1(G227gat), .A2(G233gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT33), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(G15gat), .B(G43gat), .ZN(new_n450));
  INV_X1    g249(.A(G71gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n452), .B(G99gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n447), .A2(KEYINPUT32), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT34), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT34), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n447), .A2(KEYINPUT32), .A3(new_n457), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n445), .A2(new_n446), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n456), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n460), .B1(new_n456), .B2(new_n458), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n454), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n463), .ZN(new_n465));
  INV_X1    g264(.A(new_n454), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(new_n461), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n468), .B(KEYINPUT36), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n468), .B1(new_n408), .B2(new_n412), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n368), .A2(new_n471), .A3(new_n374), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT35), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT35), .ZN(new_n474));
  INV_X1    g273(.A(new_n425), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n471), .A2(new_n474), .A3(new_n475), .A4(new_n372), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n444), .A2(new_n470), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G183gat), .B(G211gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(KEYINPUT20), .ZN(new_n479));
  XNOR2_X1  g278(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(G231gat), .ZN(new_n483));
  INV_X1    g282(.A(G233gat), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT92), .B1(G71gat), .B2(G78gat), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NOR3_X1   g286(.A1(KEYINPUT92), .A2(G71gat), .A3(G78gat), .ZN(new_n488));
  NAND3_X1  g287(.A1(KEYINPUT91), .A2(G71gat), .A3(G78gat), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT91), .B1(G71gat), .B2(G78gat), .ZN(new_n491));
  OAI22_X1  g290(.A1(new_n487), .A2(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT93), .ZN(new_n493));
  INV_X1    g292(.A(G57gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(G64gat), .ZN(new_n495));
  INV_X1    g294(.A(G64gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(G57gat), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT9), .ZN(new_n498));
  NAND2_X1  g297(.A1(G71gat), .A2(G78gat), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n495), .A2(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT92), .ZN(new_n502));
  INV_X1    g301(.A(G78gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(new_n451), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n486), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT91), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n499), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n489), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT93), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n505), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n501), .A3(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(G71gat), .A2(G78gat), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n500), .A2(new_n499), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G15gat), .B(G22gat), .ZN(new_n518));
  INV_X1    g317(.A(G1gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT16), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(G1gat), .B2(new_n518), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n522), .A2(G8gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(G8gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT21), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n517), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n523), .A2(new_n524), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(KEYINPUT21), .B2(new_n516), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n517), .A2(new_n526), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  XOR2_X1   g330(.A(G127gat), .B(G155gat), .Z(new_n532));
  OR2_X1    g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n531), .A2(new_n532), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n485), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NOR3_X1   g336(.A1(new_n534), .A2(new_n485), .A3(new_n535), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n482), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n538), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n540), .A2(new_n536), .A3(new_n481), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(G162gat), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(G29gat), .A2(G36gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT14), .ZN(new_n548));
  NAND2_X1  g347(.A1(G29gat), .A2(G36gat), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n549), .A2(KEYINPUT14), .ZN(new_n550));
  OAI211_X1 g349(.A(KEYINPUT15), .B(new_n548), .C1(new_n550), .C2(new_n547), .ZN(new_n551));
  XNOR2_X1  g350(.A(G43gat), .B(G50gat), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT15), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n547), .B1(KEYINPUT14), .B2(new_n549), .ZN(new_n556));
  INV_X1    g355(.A(new_n548), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n558), .A2(new_n551), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n554), .B1(new_n559), .B2(new_n553), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT17), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n553), .B1(new_n558), .B2(new_n551), .ZN(new_n562));
  INV_X1    g361(.A(new_n554), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT17), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G85gat), .A2(G92gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT7), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT7), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n569), .A2(G85gat), .A3(G92gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(G99gat), .A2(G106gat), .ZN(new_n572));
  INV_X1    g371(.A(G85gat), .ZN(new_n573));
  INV_X1    g372(.A(G92gat), .ZN(new_n574));
  AOI22_X1  g373(.A1(KEYINPUT8), .A2(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G99gat), .B(G106gat), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n571), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT95), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n571), .A2(new_n576), .A3(new_n575), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n576), .B1(new_n571), .B2(new_n575), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n579), .B1(new_n582), .B2(new_n578), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n561), .A2(new_n566), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G232gat), .A2(G233gat), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT41), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n575), .ZN(new_n588));
  INV_X1    g387(.A(new_n576), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n590), .A2(new_n578), .A3(new_n577), .ZN(new_n591));
  INV_X1    g390(.A(new_n579), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n587), .B1(new_n564), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT96), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI211_X1 g395(.A(KEYINPUT96), .B(new_n587), .C1(new_n564), .C2(new_n593), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n584), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(G134gat), .ZN(new_n599));
  INV_X1    g398(.A(G134gat), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n600), .B(new_n584), .C1(new_n596), .C2(new_n597), .ZN(new_n601));
  XNOR2_X1  g400(.A(G190gat), .B(G218gat), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n599), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n603), .B1(new_n599), .B2(new_n601), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n546), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n599), .A2(new_n601), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(new_n602), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n609), .A2(new_n545), .A3(new_n604), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NOR3_X1   g410(.A1(new_n477), .A2(new_n543), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G113gat), .B(G141gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(G197gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT11), .ZN(new_n615));
  INV_X1    g414(.A(G169gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT12), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G229gat), .A2(G233gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT89), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n560), .A2(KEYINPUT17), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n528), .B1(new_n622), .B2(KEYINPUT88), .ZN(new_n623));
  AOI21_X1  g422(.A(KEYINPUT88), .B1(new_n523), .B2(new_n524), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n560), .B1(new_n624), .B2(KEYINPUT17), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n621), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT18), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n560), .B(new_n525), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n621), .B(KEYINPUT13), .Z(new_n629));
  OR2_X1    g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n626), .A2(KEYINPUT18), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n619), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(KEYINPUT90), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(new_n618), .ZN(new_n635));
  OAI211_X1 g434(.A(new_n627), .B(new_n630), .C1(new_n632), .C2(KEYINPUT90), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G230gat), .A2(G233gat), .ZN(new_n639));
  NOR3_X1   g438(.A1(new_n580), .A2(new_n581), .A3(KEYINPUT95), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n511), .B(new_n515), .C1(new_n640), .C2(new_n579), .ZN(new_n641));
  INV_X1    g440(.A(new_n582), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n505), .A2(new_n508), .A3(new_n509), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n509), .B1(new_n505), .B2(new_n508), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n643), .A2(new_n644), .A3(new_n500), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n642), .B1(new_n645), .B2(new_n514), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT10), .B1(new_n641), .B2(new_n646), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n593), .A2(new_n516), .A3(KEYINPUT10), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n639), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n639), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n641), .A2(new_n646), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G120gat), .B(G148gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT97), .ZN(new_n655));
  INV_X1    g454(.A(G176gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(new_n340), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n653), .A2(KEYINPUT98), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT98), .B1(new_n653), .B2(new_n659), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n653), .A2(KEYINPUT99), .A3(new_n659), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT99), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n663), .B1(new_n652), .B2(new_n658), .ZN(new_n664));
  OAI22_X1  g463(.A1(new_n660), .A2(new_n661), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n638), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n612), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n667), .A2(new_n293), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(new_n519), .ZN(G1324gat));
  NOR2_X1   g468(.A1(new_n667), .A2(new_n372), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT16), .ZN(new_n671));
  INV_X1    g470(.A(G8gat), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n673), .B1(new_n671), .B2(new_n672), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n670), .A2(new_n672), .ZN(new_n675));
  OAI21_X1  g474(.A(KEYINPUT42), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n676), .B1(KEYINPUT42), .B2(new_n674), .ZN(G1325gat));
  INV_X1    g476(.A(G15gat), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n667), .A2(new_n678), .A3(new_n470), .ZN(new_n679));
  INV_X1    g478(.A(new_n468), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n612), .A2(new_n666), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n679), .B1(new_n678), .B2(new_n681), .ZN(G1326gat));
  NOR2_X1   g481(.A1(new_n667), .A2(new_n413), .ZN(new_n683));
  XOR2_X1   g482(.A(KEYINPUT43), .B(G22gat), .Z(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1327gat));
  INV_X1    g484(.A(new_n611), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n477), .A2(new_n686), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n542), .A2(new_n638), .A3(new_n665), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(G29gat), .ZN(new_n690));
  INV_X1    g489(.A(new_n293), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT45), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n688), .B(KEYINPUT100), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n473), .A2(new_n476), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n367), .A2(KEYINPUT83), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n373), .B1(new_n372), .B2(new_n293), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n414), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n431), .A2(new_n443), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n700), .A2(new_n701), .A3(new_n470), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n696), .B1(new_n703), .B2(new_n611), .ZN(new_n704));
  AOI211_X1 g503(.A(KEYINPUT44), .B(new_n686), .C1(new_n697), .C2(new_n702), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n695), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(KEYINPUT101), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT44), .B1(new_n477), .B2(new_n686), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n703), .A2(new_n696), .A3(new_n611), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT101), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(new_n711), .A3(new_n695), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n293), .B1(new_n707), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n693), .B1(new_n690), .B2(new_n713), .ZN(G1328gat));
  INV_X1    g513(.A(G36gat), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n689), .A2(new_n715), .A3(new_n432), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n716), .B(KEYINPUT46), .Z(new_n717));
  AOI21_X1  g516(.A(new_n372), .B1(new_n707), .B2(new_n712), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n717), .B1(new_n715), .B2(new_n718), .ZN(G1329gat));
  OAI21_X1  g518(.A(G43gat), .B1(new_n706), .B2(new_n470), .ZN(new_n720));
  INV_X1    g519(.A(G43gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n689), .A2(new_n721), .A3(new_n680), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n720), .A2(KEYINPUT47), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n711), .B1(new_n710), .B2(new_n695), .ZN(new_n724));
  AOI211_X1 g523(.A(KEYINPUT101), .B(new_n694), .C1(new_n708), .C2(new_n709), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n469), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(G43gat), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n727), .A2(new_n722), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n723), .B1(new_n728), .B2(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g528(.A(new_n413), .B1(new_n707), .B2(new_n712), .ZN(new_n730));
  INV_X1    g529(.A(G50gat), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT102), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n414), .B1(new_n724), .B2(new_n725), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT102), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n733), .A2(new_n734), .A3(G50gat), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n689), .A2(new_n731), .A3(new_n414), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n732), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT48), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(G50gat), .B1(new_n706), .B2(new_n413), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n740), .A2(KEYINPUT48), .A3(new_n736), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n741), .ZN(G1331gat));
  NAND3_X1  g541(.A1(new_n542), .A2(new_n686), .A3(new_n638), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n477), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n665), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n745), .A2(new_n293), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(new_n494), .ZN(G1332gat));
  AOI211_X1 g546(.A(new_n372), .B(new_n745), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT103), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n748), .B(KEYINPUT103), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT49), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n752), .A2(new_n753), .A3(new_n496), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n751), .A2(new_n754), .ZN(G1333gat));
  NOR3_X1   g554(.A1(new_n745), .A2(new_n451), .A3(new_n470), .ZN(new_n756));
  XOR2_X1   g555(.A(new_n756), .B(KEYINPUT104), .Z(new_n757));
  OAI21_X1  g556(.A(new_n451), .B1(new_n745), .B2(new_n468), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT50), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT50), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n757), .A2(new_n761), .A3(new_n758), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(G1334gat));
  NOR2_X1   g562(.A1(new_n745), .A2(new_n413), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(new_n503), .ZN(G1335gat));
  NOR2_X1   g564(.A1(new_n542), .A2(new_n637), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n687), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(KEYINPUT51), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n687), .A2(new_n769), .A3(new_n766), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n665), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n773), .A2(new_n573), .A3(new_n691), .ZN(new_n774));
  INV_X1    g573(.A(new_n766), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n775), .A2(new_n772), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n704), .B2(new_n705), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT105), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT105), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n710), .A2(new_n779), .A3(new_n776), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n293), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n774), .B1(new_n573), .B2(new_n781), .ZN(G1336gat));
  AOI21_X1  g581(.A(new_n372), .B1(new_n778), .B2(new_n780), .ZN(new_n783));
  OAI21_X1  g582(.A(KEYINPUT106), .B1(new_n783), .B2(new_n574), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n779), .B1(new_n710), .B2(new_n776), .ZN(new_n785));
  INV_X1    g584(.A(new_n776), .ZN(new_n786));
  AOI211_X1 g585(.A(KEYINPUT105), .B(new_n786), .C1(new_n708), .C2(new_n709), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n432), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT106), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(new_n789), .A3(G92gat), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT107), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n767), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n771), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n372), .A2(G92gat), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n767), .A2(new_n791), .A3(new_n769), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n793), .A2(new_n665), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n784), .A2(new_n790), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT52), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT52), .B1(new_n773), .B2(new_n794), .ZN(new_n799));
  OAI21_X1  g598(.A(G92gat), .B1(new_n777), .B2(new_n372), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n801), .ZN(G1337gat));
  AOI21_X1  g601(.A(G99gat), .B1(new_n773), .B2(new_n680), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n470), .B1(new_n778), .B2(new_n780), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n803), .B1(G99gat), .B2(new_n804), .ZN(G1338gat));
  OAI21_X1  g604(.A(G106gat), .B1(new_n777), .B2(new_n413), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n413), .A2(new_n772), .A3(G106gat), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n768), .A2(new_n770), .A3(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n806), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n793), .A2(new_n795), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n414), .B1(new_n785), .B2(new_n787), .ZN(new_n812));
  AOI22_X1  g611(.A1(new_n811), .A2(new_n807), .B1(G106gat), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n810), .B1(new_n813), .B2(new_n809), .ZN(G1339gat));
  INV_X1    g613(.A(KEYINPUT10), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n583), .A2(new_n516), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n582), .B1(new_n511), .B2(new_n515), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n648), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n650), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n659), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n647), .A2(new_n639), .A3(new_n648), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT108), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n823), .B1(new_n824), .B2(new_n649), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n818), .A2(new_n824), .A3(new_n819), .A4(new_n650), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT54), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n825), .A2(KEYINPUT109), .A3(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT109), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n818), .A2(new_n650), .A3(new_n819), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n830), .B1(new_n820), .B2(KEYINPUT108), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n821), .B1(new_n823), .B2(new_n824), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n829), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n822), .B1(new_n828), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OR2_X1    g635(.A1(new_n660), .A2(new_n661), .ZN(new_n837));
  OAI211_X1 g636(.A(KEYINPUT55), .B(new_n822), .C1(new_n828), .C2(new_n833), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n836), .A2(new_n637), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n623), .A2(new_n621), .A3(new_n625), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT110), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n628), .A2(new_n629), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT110), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n623), .A2(new_n843), .A3(new_n621), .A4(new_n625), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n841), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n617), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n846), .A2(KEYINPUT111), .ZN(new_n847));
  INV_X1    g646(.A(new_n636), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n619), .B1(new_n632), .B2(KEYINPUT90), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n846), .A2(KEYINPUT111), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n847), .A2(new_n850), .A3(new_n665), .A4(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n611), .B1(new_n839), .B2(new_n852), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n836), .A2(new_n611), .A3(new_n837), .A4(new_n838), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n847), .A2(new_n850), .A3(new_n851), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n543), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n743), .A2(new_n665), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n857), .A2(KEYINPUT112), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(KEYINPUT112), .B1(new_n857), .B2(new_n858), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(new_n691), .A3(new_n471), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n862), .A2(new_n432), .ZN(new_n863));
  OAI21_X1  g662(.A(G113gat), .B1(new_n863), .B2(new_n638), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n862), .B(KEYINPUT113), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n372), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n637), .A2(new_n204), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n864), .B1(new_n866), .B2(new_n867), .ZN(G1340gat));
  NAND2_X1  g667(.A1(new_n372), .A2(new_n665), .ZN(new_n869));
  OAI21_X1  g668(.A(G120gat), .B1(new_n862), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n772), .A2(new_n217), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(KEYINPUT114), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n870), .B1(new_n866), .B2(new_n872), .ZN(G1341gat));
  INV_X1    g672(.A(new_n212), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n863), .A2(new_n874), .A3(new_n543), .ZN(new_n875));
  INV_X1    g674(.A(new_n866), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n542), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n875), .B1(new_n877), .B2(new_n874), .ZN(G1342gat));
  NAND4_X1  g677(.A1(new_n865), .A2(new_n600), .A3(new_n372), .A4(new_n611), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n879), .A2(KEYINPUT56), .ZN(new_n880));
  OAI21_X1  g679(.A(G134gat), .B1(new_n863), .B2(new_n686), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(KEYINPUT56), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(G1343gat));
  NOR2_X1   g682(.A1(new_n469), .A2(new_n293), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n372), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT57), .B1(new_n861), .B2(new_n414), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n857), .A2(new_n858), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(KEYINPUT57), .A3(new_n414), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT115), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n892), .B1(new_n857), .B2(new_n858), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(KEYINPUT115), .A3(new_n414), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n886), .B1(new_n887), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(G141gat), .B1(new_n896), .B2(new_n638), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n859), .A2(new_n860), .A3(new_n413), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n372), .A3(new_n884), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n899), .A2(G141gat), .A3(new_n638), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT58), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n897), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT116), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n893), .A2(KEYINPUT115), .A3(new_n414), .ZN(new_n905));
  AOI21_X1  g704(.A(KEYINPUT115), .B1(new_n893), .B2(new_n414), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT112), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n888), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n857), .A2(KEYINPUT112), .A3(new_n858), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n909), .A2(new_n414), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n892), .ZN(new_n912));
  AOI211_X1 g711(.A(new_n904), .B(new_n885), .C1(new_n907), .C2(new_n912), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n891), .B(new_n894), .C1(new_n898), .C2(KEYINPUT57), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT116), .B1(new_n914), .B2(new_n886), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n637), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n900), .B1(new_n916), .B2(G141gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n903), .B1(new_n917), .B2(new_n902), .ZN(G1344gat));
  XOR2_X1   g717(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n919));
  NAND2_X1  g718(.A1(new_n911), .A2(KEYINPUT57), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT119), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n858), .B(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n857), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n892), .B(new_n414), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n920), .A2(new_n924), .A3(new_n665), .A4(new_n886), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n919), .B1(new_n925), .B2(G148gat), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT120), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n926), .B(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n896), .A2(new_n904), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n914), .A2(KEYINPUT116), .A3(new_n886), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n772), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(G148gat), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n932), .A2(KEYINPUT59), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n931), .A2(KEYINPUT117), .A3(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT117), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n665), .B1(new_n913), .B2(new_n915), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(new_n933), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n928), .B1(new_n935), .B2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(new_n899), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n940), .A2(new_n932), .A3(new_n665), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(G1345gat));
  NOR3_X1   g741(.A1(new_n899), .A2(G155gat), .A3(new_n543), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n542), .B1(new_n913), .B2(new_n915), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n943), .B1(new_n944), .B2(G155gat), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT121), .ZN(G1346gat));
  NAND3_X1  g745(.A1(new_n940), .A2(new_n229), .A3(new_n611), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT122), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n686), .B1(new_n929), .B2(new_n930), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n949), .B2(new_n229), .ZN(G1347gat));
  NOR3_X1   g749(.A1(new_n859), .A2(new_n860), .A3(new_n691), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT123), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n471), .A2(new_n432), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n951), .A2(new_n952), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n956), .A2(new_n616), .A3(new_n637), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n951), .A2(new_n954), .ZN(new_n958));
  OAI21_X1  g757(.A(G169gat), .B1(new_n958), .B2(new_n638), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n959), .ZN(G1348gat));
  NOR3_X1   g759(.A1(new_n958), .A2(new_n656), .A3(new_n772), .ZN(new_n961));
  XOR2_X1   g760(.A(new_n961), .B(KEYINPUT124), .Z(new_n962));
  AOI21_X1  g761(.A(G176gat), .B1(new_n956), .B2(new_n665), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n962), .A2(new_n963), .ZN(G1349gat));
  NOR2_X1   g763(.A1(new_n543), .A2(new_n304), .ZN(new_n965));
  NAND4_X1  g764(.A1(new_n953), .A2(new_n954), .A3(new_n955), .A4(new_n965), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n951), .A2(new_n542), .A3(new_n954), .ZN(new_n967));
  AOI21_X1  g766(.A(KEYINPUT125), .B1(new_n967), .B2(G183gat), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(KEYINPUT126), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n966), .A2(new_n971), .A3(new_n968), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT60), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n973), .B(new_n974), .ZN(G1350gat));
  OAI21_X1  g774(.A(G190gat), .B1(new_n958), .B2(new_n686), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n976), .B(KEYINPUT61), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n956), .A2(new_n308), .A3(new_n611), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(G1351gat));
  AND2_X1   g778(.A1(new_n920), .A2(new_n924), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n469), .A2(new_n372), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(new_n293), .ZN(new_n982));
  INV_X1    g781(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g783(.A(G197gat), .B1(new_n984), .B2(new_n638), .ZN(new_n985));
  NAND4_X1  g784(.A1(new_n953), .A2(new_n414), .A3(new_n955), .A4(new_n981), .ZN(new_n986));
  OR2_X1    g785(.A1(new_n638), .A2(G197gat), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(G1352gat));
  NOR3_X1   g787(.A1(new_n986), .A2(G204gat), .A3(new_n772), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT62), .ZN(new_n990));
  OR2_X1    g789(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n989), .A2(new_n990), .ZN(new_n992));
  AND2_X1   g791(.A1(new_n980), .A2(new_n665), .ZN(new_n993));
  AND2_X1   g792(.A1(new_n993), .A2(new_n983), .ZN(new_n994));
  OAI211_X1 g793(.A(new_n991), .B(new_n992), .C1(new_n340), .C2(new_n994), .ZN(G1353gat));
  INV_X1    g794(.A(new_n984), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n996), .A2(new_n542), .ZN(new_n997));
  AND3_X1   g796(.A1(new_n997), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n998));
  AOI21_X1  g797(.A(KEYINPUT63), .B1(new_n997), .B2(G211gat), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n542), .A2(new_n342), .ZN(new_n1000));
  OAI22_X1  g799(.A1(new_n998), .A2(new_n999), .B1(new_n986), .B2(new_n1000), .ZN(G1354gat));
  OAI21_X1  g800(.A(new_n343), .B1(new_n986), .B2(new_n686), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n611), .A2(G218gat), .ZN(new_n1003));
  OAI21_X1  g802(.A(new_n1002), .B1(new_n984), .B2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g803(.A(new_n1004), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


