//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 0 0 0 0 0 0 0 0 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 0 1 0 0 1 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n206), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  OR3_X1    g0017(.A1(new_n206), .A2(KEYINPUT64), .A3(G13), .ZN(new_n218));
  OAI21_X1  g0018(.A(KEYINPUT64), .B1(new_n206), .B2(G13), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT0), .Z(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(new_n201), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G50), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  AOI211_X1 g0028(.A(new_n217), .B(new_n222), .C1(new_n225), .C2(new_n228), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT65), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT66), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  INV_X1    g0046(.A(G274), .ZN(new_n247));
  AND2_X1   g0047(.A1(G1), .A2(G13), .ZN(new_n248));
  NAND2_X1  g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  AOI21_X1  g0049(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G41), .A2(G45), .ZN(new_n251));
  OAI21_X1  g0051(.A(KEYINPUT67), .B1(new_n251), .B2(G1), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT67), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n253), .B(new_n254), .C1(G41), .C2(G45), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n250), .A2(new_n252), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n248), .A2(new_n249), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n254), .B1(G41), .B2(G45), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(G232), .A3(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G33), .ZN(new_n264));
  INV_X1    g0064(.A(G1698), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n262), .A2(new_n264), .A3(G223), .A4(new_n265), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n262), .A2(new_n264), .A3(G226), .A4(G1698), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G87), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G179), .ZN(new_n272));
  AND3_X1   g0072(.A1(new_n260), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(G169), .B1(new_n260), .B2(new_n271), .ZN(new_n274));
  OAI21_X1  g0074(.A(KEYINPUT78), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G169), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n269), .A2(new_n270), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n256), .A2(new_n259), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT78), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n260), .A2(new_n271), .A3(new_n272), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n275), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT77), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT8), .B(G58), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT68), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n287), .B(new_n223), .C1(G1), .C2(new_n224), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT8), .ZN(new_n289));
  OR3_X1    g0089(.A1(new_n289), .A2(KEYINPUT68), .A3(G58), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n286), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n286), .A2(new_n290), .ZN(new_n292));
  INV_X1    g0092(.A(G13), .ZN(new_n293));
  NOR3_X1   g0093(.A1(new_n293), .A2(new_n224), .A3(G1), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n284), .B(new_n291), .C1(new_n292), .C2(new_n294), .ZN(new_n295));
  AND3_X1   g0095(.A1(new_n286), .A2(new_n288), .A3(new_n290), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n294), .B1(new_n286), .B2(new_n290), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT77), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT16), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT76), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n262), .A2(new_n264), .ZN(new_n302));
  AOI21_X1  g0102(.A(KEYINPUT7), .B1(new_n302), .B2(new_n224), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT7), .ZN(new_n304));
  AOI211_X1 g0104(.A(new_n304), .B(G20), .C1(new_n262), .C2(new_n264), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n301), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  XNOR2_X1  g0106(.A(KEYINPUT3), .B(G33), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n304), .B1(new_n307), .B2(G20), .ZN(new_n308));
  OAI21_X1  g0108(.A(KEYINPUT76), .B1(new_n308), .B2(KEYINPUT7), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n208), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G58), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n311), .A2(new_n208), .ZN(new_n312));
  OAI21_X1  g0112(.A(G20), .B1(new_n312), .B2(new_n201), .ZN(new_n313));
  NOR2_X1   g0113(.A1(G20), .A2(G33), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G159), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n300), .B1(new_n310), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(G68), .B1(new_n303), .B2(new_n305), .ZN(new_n318));
  INV_X1    g0118(.A(new_n316), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n318), .A2(KEYINPUT16), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n287), .A2(new_n223), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n299), .B1(new_n317), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(KEYINPUT18), .B1(new_n283), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n275), .A2(new_n282), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n295), .A2(new_n298), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n302), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n327));
  AOI21_X1  g0127(.A(KEYINPUT76), .B1(new_n308), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n302), .A2(new_n224), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n301), .B1(new_n329), .B2(new_n304), .ZN(new_n330));
  OAI21_X1  g0130(.A(G68), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT16), .B1(new_n331), .B2(new_n319), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n320), .A2(new_n321), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n326), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT18), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n325), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G200), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(new_n277), .B2(new_n278), .ZN(new_n338));
  INV_X1    g0138(.A(G190), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n260), .A2(new_n271), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n341), .B(new_n326), .C1(new_n332), .C2(new_n333), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT17), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n323), .A2(KEYINPUT17), .A3(new_n341), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n324), .A2(new_n336), .A3(new_n344), .A4(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT71), .ZN(new_n348));
  OR2_X1    g0148(.A1(new_n348), .A2(KEYINPUT10), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(KEYINPUT10), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n307), .A2(G222), .A3(new_n265), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n307), .A2(G223), .A3(G1698), .ZN(new_n352));
  INV_X1    g0152(.A(G77), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n351), .B(new_n352), .C1(new_n353), .C2(new_n307), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n270), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n257), .A2(G226), .A3(new_n258), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n256), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT70), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(new_n360), .A3(G200), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n357), .B1(new_n354), .B2(new_n270), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT70), .B1(new_n362), .B2(new_n337), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(G50), .B1(new_n224), .B2(G1), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n365), .B(KEYINPUT69), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n294), .A2(new_n321), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n366), .A2(new_n367), .B1(new_n202), .B2(new_n294), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n261), .A2(G20), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n286), .A2(new_n369), .A3(new_n290), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n314), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n321), .ZN(new_n373));
  OAI211_X1 g0173(.A(KEYINPUT9), .B(new_n368), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n362), .A2(G190), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT9), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n373), .B1(new_n370), .B2(new_n371), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT69), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n365), .B(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n293), .A2(G1), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(G20), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n373), .A2(new_n381), .ZN(new_n382));
  OAI22_X1  g0182(.A1(new_n379), .A2(new_n382), .B1(G50), .B2(new_n381), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n376), .B1(new_n377), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n374), .A2(new_n375), .A3(new_n384), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n349), .B(new_n350), .C1(new_n364), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n294), .A2(new_n353), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n353), .B2(new_n288), .ZN(new_n388));
  XOR2_X1   g0188(.A(KEYINPUT15), .B(G87), .Z(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n369), .ZN(new_n390));
  INV_X1    g0190(.A(new_n314), .ZN(new_n391));
  OAI221_X1 g0191(.A(new_n390), .B1(new_n224), .B2(new_n353), .C1(new_n391), .C2(new_n285), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n388), .B1(new_n392), .B2(new_n321), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n307), .A2(G232), .A3(new_n265), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n307), .A2(G238), .A3(G1698), .ZN(new_n395));
  INV_X1    g0195(.A(G107), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n394), .B(new_n395), .C1(new_n396), .C2(new_n307), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n270), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n257), .A2(new_n258), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G244), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(new_n256), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n393), .B1(new_n401), .B2(new_n276), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(G179), .B2(new_n401), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n377), .A2(new_n383), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n404), .B1(new_n276), .B2(new_n359), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(G179), .B2(new_n359), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n401), .A2(G200), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n407), .B(new_n393), .C1(new_n339), .C2(new_n401), .ZN(new_n408));
  AND3_X1   g0208(.A1(new_n403), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n361), .A2(new_n363), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n374), .A2(new_n375), .A3(new_n384), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n410), .A2(new_n348), .A3(KEYINPUT10), .A4(new_n411), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n347), .A2(new_n386), .A3(new_n409), .A4(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n307), .A2(G232), .A3(G1698), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n307), .A2(G226), .A3(new_n265), .ZN(new_n415));
  NAND2_X1  g0215(.A1(G33), .A2(G97), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n270), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n250), .A2(new_n252), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n419), .A2(new_n255), .B1(G238), .B2(new_n399), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT13), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT72), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT13), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n418), .A2(new_n420), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n422), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n418), .A2(new_n420), .A3(KEYINPUT72), .A4(new_n424), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n426), .A2(G169), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT14), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT73), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n422), .A2(new_n430), .A3(new_n425), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n421), .A2(KEYINPUT73), .A3(KEYINPUT13), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(G179), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT14), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n426), .A2(new_n435), .A3(G169), .A4(new_n427), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n429), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n288), .A2(new_n208), .ZN(new_n438));
  XNOR2_X1  g0238(.A(new_n438), .B(KEYINPUT74), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n294), .A2(new_n208), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n440), .B(KEYINPUT12), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT75), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n369), .A2(G77), .ZN(new_n445));
  OAI221_X1 g0245(.A(new_n445), .B1(new_n224), .B2(G68), .C1(new_n202), .C2(new_n391), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n321), .ZN(new_n447));
  XNOR2_X1  g0247(.A(new_n447), .B(KEYINPUT11), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n439), .A2(KEYINPUT75), .A3(new_n441), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n444), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n437), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n450), .B1(new_n433), .B2(G190), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n426), .A2(G200), .A3(new_n427), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n413), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n262), .A2(new_n264), .A3(G244), .A4(new_n265), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT4), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n307), .A2(KEYINPUT4), .A3(G244), .A4(new_n265), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n307), .A2(G250), .A3(G1698), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n460), .A2(new_n461), .A3(new_n462), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n270), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT5), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT81), .B1(new_n467), .B2(G41), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT81), .ZN(new_n469));
  INV_X1    g0269(.A(G41), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n469), .A2(new_n470), .A3(KEYINPUT5), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n467), .A2(G41), .ZN(new_n472));
  INV_X1    g0272(.A(G45), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(G1), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n468), .A2(new_n471), .A3(new_n472), .A4(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n475), .A2(G257), .A3(new_n257), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT82), .ZN(new_n477));
  INV_X1    g0277(.A(new_n250), .ZN(new_n478));
  OR2_X1    g0278(.A1(new_n478), .A2(new_n475), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT82), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n475), .A2(new_n480), .A3(G257), .A4(new_n257), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n276), .B1(new_n466), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(G107), .B1(new_n328), .B2(new_n330), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT6), .ZN(new_n485));
  INV_X1    g0285(.A(G97), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(new_n396), .ZN(new_n487));
  NOR2_X1   g0287(.A1(G97), .A2(G107), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n396), .A2(KEYINPUT6), .A3(G97), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n491), .A2(G20), .B1(G77), .B2(new_n314), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n373), .B1(new_n484), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n367), .B1(G1), .B2(new_n261), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT79), .B1(new_n381), .B2(G97), .ZN(new_n496));
  OR3_X1    g0296(.A1(new_n381), .A2(KEYINPUT79), .A3(G97), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n495), .A2(G97), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n483), .B1(new_n493), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n465), .A2(KEYINPUT80), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT80), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n464), .A2(new_n502), .A3(new_n270), .ZN(new_n503));
  AOI211_X1 g0303(.A(G179), .B(new_n482), .C1(new_n501), .C2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT83), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n500), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n396), .B1(new_n306), .B2(new_n309), .ZN(new_n507));
  INV_X1    g0307(.A(new_n492), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n321), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n465), .A2(new_n477), .A3(new_n479), .A4(new_n481), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n509), .A2(new_n498), .B1(new_n276), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n501), .A2(new_n503), .ZN(new_n512));
  INV_X1    g0312(.A(new_n482), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n512), .A2(new_n272), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT83), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n506), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT88), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n493), .A2(new_n499), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n466), .A2(new_n482), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G190), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n482), .B1(new_n501), .B2(new_n503), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n518), .B(new_n520), .C1(new_n337), .C2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n307), .A2(G238), .A3(new_n265), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n307), .A2(G244), .A3(G1698), .ZN(new_n524));
  OR2_X1    g0324(.A1(KEYINPUT85), .A2(G116), .ZN(new_n525));
  NAND2_X1  g0325(.A1(KEYINPUT85), .A2(G116), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G33), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n523), .A2(new_n524), .A3(new_n528), .ZN(new_n529));
  AND2_X1   g0329(.A1(new_n529), .A2(new_n270), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n250), .A2(new_n474), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n474), .A2(new_n211), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n532), .A2(KEYINPUT84), .A3(new_n257), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(KEYINPUT84), .B1(new_n532), .B2(new_n257), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n531), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(G200), .B1(new_n530), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n495), .A2(KEYINPUT87), .A3(G87), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT87), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n494), .B2(new_n210), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n307), .A2(new_n224), .A3(G68), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT86), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT86), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n307), .A2(new_n544), .A3(new_n224), .A4(G68), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT19), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n369), .A2(new_n546), .A3(G97), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n488), .A2(new_n210), .B1(new_n416), .B2(new_n224), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n547), .B1(new_n548), .B2(new_n546), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n543), .A2(new_n545), .A3(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n389), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n550), .A2(new_n321), .B1(new_n294), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n532), .A2(new_n257), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT84), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n555), .A2(new_n533), .B1(new_n474), .B2(new_n250), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n529), .A2(new_n270), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(G190), .A3(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n537), .A2(new_n541), .A3(new_n552), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n550), .A2(new_n321), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n495), .A2(new_n389), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n551), .A2(new_n294), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n276), .B1(new_n530), .B2(new_n536), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n556), .A2(new_n272), .A3(new_n557), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n559), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n516), .A2(new_n517), .A3(new_n522), .A4(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n505), .B1(new_n500), .B2(new_n504), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n509), .A2(new_n498), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n514), .A2(new_n570), .A3(KEYINPUT83), .A4(new_n483), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n569), .A2(new_n571), .A3(new_n522), .A4(new_n567), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(KEYINPUT88), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n262), .A2(new_n264), .A3(new_n224), .A4(G87), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT22), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n576), .A2(KEYINPUT90), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n307), .A2(new_n224), .A3(G87), .A4(new_n577), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n527), .A2(new_n224), .A3(G33), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT23), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n224), .B2(G107), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n396), .A2(KEYINPUT23), .A3(G20), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n579), .A2(new_n580), .A3(new_n581), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT24), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n261), .B1(new_n525), .B2(new_n526), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n588), .A2(new_n224), .B1(new_n583), .B2(new_n584), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT24), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n589), .A2(new_n590), .A3(new_n580), .A4(new_n579), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n321), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT25), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n381), .B2(G107), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n294), .A2(KEYINPUT25), .A3(new_n396), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n494), .B2(new_n396), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n262), .A2(new_n264), .A3(G257), .A4(G1698), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n262), .A2(new_n264), .A3(G250), .A4(new_n265), .ZN(new_n602));
  NAND2_X1  g0402(.A1(G33), .A2(G294), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n270), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n475), .A2(G264), .A3(new_n257), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n479), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n276), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n605), .A2(new_n479), .A3(new_n272), .A4(new_n606), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n600), .A2(new_n610), .A3(KEYINPUT91), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT91), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n598), .B1(new_n592), .B2(new_n321), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n608), .A2(new_n609), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OR2_X1    g0415(.A1(new_n607), .A2(new_n339), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n607), .A2(G200), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n613), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n611), .A2(new_n615), .A3(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT92), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n611), .A2(new_n615), .A3(KEYINPUT92), .A4(new_n618), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(G116), .ZN(new_n624));
  OAI22_X1  g0424(.A1(new_n494), .A2(new_n624), .B1(new_n381), .B2(new_n527), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n462), .B(new_n224), .C1(G33), .C2(new_n486), .ZN(new_n627));
  XNOR2_X1  g0427(.A(new_n627), .B(KEYINPUT89), .ZN(new_n628));
  INV_X1    g0428(.A(new_n527), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n373), .B1(new_n629), .B2(G20), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n628), .A2(new_n630), .A3(KEYINPUT20), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(KEYINPUT20), .B1(new_n628), .B2(new_n630), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n626), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n307), .A2(G257), .A3(new_n265), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n307), .A2(G264), .A3(G1698), .ZN(new_n636));
  INV_X1    g0436(.A(G303), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n635), .B(new_n636), .C1(new_n637), .C2(new_n307), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n270), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n475), .A2(G270), .A3(new_n257), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(new_n479), .A3(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n634), .A2(KEYINPUT21), .A3(G169), .A4(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n272), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n634), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT21), .ZN(new_n646));
  INV_X1    g0446(.A(new_n633), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n625), .B1(new_n647), .B2(new_n631), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n641), .A2(G169), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n641), .A2(G200), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n648), .B(new_n651), .C1(new_n339), .C2(new_n641), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n645), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  NOR4_X1   g0453(.A1(new_n457), .A2(new_n574), .A3(new_n623), .A4(new_n653), .ZN(G372));
  NOR2_X1   g0454(.A1(new_n500), .A2(new_n504), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT26), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(new_n567), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n566), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n567), .B1(new_n506), .B2(new_n515), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n658), .B1(KEYINPUT26), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n618), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n600), .A2(new_n610), .ZN(new_n662));
  AND4_X1   g0462(.A1(new_n662), .A2(new_n650), .A3(new_n644), .A4(new_n642), .ZN(new_n663));
  OR3_X1    g0463(.A1(new_n572), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n456), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n324), .A2(new_n336), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n451), .A2(new_n403), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n345), .A2(new_n344), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n669), .A2(new_n454), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n667), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n412), .A2(new_n386), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT93), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n412), .A2(new_n386), .A3(KEYINPUT93), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n406), .B1(new_n671), .B2(new_n677), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n666), .A2(new_n678), .ZN(G369));
  NAND2_X1  g0479(.A1(new_n380), .A2(new_n224), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(new_n682), .A3(G213), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n648), .A2(new_n686), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n653), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n645), .A2(new_n650), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n687), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G330), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n662), .A2(new_n686), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n621), .A2(new_n622), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n600), .A2(new_n685), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n689), .A2(new_n686), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n623), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n662), .A2(new_n685), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n698), .A2(new_n702), .ZN(G399));
  INV_X1    g0503(.A(new_n220), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G41), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n488), .A2(new_n210), .A3(new_n624), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n705), .A2(new_n254), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n228), .B2(new_n705), .ZN(new_n708));
  XNOR2_X1  g0508(.A(KEYINPUT94), .B(KEYINPUT28), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n708), .B(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT29), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n665), .A2(new_n711), .A3(new_n686), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n659), .A2(KEYINPUT96), .A3(new_n656), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT96), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n559), .A2(new_n566), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n715), .B1(new_n569), .B2(new_n571), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n714), .B1(new_n716), .B2(KEYINPUT26), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n655), .A2(new_n567), .A3(KEYINPUT26), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n713), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n566), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n572), .A2(new_n661), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n611), .A2(new_n615), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(new_n650), .A3(new_n645), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n720), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n685), .B1(new_n719), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n712), .B1(new_n725), .B2(new_n711), .ZN(new_n726));
  INV_X1    g0526(.A(G330), .ZN(new_n727));
  AND4_X1   g0527(.A1(new_n557), .A2(new_n556), .A3(new_n606), .A4(new_n605), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n643), .A2(new_n728), .A3(new_n519), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n643), .A2(new_n728), .A3(new_n519), .A4(KEYINPUT30), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n556), .A2(new_n557), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n641), .A2(new_n733), .A3(new_n272), .A4(new_n607), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n731), .B(new_n732), .C1(new_n521), .C2(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n685), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(KEYINPUT95), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT95), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n735), .A2(new_n738), .A3(KEYINPUT31), .A4(new_n685), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n735), .A2(new_n685), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT31), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n737), .A2(new_n739), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n653), .B1(new_n621), .B2(new_n622), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n744), .A2(new_n568), .A3(new_n573), .A4(new_n686), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n727), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n726), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n710), .B1(new_n747), .B2(G1), .ZN(G364));
  XOR2_X1   g0548(.A(new_n692), .B(KEYINPUT97), .Z(new_n749));
  NOR2_X1   g0549(.A1(new_n293), .A2(G20), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n254), .B1(new_n750), .B2(G45), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n705), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n749), .B(new_n754), .C1(G330), .C2(new_n691), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n220), .A2(G355), .A3(new_n307), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(G116), .B2(new_n220), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n220), .A2(new_n302), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(new_n473), .B2(new_n228), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n245), .A2(G45), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n757), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n223), .B1(G20), .B2(new_n276), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT98), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n753), .B1(new_n761), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n224), .A2(G179), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G190), .A2(G200), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n307), .B1(new_n772), .B2(G329), .ZN(new_n773));
  INV_X1    g0573(.A(G283), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n769), .A2(new_n339), .A3(G200), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n339), .A2(G200), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n224), .A2(new_n272), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n778), .A2(KEYINPUT99), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(KEYINPUT99), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n777), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n776), .B1(new_n782), .B2(G322), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n778), .A2(G200), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(G190), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  XOR2_X1   g0586(.A(KEYINPUT33), .B(G317), .Z(new_n787));
  NOR2_X1   g0587(.A1(new_n784), .A2(new_n339), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G326), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n786), .A2(new_n787), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n777), .A2(new_n272), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G294), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n769), .A2(G190), .A3(G200), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n794), .A2(new_n795), .B1(new_n796), .B2(new_n637), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n791), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G311), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n770), .B1(new_n779), .B2(new_n780), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n783), .B(new_n798), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n800), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G58), .A2(new_n782), .B1(new_n802), .B2(G77), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n796), .A2(new_n210), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n307), .B1(new_n775), .B2(new_n396), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n804), .B(new_n805), .C1(G68), .C2(new_n785), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n794), .A2(new_n486), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(G50), .B2(new_n788), .ZN(new_n808));
  INV_X1    g0608(.A(G159), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n771), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT32), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n803), .A2(new_n806), .A3(new_n808), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n801), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n768), .B1(new_n813), .B2(new_n765), .ZN(new_n814));
  INV_X1    g0614(.A(new_n764), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n814), .B1(new_n691), .B2(new_n815), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n755), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(G396));
  NAND2_X1  g0618(.A1(new_n665), .A2(new_n686), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n403), .A2(new_n685), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n408), .B1(new_n393), .B2(new_n686), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n403), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n819), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n824), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n566), .B(new_n657), .C1(new_n716), .C2(new_n656), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n572), .A2(new_n661), .A3(new_n663), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n686), .B(new_n826), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n746), .B1(new_n825), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(new_n753), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n825), .A2(new_n746), .A3(new_n829), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n765), .A2(new_n762), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n754), .B1(new_n353), .B2(new_n834), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n307), .B(new_n807), .C1(G311), .C2(new_n772), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n836), .B1(new_n795), .B2(new_n781), .C1(new_n629), .C2(new_n800), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n210), .A2(new_n775), .B1(new_n796), .B2(new_n396), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n786), .A2(new_n774), .B1(new_n789), .B2(new_n637), .ZN(new_n839));
  NOR3_X1   g0639(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G137), .A2(new_n788), .B1(new_n785), .B2(G150), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT100), .ZN(new_n842));
  INV_X1    g0642(.A(G143), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n842), .B1(new_n843), .B2(new_n781), .C1(new_n809), .C2(new_n800), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT34), .ZN(new_n845));
  INV_X1    g0645(.A(G132), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n307), .B1(new_n771), .B2(new_n846), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n202), .A2(new_n796), .B1(new_n775), .B2(new_n208), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n847), .B(new_n848), .C1(G58), .C2(new_n793), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n840), .B1(new_n845), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n765), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n835), .B1(new_n826), .B2(new_n763), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n833), .A2(new_n852), .ZN(G384));
  OR2_X1    g0653(.A1(new_n491), .A2(KEYINPUT35), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n491), .A2(KEYINPUT35), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n854), .A2(G116), .A3(new_n225), .A4(new_n855), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT36), .Z(new_n857));
  OR3_X1    g0657(.A1(new_n227), .A2(new_n353), .A3(new_n312), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n202), .A2(G68), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n254), .B(G13), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n678), .B1(new_n726), .B2(new_n456), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT106), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n208), .B1(new_n308), .B2(new_n327), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n300), .B1(new_n864), .B2(new_n316), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n320), .A2(new_n865), .A3(new_n321), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n326), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT102), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n683), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n326), .A2(new_n866), .A3(KEYINPUT102), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n869), .A2(new_n325), .A3(new_n871), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n872), .A2(new_n873), .A3(new_n342), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(KEYINPUT37), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n325), .A2(new_n334), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n334), .A2(new_n870), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT37), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n876), .A2(new_n877), .A3(new_n878), .A4(new_n342), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n879), .A2(KEYINPUT103), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n879), .A2(KEYINPUT103), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n875), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  INV_X1    g0683(.A(new_n872), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n883), .B1(new_n346), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n325), .A2(new_n334), .A3(new_n335), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n335), .B1(new_n325), .B2(new_n334), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n872), .B1(new_n889), .B2(new_n669), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n317), .A2(new_n322), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n891), .A2(new_n326), .B1(new_n275), .B2(new_n282), .ZN(new_n892));
  INV_X1    g0692(.A(new_n342), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT103), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n894), .A2(new_n895), .A3(new_n878), .A4(new_n877), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n879), .A2(KEYINPUT103), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n890), .B1(new_n898), .B2(new_n875), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n886), .B1(new_n899), .B2(KEYINPUT38), .ZN(new_n900));
  XOR2_X1   g0700(.A(new_n820), .B(KEYINPUT101), .Z(new_n901));
  NAND2_X1  g0701(.A1(new_n829), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n454), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n450), .B(new_n685), .C1(new_n903), .C2(new_n437), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n450), .A2(new_n685), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n451), .A2(new_n454), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n900), .A2(new_n902), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n667), .A2(new_n683), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(KEYINPUT104), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT39), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n896), .A2(new_n897), .B1(KEYINPUT37), .B2(new_n874), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n346), .A2(new_n884), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT38), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n912), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n876), .A2(new_n877), .A3(new_n342), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(KEYINPUT37), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n880), .B2(new_n881), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n346), .A2(new_n334), .A3(new_n870), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT38), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT105), .B1(new_n916), .B2(new_n921), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n896), .A2(new_n897), .B1(KEYINPUT37), .B2(new_n917), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n347), .A2(new_n877), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n883), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT105), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n925), .A2(new_n926), .A3(new_n912), .A4(new_n886), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT38), .B1(new_n882), .B2(new_n914), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n913), .A2(new_n915), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT39), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n922), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n451), .A2(new_n685), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT104), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n908), .A2(new_n934), .A3(new_n909), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n911), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n863), .B(new_n936), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n685), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT31), .B1(new_n735), .B2(new_n685), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n653), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n694), .A2(new_n941), .A3(new_n686), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n940), .B1(new_n574), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n824), .B1(new_n904), .B2(new_n906), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n943), .B(new_n944), .C1(new_n928), .C2(new_n929), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT40), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n925), .A2(new_n886), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n948), .A2(KEYINPUT40), .A3(new_n943), .A4(new_n944), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n943), .A2(new_n456), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n951), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n952), .A2(G330), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n937), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n254), .B2(new_n750), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n937), .A2(new_n954), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n861), .B1(new_n956), .B2(new_n957), .ZN(G367));
  INV_X1    g0758(.A(new_n767), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n220), .B2(new_n551), .ZN(new_n960));
  AND3_X1   g0760(.A1(new_n237), .A2(new_n220), .A3(new_n302), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n753), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n775), .A2(new_n486), .ZN(new_n963));
  NAND2_X1  g0763(.A1(KEYINPUT46), .A2(G116), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n786), .A2(new_n795), .B1(new_n796), .B2(new_n964), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n963), .B(new_n965), .C1(G107), .C2(new_n793), .ZN(new_n966));
  INV_X1    g0766(.A(G317), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n302), .B1(new_n771), .B2(new_n967), .C1(new_n789), .C2(new_n799), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(new_n782), .B2(G303), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n802), .A2(G283), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT46), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n629), .B2(new_n796), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n966), .A2(new_n969), .A3(new_n970), .A4(new_n972), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n786), .A2(new_n809), .B1(new_n789), .B2(new_n843), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n793), .A2(G68), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n353), .B2(new_n775), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(G137), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n307), .B1(new_n771), .B2(new_n978), .C1(new_n311), .C2(new_n796), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(new_n802), .B2(G50), .ZN(new_n980));
  INV_X1    g0780(.A(G150), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n977), .B(new_n980), .C1(new_n981), .C2(new_n781), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n973), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT47), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n962), .B1(new_n984), .B2(new_n765), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n541), .A2(new_n552), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n685), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n567), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n566), .B2(new_n987), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n985), .B1(new_n989), .B2(new_n815), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n705), .B(KEYINPUT41), .Z(new_n991));
  NAND2_X1  g0791(.A1(new_n696), .A2(new_n699), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n623), .B2(new_n699), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n993), .A2(new_n692), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n994), .B1(new_n749), .B2(new_n993), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n747), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n516), .B(new_n522), .C1(new_n518), .C2(new_n686), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n655), .A2(new_n685), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n702), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT45), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1002), .B(new_n1003), .ZN(new_n1004));
  AND2_X1   g0804(.A1(new_n999), .A2(new_n1000), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n700), .B2(new_n701), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT44), .ZN(new_n1007));
  AND2_X1   g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1004), .B(new_n698), .C1(new_n1008), .C2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1004), .B1(new_n1010), .B2(new_n1008), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n697), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n998), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n991), .B1(new_n1014), .B2(new_n747), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1015), .A2(new_n752), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1001), .A2(new_n700), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT42), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n516), .B1(new_n1005), .B2(new_n722), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n686), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n989), .A2(KEYINPUT43), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1022), .A2(KEYINPUT107), .A3(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1019), .A2(new_n1023), .A3(new_n1021), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT107), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n989), .B(KEYINPUT43), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1024), .B(new_n1027), .C1(new_n1022), .C2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n697), .A2(new_n1001), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1029), .B(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n990), .B1(new_n1016), .B2(new_n1031), .ZN(G387));
  INV_X1    g0832(.A(new_n998), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n996), .A2(new_n997), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1033), .A2(new_n705), .A3(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n794), .A2(new_n551), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n782), .B2(G50), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT109), .Z(new_n1038));
  AOI211_X1 g0838(.A(new_n302), .B(new_n963), .C1(G159), .C2(new_n788), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n802), .A2(G68), .B1(new_n292), .B2(new_n785), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n796), .A2(new_n353), .B1(new_n771), .B2(new_n981), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT108), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .A4(new_n1042), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G311), .A2(new_n785), .B1(new_n788), .B2(G322), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n637), .B2(new_n800), .C1(new_n967), .C2(new_n781), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT48), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n796), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G294), .A2(new_n1049), .B1(new_n793), .B2(G283), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1047), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT49), .Z(new_n1052));
  OAI221_X1 g0852(.A(new_n302), .B1(new_n771), .B2(new_n790), .C1(new_n629), .C2(new_n775), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1043), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n765), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n234), .A2(G45), .A3(new_n302), .ZN(new_n1056));
  OAI21_X1  g0856(.A(KEYINPUT50), .B1(new_n285), .B2(G50), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1057), .B(new_n473), .C1(new_n208), .C2(new_n353), .ZN(new_n1058));
  NOR3_X1   g0858(.A1(new_n285), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n302), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n706), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n704), .B1(new_n1056), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n959), .B1(new_n396), .B2(new_n220), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1055), .B(new_n753), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n696), .B2(new_n764), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT110), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1035), .B(new_n1067), .C1(new_n751), .C2(new_n996), .ZN(G393));
  NAND3_X1  g0868(.A1(new_n1013), .A2(new_n1011), .A3(new_n752), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n782), .A2(G311), .B1(G317), .B2(new_n788), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT52), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n796), .A2(new_n774), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n786), .A2(new_n637), .B1(new_n794), .B2(new_n629), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n307), .B1(new_n772), .B2(G322), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1074), .B1(new_n396), .B2(new_n775), .C1(new_n800), .C2(new_n795), .ZN(new_n1075));
  OR4_X1    g0875(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .A4(new_n1075), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n781), .A2(new_n809), .B1(new_n789), .B2(new_n981), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT51), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n786), .A2(new_n202), .B1(new_n794), .B2(new_n353), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(G68), .B2(new_n1049), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n307), .B1(new_n771), .B2(new_n843), .C1(new_n210), .C2(new_n775), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n285), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1081), .B1(new_n802), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1078), .A2(new_n1080), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n851), .B1(new_n1076), .B2(new_n1084), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n242), .A2(new_n758), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n767), .B1(G97), .B2(new_n704), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n754), .B(new_n1085), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n1001), .B2(new_n815), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1069), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(KEYINPUT111), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT111), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1069), .A2(new_n1092), .A3(new_n1089), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1013), .A2(new_n1011), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1033), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1096), .A2(new_n1014), .A3(new_n705), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1094), .A2(new_n1097), .ZN(G390));
  AOI21_X1  g0898(.A(new_n932), .B1(new_n902), .B2(new_n907), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n907), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n719), .A2(new_n724), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1101), .A2(new_n686), .A3(new_n823), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1100), .B1(new_n1102), .B2(new_n821), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n932), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n948), .A2(new_n1104), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n931), .A2(new_n1099), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n943), .A2(G330), .A3(new_n944), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n820), .B1(new_n725), .B2(new_n823), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1104), .B(new_n948), .C1(new_n1109), .C2(new_n1100), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n746), .A2(new_n826), .A3(new_n907), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1110), .B(new_n1111), .C1(new_n931), .C2(new_n1099), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1108), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n907), .B1(new_n746), .B2(new_n826), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n902), .B1(new_n1114), .B2(new_n1107), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n943), .A2(G330), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1100), .B1(new_n1116), .B2(new_n824), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1117), .A2(new_n1111), .A3(new_n1109), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  AND3_X1   g0919(.A1(new_n943), .A2(G330), .A3(new_n456), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n678), .B(new_n1120), .C1(new_n726), .C2(new_n456), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1113), .A2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1108), .A2(new_n1112), .A3(new_n1121), .A4(new_n1119), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1123), .A2(new_n705), .A3(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1108), .A2(new_n752), .A3(new_n1112), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n834), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n753), .B1(new_n292), .B2(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT112), .ZN(new_n1129));
  INV_X1    g0929(.A(G128), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n789), .A2(new_n1130), .B1(new_n794), .B2(new_n809), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(G137), .B2(new_n785), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n302), .B1(new_n772), .B2(G125), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n202), .B2(new_n775), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(new_n782), .B2(G132), .ZN(new_n1135));
  XOR2_X1   g0935(.A(KEYINPUT54), .B(G143), .Z(new_n1136));
  NAND2_X1  g0936(.A1(new_n802), .A2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n796), .A2(new_n981), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT53), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1132), .A2(new_n1135), .A3(new_n1137), .A4(new_n1139), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n802), .A2(G97), .B1(G107), .B2(new_n785), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1141), .A2(KEYINPUT113), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n781), .A2(new_n624), .B1(new_n794), .B2(new_n353), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1142), .B1(KEYINPUT114), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1144), .B1(KEYINPUT114), .B2(new_n1143), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1141), .A2(KEYINPUT113), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n307), .B(new_n804), .C1(G294), .C2(new_n772), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n775), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n788), .A2(G283), .B1(new_n1148), .B2(G68), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1146), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1140), .B1(new_n1145), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1129), .B1(new_n1151), .B2(new_n765), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n931), .B2(new_n763), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1125), .A2(new_n1126), .A3(new_n1153), .ZN(G378));
  NAND3_X1  g0954(.A1(new_n947), .A2(G330), .A3(new_n949), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT117), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n404), .A2(new_n683), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n676), .B2(new_n406), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n412), .A2(new_n386), .A3(KEYINPUT93), .ZN(new_n1162));
  AOI21_X1  g0962(.A(KEYINPUT93), .B1(new_n412), .B2(new_n386), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n406), .B(new_n1160), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1158), .B1(new_n1161), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n406), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n1159), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1168), .A2(new_n1164), .A3(new_n1157), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1155), .A2(new_n1156), .A3(new_n1170), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n1166), .A2(KEYINPUT116), .A3(new_n1169), .ZN(new_n1172));
  AOI21_X1  g0972(.A(KEYINPUT116), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1174), .A2(G330), .A3(new_n947), .A4(new_n949), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1171), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1156), .B1(new_n1155), .B2(new_n1170), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n936), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1155), .A2(new_n1170), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(KEYINPUT117), .ZN(new_n1180));
  AND3_X1   g0980(.A1(new_n911), .A2(new_n933), .A3(new_n935), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1180), .A2(new_n1181), .A3(new_n1175), .A4(new_n1171), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1178), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT57), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n1124), .B2(new_n1121), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1178), .A2(new_n1182), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n705), .C1(KEYINPUT57), .C2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n753), .B1(G50), .B2(new_n1127), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1174), .A2(new_n763), .ZN(new_n1190));
  AOI211_X1 g0990(.A(G41), .B(new_n307), .C1(new_n772), .C2(G283), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1191), .B1(new_n311), .B2(new_n775), .C1(new_n353), .C2(new_n796), .ZN(new_n1192));
  XOR2_X1   g0992(.A(new_n1192), .B(KEYINPUT115), .Z(new_n1193));
  OAI221_X1 g0993(.A(new_n975), .B1(new_n789), .B2(new_n624), .C1(new_n486), .C2(new_n786), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n396), .A2(new_n781), .B1(new_n800), .B2(new_n551), .ZN(new_n1195));
  NOR3_X1   g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT58), .Z(new_n1197));
  AOI21_X1  g0997(.A(G50), .B1(new_n261), .B2(new_n470), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n307), .B2(G41), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G128), .A2(new_n782), .B1(new_n802), .B2(G137), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n788), .A2(G125), .B1(new_n793), .B2(G150), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n785), .A2(G132), .B1(new_n1049), .B2(new_n1136), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1204), .A2(KEYINPUT59), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(KEYINPUT59), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1148), .A2(G159), .ZN(new_n1207));
  AOI211_X1 g1007(.A(G33), .B(G41), .C1(new_n772), .C2(G124), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1197), .B(new_n1199), .C1(new_n1205), .C2(new_n1209), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1189), .B(new_n1190), .C1(new_n765), .C2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n1183), .B2(new_n752), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1188), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT118), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1213), .B(new_n1214), .ZN(G375));
  NAND2_X1  g1015(.A1(new_n1119), .A2(new_n752), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n753), .B1(G68), .B2(new_n1127), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n629), .A2(new_n786), .B1(new_n789), .B2(new_n795), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1036), .B(new_n1218), .C1(G97), .C2(new_n1049), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n302), .B1(new_n771), .B2(new_n637), .C1(new_n353), .C2(new_n775), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n782), .B2(G283), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1219), .B(new_n1221), .C1(new_n396), .C2(new_n800), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n307), .B1(new_n771), .B2(new_n1130), .C1(new_n311), .C2(new_n775), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n794), .A2(new_n202), .B1(new_n796), .B2(new_n809), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(G150), .C2(new_n802), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT120), .Z(new_n1226));
  AOI22_X1  g1026(.A1(G132), .A2(new_n788), .B1(new_n785), .B2(new_n1136), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n978), .B2(new_n781), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT119), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1222), .B1(new_n1226), .B2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1217), .B1(new_n1230), .B2(new_n765), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n907), .B2(new_n763), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1216), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n862), .B1(new_n457), .B2(new_n1116), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1235), .A2(new_n1115), .A3(new_n1118), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n991), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1122), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1234), .A2(new_n1238), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(KEYINPUT121), .ZN(G381));
  NOR4_X1   g1040(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1031), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(new_n1015), .B2(new_n752), .ZN(new_n1243));
  INV_X1    g1043(.A(G378), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1241), .A2(new_n1243), .A3(new_n990), .A4(new_n1244), .ZN(new_n1245));
  OR3_X1    g1045(.A1(new_n1245), .A2(G375), .A3(G381), .ZN(G407));
  INV_X1    g1046(.A(G213), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1247), .A2(G343), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(G375), .A2(G378), .A3(new_n1249), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT122), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1251), .A2(G213), .A3(G407), .ZN(G409));
  NAND2_X1  g1052(.A1(new_n1186), .A2(new_n705), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1124), .A2(new_n1121), .ZN(new_n1254));
  AOI21_X1  g1054(.A(KEYINPUT57), .B1(new_n1183), .B2(new_n1254), .ZN(new_n1255));
  OAI211_X1 g1055(.A(G378), .B(new_n1212), .C1(new_n1253), .C2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT123), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1188), .A2(KEYINPUT123), .A3(G378), .A4(new_n1212), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1187), .A2(new_n1237), .ZN(new_n1261));
  AOI21_X1  g1061(.A(G378), .B1(new_n1261), .B2(new_n1212), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1260), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(G384), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1122), .A2(new_n705), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT124), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT60), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1267), .B(KEYINPUT60), .C1(new_n1119), .C2(new_n1121), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1266), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1265), .B1(new_n1272), .B2(new_n1233), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1266), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1271), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT60), .B1(new_n1236), .B2(new_n1267), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1274), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1277), .A2(G384), .A3(new_n1234), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1273), .A2(new_n1278), .A3(KEYINPUT125), .ZN(new_n1279));
  AOI21_X1  g1079(.A(KEYINPUT125), .B1(new_n1273), .B2(new_n1278), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT63), .ZN(new_n1281));
  NOR3_X1   g1081(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1264), .A2(new_n1249), .A3(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1248), .A2(G2897), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1284), .B1(new_n1273), .B2(new_n1278), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1285), .B1(new_n1286), .B2(new_n1284), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1262), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1287), .B1(new_n1288), .B2(new_n1248), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT61), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(G387), .A2(new_n1094), .A3(new_n1097), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1243), .A2(G390), .A3(new_n990), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(G393), .B(new_n817), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1291), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1293), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1283), .A2(new_n1289), .A3(new_n1290), .A4(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1288), .A2(new_n1248), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT63), .B1(new_n1299), .B2(new_n1286), .ZN(new_n1300));
  OAI21_X1  g1100(.A(KEYINPUT126), .B1(new_n1298), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1264), .A2(new_n1249), .ZN(new_n1302));
  AOI21_X1  g1102(.A(KEYINPUT61), .B1(new_n1302), .B2(new_n1287), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1293), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1294), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1307), .B1(new_n1299), .B2(new_n1282), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1264), .A2(new_n1249), .A3(new_n1286), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1281), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT126), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1303), .A2(new_n1308), .A3(new_n1310), .A4(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1301), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT127), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1309), .A2(new_n1314), .A3(KEYINPUT62), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n1303), .ZN(new_n1316));
  XOR2_X1   g1116(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1317));
  NOR2_X1   g1117(.A1(new_n1309), .A2(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1307), .B1(new_n1316), .B2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1313), .A2(new_n1319), .ZN(G405));
  NAND2_X1  g1120(.A1(G375), .A2(new_n1244), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1273), .A2(new_n1278), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1321), .A2(new_n1260), .A3(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1286), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1324), .B1(new_n1321), .B2(new_n1260), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1323), .A2(new_n1325), .ZN(new_n1326));
  XNOR2_X1  g1126(.A(new_n1326), .B(new_n1297), .ZN(G402));
endmodule


