//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 1 1 1 0 1 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n569, new_n571, new_n572, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n626, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1240;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT64), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n462), .B1(new_n463), .B2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(KEYINPUT64), .A3(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(G101), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT65), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT65), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n464), .A2(new_n466), .A3(new_n469), .A4(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n472), .A2(new_n474), .A3(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n472), .A2(new_n474), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G137), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n471), .A2(new_n478), .A3(new_n481), .ZN(G160));
  OAI21_X1  g057(.A(KEYINPUT66), .B1(new_n479), .B2(new_n465), .ZN(new_n483));
  XNOR2_X1  g058(.A(KEYINPUT3), .B(G2104), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT66), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n484), .A2(new_n485), .A3(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  AOI22_X1  g062(.A1(new_n487), .A2(G124), .B1(G136), .B2(new_n480), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT67), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n488), .A2(new_n493), .A3(new_n490), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(G162));
  NAND4_X1  g070(.A1(new_n472), .A2(new_n474), .A3(G138), .A4(new_n465), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AND3_X1   g073(.A1(new_n465), .A2(KEYINPUT4), .A3(G138), .ZN(new_n499));
  AND2_X1   g074(.A1(G126), .A2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n484), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT68), .B1(new_n465), .B2(G114), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT68), .ZN(new_n503));
  INV_X1    g078(.A(G114), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(new_n504), .A3(G2105), .ZN(new_n505));
  OR2_X1    g080(.A1(G102), .A2(G2105), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n502), .A2(new_n505), .A3(G2104), .A4(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n498), .A2(new_n501), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n510));
  AND3_X1   g085(.A1(KEYINPUT69), .A2(KEYINPUT6), .A3(G651), .ZN(new_n511));
  AOI21_X1  g086(.A(KEYINPUT6), .B1(KEYINPUT69), .B2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n510), .B1(new_n513), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT69), .A2(G651), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT6), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(KEYINPUT69), .A2(KEYINPUT6), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT5), .B(G543), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n524), .A2(KEYINPUT70), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n519), .A2(G88), .A3(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n513), .A2(new_n514), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G50), .ZN(new_n529));
  INV_X1    g104(.A(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(G75), .A2(G543), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(KEYINPUT71), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT71), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n533), .A2(G75), .A3(G543), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n515), .A2(new_n517), .A3(G62), .ZN(new_n536));
  AOI211_X1 g111(.A(KEYINPUT72), .B(new_n530), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT72), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n536), .A2(new_n532), .A3(new_n534), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n538), .B1(new_n539), .B2(G651), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n527), .B(new_n529), .C1(new_n537), .C2(new_n540), .ZN(G303));
  INV_X1    g116(.A(G303), .ZN(G166));
  NAND3_X1  g117(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT73), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n528), .A2(G51), .ZN(new_n545));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT7), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n519), .A2(G89), .A3(new_n526), .ZN(new_n548));
  NAND4_X1  g123(.A1(new_n544), .A2(new_n545), .A3(new_n547), .A4(new_n548), .ZN(G286));
  INV_X1    g124(.A(G286), .ZN(G168));
  NAND2_X1  g125(.A1(G77), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G64), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n518), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(G52), .A2(new_n528), .B1(new_n553), .B2(G651), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n519), .A2(G90), .A3(new_n526), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(G301));
  INV_X1    g131(.A(G301), .ZN(G171));
  NAND3_X1  g132(.A1(new_n519), .A2(G81), .A3(new_n526), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n528), .A2(G43), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n558), .A2(KEYINPUT74), .A3(new_n559), .ZN(new_n563));
  NAND2_X1  g138(.A1(G68), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G56), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n518), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n562), .A2(new_n563), .B1(G651), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  AND3_X1   g143(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G36), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n569), .A2(new_n572), .ZN(G188));
  OAI211_X1 g148(.A(G53), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n524), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(KEYINPUT75), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT75), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n576), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n519), .A2(G91), .A3(new_n526), .ZN(new_n583));
  NAND2_X1  g158(.A1(G78), .A2(G543), .ZN(new_n584));
  XOR2_X1   g159(.A(KEYINPUT76), .B(G65), .Z(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n585), .B2(new_n518), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G651), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n582), .A2(new_n589), .ZN(G299));
  NAND3_X1  g165(.A1(new_n519), .A2(G87), .A3(new_n526), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n528), .A2(G49), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(G288));
  NAND3_X1  g169(.A1(new_n519), .A2(G86), .A3(new_n526), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT77), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n528), .A2(new_n596), .A3(G48), .ZN(new_n597));
  NAND2_X1  g172(.A1(G73), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G61), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n518), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G651), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n524), .A2(G48), .A3(G543), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(KEYINPUT77), .ZN(new_n603));
  NAND4_X1  g178(.A1(new_n595), .A2(new_n597), .A3(new_n601), .A4(new_n603), .ZN(G305));
  AND2_X1   g179(.A1(new_n519), .A2(new_n526), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G85), .ZN(new_n606));
  NAND2_X1  g181(.A1(G72), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G60), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n518), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(G47), .A2(new_n528), .B1(new_n609), .B2(G651), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n606), .A2(new_n610), .ZN(G290));
  NAND2_X1  g186(.A1(G301), .A2(G868), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n605), .A2(new_n613), .A3(G92), .ZN(new_n614));
  NAND2_X1  g189(.A1(G79), .A2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G66), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n518), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(G54), .A2(new_n528), .B1(new_n617), .B2(G651), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n519), .A2(new_n526), .ZN(new_n619));
  INV_X1    g194(.A(G92), .ZN(new_n620));
  OAI21_X1  g195(.A(KEYINPUT10), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AND3_X1   g196(.A1(new_n614), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n612), .B1(new_n622), .B2(G868), .ZN(G284));
  OAI21_X1  g198(.A(new_n612), .B1(new_n622), .B2(G868), .ZN(G321));
  NAND2_X1  g199(.A1(G286), .A2(G868), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n588), .B1(new_n579), .B2(new_n581), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G868), .ZN(G297));
  OAI21_X1  g202(.A(new_n625), .B1(new_n626), .B2(G868), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n622), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND2_X1  g205(.A1(new_n566), .A2(G651), .ZN(new_n631));
  INV_X1    g206(.A(new_n563), .ZN(new_n632));
  AOI21_X1  g207(.A(KEYINPUT74), .B1(new_n558), .B2(new_n559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(G868), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n622), .A2(new_n629), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n636), .B1(new_n638), .B2(new_n635), .ZN(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g215(.A1(new_n464), .A2(new_n466), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(new_n484), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT12), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT13), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2100), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n487), .A2(G123), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n480), .A2(G135), .ZN(new_n647));
  NOR2_X1   g222(.A1(G99), .A2(G2105), .ZN(new_n648));
  OAI21_X1  g223(.A(G2104), .B1(new_n465), .B2(G111), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n646), .B(new_n647), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(G2096), .Z(new_n651));
  NAND2_X1  g226(.A1(new_n645), .A2(new_n651), .ZN(G156));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2430), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2435), .ZN(new_n654));
  XOR2_X1   g229(.A(G2427), .B(G2438), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(KEYINPUT14), .ZN(new_n657));
  XOR2_X1   g232(.A(G2451), .B(G2454), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n659), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n663), .B(new_n664), .Z(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(G14), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(G401));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  XOR2_X1   g243(.A(G2067), .B(G2678), .Z(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2084), .B(G2090), .Z(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n668), .B1(new_n672), .B2(KEYINPUT18), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT80), .ZN(new_n674));
  XOR2_X1   g249(.A(G2096), .B(G2100), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n670), .A2(new_n671), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT79), .B(KEYINPUT17), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n670), .B2(new_n671), .ZN(new_n679));
  AOI21_X1  g254(.A(KEYINPUT18), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n676), .B(new_n680), .ZN(G227));
  XOR2_X1   g256(.A(G1956), .B(G2474), .Z(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1971), .B(G1976), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n682), .A2(new_n683), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT20), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n688), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n685), .A2(new_n687), .A3(new_n689), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n692), .B(new_n693), .C1(new_n691), .C2(new_n690), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT21), .B(G1986), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(G1991), .B(G1996), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT22), .B(G1981), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(G229));
  OR2_X1    g275(.A1(G16), .A2(G21), .ZN(new_n701));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n701), .B1(G286), .B2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT92), .ZN(new_n704));
  INV_X1    g279(.A(G1966), .ZN(new_n705));
  OR3_X1    g280(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n704), .B1(new_n703), .B2(new_n705), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G26), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n487), .A2(G128), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n480), .A2(G140), .ZN(new_n712));
  OAI21_X1  g287(.A(G2104), .B1(new_n465), .B2(G116), .ZN(new_n713));
  NOR2_X1   g288(.A1(G104), .A2(G2105), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT86), .Z(new_n715));
  OAI21_X1  g290(.A(new_n712), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(G29), .B1(new_n711), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(new_n710), .ZN(new_n718));
  MUX2_X1   g293(.A(new_n710), .B(new_n718), .S(KEYINPUT28), .Z(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G2067), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n709), .B1(new_n492), .B2(new_n494), .ZN(new_n721));
  NOR2_X1   g296(.A1(G29), .A2(G35), .ZN(new_n722));
  OAI21_X1  g297(.A(KEYINPUT29), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n494), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n493), .B1(new_n488), .B2(new_n490), .ZN(new_n725));
  OAI21_X1  g300(.A(G29), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT29), .ZN(new_n727));
  INV_X1    g302(.A(new_n722), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(G2090), .B1(new_n723), .B2(new_n729), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n708), .B(new_n720), .C1(new_n730), .C2(KEYINPUT95), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n719), .A2(G2067), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n487), .A2(G129), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT90), .ZN(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT26), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n641), .A2(G105), .ZN(new_n738));
  AOI211_X1 g313(.A(new_n737), .B(new_n738), .C1(G141), .C2(new_n480), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n735), .A2(G29), .A3(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT91), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G29), .B2(G32), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n741), .B2(new_n740), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT27), .B(G1996), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n746), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n744), .B(new_n748), .C1(new_n741), .C2(new_n740), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n702), .A2(G4), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n622), .B2(new_n702), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n752), .A2(G1348), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n752), .A2(G1348), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G34), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(new_n709), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n471), .A2(new_n478), .A3(new_n481), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n758), .B2(new_n709), .ZN(new_n759));
  INV_X1    g334(.A(G2084), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR3_X1   g336(.A1(new_n753), .A2(new_n754), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n759), .A2(new_n760), .ZN(new_n763));
  AND3_X1   g338(.A1(new_n750), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n702), .A2(G5), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G171), .B2(new_n702), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G1961), .ZN(new_n767));
  AND2_X1   g342(.A1(KEYINPUT81), .A2(G16), .ZN(new_n768));
  NOR2_X1   g343(.A1(KEYINPUT81), .A2(G16), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n771), .A2(KEYINPUT23), .A3(G20), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT23), .ZN(new_n773));
  INV_X1    g348(.A(G20), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n770), .B2(new_n774), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n772), .B(new_n775), .C1(new_n626), .C2(new_n702), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G1956), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n767), .B(new_n777), .C1(new_n730), .C2(KEYINPUT95), .ZN(new_n778));
  OR2_X1    g353(.A1(G29), .A2(G33), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT87), .Z(new_n781));
  OR2_X1    g356(.A1(new_n781), .A2(KEYINPUT25), .ZN(new_n782));
  NAND2_X1  g357(.A1(G115), .A2(G2104), .ZN(new_n783));
  INV_X1    g358(.A(G127), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n479), .B2(new_n784), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n785), .A2(G2105), .B1(new_n480), .B2(G139), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n781), .A2(KEYINPUT25), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n782), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  OAI211_X1 g363(.A(G2072), .B(new_n779), .C1(new_n788), .C2(new_n709), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT89), .Z(new_n790));
  NAND2_X1  g365(.A1(new_n709), .A2(G27), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G164), .B2(new_n709), .ZN(new_n792));
  INV_X1    g367(.A(G2078), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n650), .A2(new_n709), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT30), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n709), .B1(new_n796), .B2(G28), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT93), .Z(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n796), .B2(G28), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n779), .B1(new_n788), .B2(new_n709), .ZN(new_n800));
  INV_X1    g375(.A(G2072), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n790), .A2(new_n794), .A3(new_n795), .A4(new_n802), .ZN(new_n803));
  AND3_X1   g378(.A1(new_n723), .A2(G2090), .A3(new_n729), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n733), .A2(new_n764), .A3(new_n778), .A4(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT36), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n807), .A2(KEYINPUT85), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n771), .A2(G24), .ZN(new_n809));
  INV_X1    g384(.A(G290), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n810), .B2(new_n771), .ZN(new_n811));
  INV_X1    g386(.A(G1986), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n487), .A2(G119), .B1(G131), .B2(new_n480), .ZN(new_n815));
  OR2_X1    g390(.A1(G95), .A2(G2105), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n816), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(new_n709), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G25), .B2(new_n709), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT35), .B(G1991), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n821), .B(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(G16), .A2(G23), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(G288), .A2(KEYINPUT83), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT83), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n591), .A2(new_n828), .A3(new_n592), .A4(new_n593), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n826), .B1(new_n831), .B2(new_n702), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT33), .B(G1976), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT84), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n834), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n836), .B(new_n826), .C1(new_n831), .C2(new_n702), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n771), .A2(G22), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(G166), .B2(new_n771), .ZN(new_n839));
  INV_X1    g414(.A(G1971), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI211_X1 g416(.A(G1971), .B(new_n838), .C1(G166), .C2(new_n771), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AND3_X1   g418(.A1(new_n835), .A2(new_n837), .A3(new_n843), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT32), .B(G1981), .Z(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(G305), .A2(G16), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT82), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n702), .A2(G6), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n848), .B1(new_n847), .B2(new_n849), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n846), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n852), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n854), .A2(new_n845), .A3(new_n850), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n844), .A2(KEYINPUT34), .A3(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT34), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n835), .A2(new_n837), .A3(new_n843), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n859), .B1(new_n860), .B2(new_n856), .ZN(new_n861));
  AOI211_X1 g436(.A(new_n814), .B(new_n824), .C1(new_n858), .C2(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n806), .B1(new_n808), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n771), .A2(G19), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n567), .B2(new_n771), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(G1341), .Z(new_n866));
  XNOR2_X1  g441(.A(KEYINPUT31), .B(G11), .ZN(new_n867));
  INV_X1    g442(.A(new_n824), .ZN(new_n868));
  AOI21_X1  g443(.A(KEYINPUT34), .B1(new_n844), .B2(new_n857), .ZN(new_n869));
  NOR3_X1   g444(.A1(new_n860), .A2(new_n856), .A3(new_n859), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n813), .B(new_n868), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n808), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n807), .A2(KEYINPUT85), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n863), .A2(new_n866), .A3(new_n867), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n703), .A2(new_n705), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(KEYINPUT94), .Z(new_n877));
  NOR2_X1   g452(.A1(new_n875), .A2(new_n877), .ZN(G311));
  INV_X1    g453(.A(KEYINPUT96), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n879), .B1(new_n875), .B2(new_n877), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n862), .A2(new_n808), .ZN(new_n881));
  INV_X1    g456(.A(new_n806), .ZN(new_n882));
  AND4_X1   g457(.A1(new_n867), .A2(new_n881), .A3(new_n874), .A4(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n877), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n883), .A2(KEYINPUT96), .A3(new_n884), .A4(new_n866), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n880), .A2(new_n885), .ZN(G150));
  NAND2_X1  g461(.A1(new_n605), .A2(G93), .ZN(new_n887));
  NAND2_X1  g462(.A1(G80), .A2(G543), .ZN(new_n888));
  INV_X1    g463(.A(G67), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n888), .B1(new_n518), .B2(new_n889), .ZN(new_n890));
  AOI22_X1  g465(.A1(G55), .A2(new_n528), .B1(new_n890), .B2(G651), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(G860), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n893), .B(KEYINPUT37), .Z(new_n894));
  NAND3_X1  g469(.A1(new_n614), .A2(new_n618), .A3(new_n621), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n895), .A2(new_n629), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT98), .ZN(new_n897));
  XNOR2_X1  g472(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n897), .B(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n634), .A2(new_n887), .A3(new_n891), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n567), .A2(new_n892), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT39), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n899), .B(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n894), .B1(new_n904), .B2(G860), .ZN(G145));
  NOR2_X1   g480(.A1(new_n711), .A2(new_n716), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(new_n508), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n735), .A2(new_n739), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n907), .B(new_n908), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n909), .A2(new_n788), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n788), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI22_X1  g487(.A1(new_n487), .A2(G130), .B1(G142), .B2(new_n480), .ZN(new_n913));
  OR2_X1    g488(.A1(G106), .A2(G2105), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n914), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(new_n643), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(new_n818), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(KEYINPUT99), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n912), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n910), .A2(new_n911), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n919), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n650), .B(G160), .ZN(new_n925));
  XOR2_X1   g500(.A(new_n925), .B(G162), .Z(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(G37), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n922), .A2(new_n918), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n921), .A2(new_n926), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g507(.A(KEYINPUT100), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n902), .A2(new_n638), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n900), .A2(new_n901), .A3(new_n637), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n622), .A2(new_n626), .ZN(new_n937));
  NAND2_X1  g512(.A1(G299), .A2(new_n895), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n936), .A2(new_n940), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n937), .A2(KEYINPUT41), .A3(new_n938), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT41), .B1(new_n937), .B2(new_n938), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n944), .A2(new_n935), .A3(new_n934), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n933), .B1(new_n941), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT100), .B1(new_n936), .B2(new_n940), .ZN(new_n947));
  OR3_X1    g522(.A1(new_n946), .A2(KEYINPUT42), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT42), .B1(new_n946), .B2(new_n947), .ZN(new_n949));
  XOR2_X1   g524(.A(G303), .B(G305), .Z(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n810), .ZN(new_n951));
  OR2_X1    g526(.A1(G166), .A2(G305), .ZN(new_n952));
  NAND2_X1  g527(.A1(G166), .A2(G305), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(G290), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n951), .A2(new_n831), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n831), .B1(new_n951), .B2(new_n954), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n948), .A2(new_n949), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n958), .B1(new_n948), .B2(new_n949), .ZN(new_n960));
  OAI21_X1  g535(.A(G868), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n892), .A2(new_n635), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(G295));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n962), .ZN(G331));
  INV_X1    g539(.A(KEYINPUT101), .ZN(new_n965));
  NAND3_X1  g540(.A1(G168), .A2(new_n965), .A3(G171), .ZN(new_n966));
  NAND2_X1  g541(.A1(G301), .A2(KEYINPUT101), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n554), .A2(new_n965), .A3(new_n555), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(G286), .A3(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n902), .A2(new_n966), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n966), .A2(new_n969), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n971), .A2(new_n900), .A3(new_n901), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n970), .A2(new_n940), .A3(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT102), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n970), .A2(new_n972), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n973), .A2(new_n974), .B1(new_n975), .B2(new_n944), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n970), .A2(KEYINPUT102), .A3(new_n940), .A4(new_n972), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT103), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n978), .B1(new_n956), .B2(new_n957), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n951), .A2(new_n954), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n830), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n981), .A2(KEYINPUT103), .A3(new_n955), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n976), .A2(new_n977), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT104), .B1(new_n983), .B2(G37), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n979), .A2(new_n982), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n973), .A2(new_n974), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n975), .A2(new_n944), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n986), .A2(new_n977), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT104), .ZN(new_n990));
  INV_X1    g565(.A(G37), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n976), .A2(new_n958), .A3(new_n977), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n984), .A2(new_n992), .A3(KEYINPUT43), .A4(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT43), .ZN(new_n996));
  INV_X1    g571(.A(new_n973), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n975), .A2(new_n944), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT105), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n987), .A2(KEYINPUT105), .ZN(new_n1001));
  AOI22_X1  g576(.A1(new_n1000), .A2(new_n1001), .B1(new_n982), .B2(new_n979), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n993), .A2(new_n991), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n996), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n994), .A2(new_n995), .A3(new_n1004), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n1002), .A2(new_n1003), .A3(new_n996), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n984), .A2(new_n993), .A3(new_n992), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1006), .B1(new_n996), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1005), .B1(new_n1008), .B2(new_n995), .ZN(G397));
  AND2_X1   g584(.A1(new_n501), .A2(new_n507), .ZN(new_n1010));
  AOI21_X1  g585(.A(G1384), .B1(new_n1010), .B2(new_n498), .ZN(new_n1011));
  NAND4_X1  g586(.A1(G160), .A2(new_n1011), .A3(KEYINPUT121), .A4(G40), .ZN(new_n1012));
  INV_X1    g587(.A(G2067), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT121), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n471), .A2(G40), .A3(new_n478), .A4(new_n481), .ZN(new_n1015));
  INV_X1    g590(.A(G1384), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n508), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1014), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1012), .A2(new_n1013), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1015), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1017), .A2(KEYINPUT50), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n508), .A2(new_n1022), .A3(new_n1016), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1020), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1019), .B(new_n622), .C1(new_n1025), .C2(G1348), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1026), .A2(KEYINPUT60), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n1012), .A2(new_n1013), .A3(new_n1018), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1022), .B1(new_n508), .B2(new_n1016), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(new_n1015), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1348), .B1(new_n1030), .B2(new_n1023), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n895), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1032), .A2(KEYINPUT60), .A3(new_n1026), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1027), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1017), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n508), .A2(KEYINPUT45), .A3(new_n1016), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1036), .A2(G40), .A3(G160), .A4(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g613(.A(KEYINPUT56), .B(G2072), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  OAI22_X1  g615(.A1(new_n1025), .A2(G1956), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT119), .B1(G299), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT119), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n626), .A2(new_n1044), .A3(KEYINPUT57), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n588), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n578), .A2(KEYINPUT116), .ZN(new_n1049));
  OR2_X1    g624(.A1(new_n578), .A2(KEYINPUT116), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n583), .A2(new_n587), .A3(KEYINPUT117), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1052), .A2(KEYINPUT118), .A3(new_n1042), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT118), .B1(new_n1052), .B2(new_n1042), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1041), .B(new_n1046), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT61), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1046), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1041), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1034), .B1(new_n1055), .B2(new_n1059), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1012), .A2(new_n1018), .ZN(new_n1061));
  XNOR2_X1  g636(.A(KEYINPUT58), .B(G1341), .ZN(new_n1062));
  OAI22_X1  g637(.A1(new_n1061), .A2(new_n1062), .B1(G1996), .B2(new_n1038), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n567), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n1064), .B(KEYINPUT59), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1057), .A2(new_n1066), .A3(new_n1058), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1066), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1055), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1060), .B(new_n1065), .C1(new_n1070), .C2(KEYINPUT61), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n622), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1055), .A2(new_n1072), .ZN(new_n1073));
  OR3_X1    g648(.A1(new_n1073), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT45), .B1(new_n508), .B2(new_n1016), .ZN(new_n1076));
  INV_X1    g651(.A(G40), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1076), .A2(new_n758), .A3(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1037), .B1(new_n1078), .B2(KEYINPUT112), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1077), .B1(new_n1017), .B2(new_n1035), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1080), .A2(KEYINPUT112), .A3(G160), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n705), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1083));
  XNOR2_X1  g658(.A(KEYINPUT113), .B(G2084), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1025), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT114), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1025), .A2(KEYINPUT114), .A3(new_n1084), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1083), .A2(new_n1087), .A3(G168), .A4(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(G8), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G1961), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1024), .A2(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n1094), .B(KEYINPUT123), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1080), .A2(new_n793), .A3(G160), .A4(new_n1037), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n471), .A2(new_n481), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT124), .ZN(new_n1100));
  AND4_X1   g675(.A1(new_n478), .A2(new_n1080), .A3(new_n1037), .A4(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1097), .A2(G2078), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1101), .B(new_n1102), .C1(KEYINPUT124), .C2(new_n1099), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1095), .A2(new_n1098), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(G171), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1036), .A2(G40), .A3(G160), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT112), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1108), .A2(new_n1102), .A3(new_n1081), .A4(new_n1037), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1096), .A2(new_n1097), .B1(new_n1024), .B2(new_n1093), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1105), .B(KEYINPUT54), .C1(G171), .C2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1083), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(G286), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1114), .A2(KEYINPUT51), .A3(G8), .A4(new_n1089), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT111), .ZN(new_n1116));
  AOI21_X1  g691(.A(G1971), .B1(new_n1078), .B2(new_n1037), .ZN(new_n1117));
  INV_X1    g692(.A(G2090), .ZN(new_n1118));
  AND4_X1   g693(.A1(new_n1118), .A2(new_n1020), .A3(new_n1021), .A4(new_n1023), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1116), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1038), .A2(new_n840), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1030), .A2(new_n1118), .A3(new_n1023), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1121), .A2(KEYINPUT111), .A3(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1120), .A2(G8), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(G303), .A2(G8), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT55), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT109), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT109), .ZN(new_n1129));
  AOI211_X1 g704(.A(new_n1129), .B(KEYINPUT55), .C1(G303), .C2(G8), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT108), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g709(.A1(G303), .A2(KEYINPUT108), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1128), .A2(new_n1131), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1124), .A2(new_n1136), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1135), .ZN(new_n1139));
  OAI22_X1  g714(.A1(new_n1138), .A2(new_n1139), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT107), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT107), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1121), .A2(new_n1142), .A3(new_n1122), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1140), .A2(new_n1141), .A3(G8), .A4(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(G305), .A2(G1981), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n602), .B(new_n596), .ZN(new_n1146));
  INV_X1    g721(.A(G1981), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1146), .A2(new_n1147), .A3(new_n595), .A4(new_n601), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT49), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(G8), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1145), .A2(new_n1148), .A3(KEYINPUT49), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1151), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(G1976), .ZN(new_n1156));
  AOI21_X1  g731(.A(KEYINPUT52), .B1(G288), .B2(new_n1156), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1153), .B(new_n1157), .C1(new_n831), .C2(new_n1156), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1156), .B1(new_n827), .B2(new_n829), .ZN(new_n1159));
  OAI21_X1  g734(.A(KEYINPUT52), .B1(new_n1159), .B2(new_n1152), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1155), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1137), .A2(new_n1144), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1162), .ZN(new_n1163));
  AND4_X1   g738(.A1(new_n1092), .A2(new_n1112), .A3(new_n1115), .A4(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1111), .A2(G171), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1095), .A2(G301), .A3(new_n1098), .A4(new_n1103), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1111), .A2(KEYINPUT122), .A3(G171), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT54), .ZN(new_n1172));
  AND3_X1   g747(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1171), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1075), .A2(new_n1164), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT63), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1113), .A2(G8), .A3(G168), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1177), .B1(new_n1162), .B2(new_n1178), .ZN(new_n1179));
  AND3_X1   g754(.A1(new_n1113), .A2(G8), .A3(G168), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1141), .A2(new_n1143), .A3(G8), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1177), .B1(new_n1181), .B2(new_n1136), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1180), .A2(new_n1182), .A3(new_n1144), .A4(new_n1161), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1179), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1181), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1185), .A2(new_n1161), .A3(new_n1140), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1148), .B1(new_n1187), .B2(G288), .ZN(new_n1188));
  OR2_X1    g763(.A1(new_n1188), .A2(KEYINPUT110), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(KEYINPUT110), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1189), .A2(new_n1153), .A3(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1184), .A2(new_n1186), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT115), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT62), .ZN(new_n1196));
  AND3_X1   g771(.A1(new_n1115), .A2(new_n1196), .A3(new_n1092), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1196), .B1(new_n1115), .B2(new_n1092), .ZN(new_n1198));
  OAI211_X1 g773(.A(new_n1195), .B(new_n1163), .C1(new_n1197), .C2(new_n1198), .ZN(new_n1199));
  NAND4_X1  g774(.A1(new_n1184), .A2(KEYINPUT115), .A3(new_n1186), .A4(new_n1191), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1176), .A2(new_n1194), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(G1996), .ZN(new_n1202));
  OR2_X1    g777(.A1(new_n908), .A2(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n906), .B(G2067), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n908), .A2(new_n1202), .ZN(new_n1205));
  AND3_X1   g780(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n819), .A2(new_n823), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n818), .A2(new_n822), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1209), .B1(G1986), .B2(G290), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1210), .B1(G1986), .B2(G290), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1020), .A2(new_n1076), .ZN(new_n1212));
  XOR2_X1   g787(.A(new_n1212), .B(KEYINPUT106), .Z(new_n1213));
  NAND2_X1  g788(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1201), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(new_n1213), .ZN(new_n1216));
  XOR2_X1   g791(.A(new_n1207), .B(KEYINPUT126), .Z(new_n1217));
  NAND2_X1  g792(.A1(new_n1206), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n906), .A2(new_n1013), .ZN(new_n1219));
  AOI21_X1  g794(.A(new_n1216), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g795(.A(KEYINPUT46), .ZN(new_n1221));
  OAI22_X1  g796(.A1(new_n1216), .A2(G1996), .B1(KEYINPUT127), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1204), .A2(new_n908), .ZN(new_n1223));
  AOI22_X1  g798(.A1(new_n1213), .A2(new_n1223), .B1(KEYINPUT127), .B2(new_n1221), .ZN(new_n1224));
  NOR2_X1   g799(.A1(new_n1221), .A2(KEYINPUT127), .ZN(new_n1225));
  NAND3_X1  g800(.A1(new_n1213), .A2(new_n1202), .A3(new_n1225), .ZN(new_n1226));
  NAND3_X1  g801(.A1(new_n1222), .A2(new_n1224), .A3(new_n1226), .ZN(new_n1227));
  XOR2_X1   g802(.A(new_n1227), .B(KEYINPUT47), .Z(new_n1228));
  NAND2_X1  g803(.A1(new_n1209), .A2(new_n1213), .ZN(new_n1229));
  NAND3_X1  g804(.A1(new_n1213), .A2(new_n812), .A3(new_n810), .ZN(new_n1230));
  XNOR2_X1  g805(.A(new_n1230), .B(KEYINPUT48), .ZN(new_n1231));
  AOI211_X1 g806(.A(new_n1220), .B(new_n1228), .C1(new_n1229), .C2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1215), .A2(new_n1232), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g808(.A(new_n460), .B1(new_n928), .B2(new_n930), .ZN(new_n1235));
  INV_X1    g809(.A(new_n1235), .ZN(new_n1236));
  NOR2_X1   g810(.A1(G229), .A2(G227), .ZN(new_n1237));
  NAND4_X1  g811(.A1(new_n994), .A2(new_n666), .A3(new_n1004), .A4(new_n1237), .ZN(new_n1238));
  NOR2_X1   g812(.A1(new_n1236), .A2(new_n1238), .ZN(G308));
  AND2_X1   g813(.A1(new_n994), .A2(new_n1004), .ZN(new_n1240));
  NAND4_X1  g814(.A1(new_n1240), .A2(new_n666), .A3(new_n1235), .A4(new_n1237), .ZN(G225));
endmodule


