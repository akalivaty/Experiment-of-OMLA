//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 1 1 0 1 0 0 0 0 1 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n600, new_n601,
    new_n602, new_n603, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964;
  XNOR2_X1  g000(.A(KEYINPUT69), .B(G119), .ZN(new_n187));
  INV_X1    g001(.A(G128), .ZN(new_n188));
  AOI21_X1  g002(.A(KEYINPUT23), .B1(new_n187), .B2(new_n188), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(G119), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n190), .B1(new_n187), .B2(new_n188), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n189), .B1(KEYINPUT23), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G110), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT24), .B(G110), .Z(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  AOI22_X1  g009(.A1(new_n192), .A2(new_n193), .B1(new_n191), .B2(new_n195), .ZN(new_n196));
  XOR2_X1   g010(.A(new_n196), .B(KEYINPUT78), .Z(new_n197));
  XOR2_X1   g011(.A(G125), .B(G140), .Z(new_n198));
  INV_X1    g012(.A(KEYINPUT16), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G125), .ZN(new_n200));
  OAI22_X1  g014(.A1(new_n198), .A2(new_n199), .B1(G140), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  OR2_X1    g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  OR2_X1    g017(.A1(new_n198), .A2(G146), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n197), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(new_n201), .B(new_n202), .ZN(new_n206));
  OAI221_X1 g020(.A(new_n206), .B1(new_n193), .B2(new_n192), .C1(new_n191), .C2(new_n195), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT22), .B(G137), .ZN(new_n208));
  INV_X1    g022(.A(G953), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(G221), .A3(G234), .ZN(new_n210));
  XNOR2_X1  g024(.A(new_n208), .B(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n205), .A2(new_n207), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n205), .A2(new_n207), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n213), .B(KEYINPUT79), .ZN(new_n214));
  XOR2_X1   g028(.A(new_n211), .B(KEYINPUT80), .Z(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT25), .B1(new_n217), .B2(G902), .ZN(new_n218));
  INV_X1    g032(.A(G217), .ZN(new_n219));
  INV_X1    g033(.A(G902), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n219), .B1(G234), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT79), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n213), .B(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n215), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT25), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n224), .A2(new_n225), .A3(new_n220), .A4(new_n212), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n218), .A2(new_n221), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n217), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n221), .A2(G902), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT81), .B(G104), .ZN(new_n233));
  INV_X1    g047(.A(G107), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT3), .ZN(new_n236));
  OR2_X1    g050(.A1(new_n233), .A2(new_n234), .ZN(new_n237));
  INV_X1    g051(.A(G104), .ZN(new_n238));
  OR3_X1    g052(.A1(new_n238), .A2(KEYINPUT3), .A3(G107), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n236), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G101), .ZN(new_n241));
  INV_X1    g055(.A(G101), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n236), .A2(new_n237), .A3(new_n242), .A4(new_n239), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n241), .A2(KEYINPUT4), .A3(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n202), .A2(G143), .ZN(new_n245));
  AND2_X1   g059(.A1(KEYINPUT64), .A2(G143), .ZN(new_n246));
  NOR2_X1   g060(.A1(KEYINPUT64), .A2(G143), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n245), .B1(new_n248), .B2(new_n202), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT0), .B(G128), .ZN(new_n250));
  OAI21_X1  g064(.A(KEYINPUT65), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G143), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(G146), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT64), .B(G143), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n253), .B1(new_n254), .B2(G146), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(KEYINPUT0), .A3(G128), .ZN(new_n256));
  INV_X1    g070(.A(new_n250), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT65), .ZN(new_n258));
  NOR3_X1   g072(.A1(new_n246), .A2(new_n247), .A3(G146), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n257), .B(new_n258), .C1(new_n259), .C2(new_n245), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n251), .A2(new_n256), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n240), .A2(new_n263), .A3(G101), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n244), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT82), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n266), .B1(new_n238), .B2(G107), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n235), .A2(new_n267), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n268), .B(G101), .C1(KEYINPUT82), .C2(new_n235), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n243), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT1), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n255), .A2(new_n272), .A3(G128), .ZN(new_n273));
  OAI21_X1  g087(.A(G128), .B1(new_n253), .B2(new_n272), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n274), .B1(new_n259), .B2(new_n245), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n271), .A2(KEYINPUT10), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT11), .ZN(new_n278));
  INV_X1    g092(.A(G134), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n278), .B1(new_n279), .B2(G137), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(G137), .ZN(new_n281));
  INV_X1    g095(.A(G137), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(KEYINPUT11), .A3(G134), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n280), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n284), .B(G131), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n248), .A2(new_n202), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n188), .B1(new_n287), .B2(KEYINPUT1), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n273), .B1(new_n288), .B2(new_n255), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(new_n243), .A3(new_n269), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT10), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n265), .A2(new_n277), .A3(new_n286), .A4(new_n292), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n273), .A2(new_n275), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n270), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n290), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT12), .B1(new_n296), .B2(new_n285), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT12), .ZN(new_n298));
  AOI211_X1 g112(.A(new_n298), .B(new_n286), .C1(new_n295), .C2(new_n290), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n293), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(G110), .B(G140), .ZN(new_n301));
  AND2_X1   g115(.A1(new_n209), .A2(G227), .ZN(new_n302));
  XOR2_X1   g116(.A(new_n301), .B(new_n302), .Z(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n265), .A2(new_n277), .A3(new_n292), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n285), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(new_n293), .A3(new_n303), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n305), .A2(KEYINPUT83), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT83), .B1(new_n305), .B2(new_n308), .ZN(new_n311));
  OAI21_X1  g125(.A(G469), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G469), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n313), .A2(new_n220), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  OR2_X1    g129(.A1(new_n297), .A2(new_n299), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n316), .A2(new_n293), .A3(new_n303), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n303), .B1(new_n307), .B2(new_n293), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n313), .B(new_n220), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n312), .A2(new_n315), .A3(new_n319), .ZN(new_n320));
  XOR2_X1   g134(.A(KEYINPUT9), .B(G234), .Z(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(G221), .B1(new_n322), .B2(G902), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT84), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n320), .A2(KEYINPUT84), .A3(new_n323), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n261), .A2(G125), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n329), .B1(G125), .B2(new_n276), .ZN(new_n330));
  INV_X1    g144(.A(G224), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(G953), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n330), .B(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n333), .B1(KEYINPUT7), .B2(new_n332), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT7), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n330), .B(new_n335), .C1(new_n331), .C2(G953), .ZN(new_n336));
  INV_X1    g150(.A(G116), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G119), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  XOR2_X1   g153(.A(KEYINPUT69), .B(G119), .Z(new_n340));
  AOI21_X1  g154(.A(new_n339), .B1(new_n340), .B2(G116), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT68), .ZN(new_n342));
  OR3_X1    g156(.A1(new_n342), .A2(KEYINPUT2), .A3(G113), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n342), .B1(KEYINPUT2), .B2(G113), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n343), .A2(new_n344), .B1(KEYINPUT2), .B2(G113), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n341), .A2(new_n345), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT70), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT70), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n341), .A2(new_n345), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n346), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(new_n264), .A3(new_n244), .ZN(new_n353));
  XOR2_X1   g167(.A(KEYINPUT85), .B(KEYINPUT5), .Z(new_n354));
  NAND3_X1  g168(.A1(new_n340), .A2(new_n354), .A3(G116), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n355), .A2(G113), .ZN(new_n356));
  INV_X1    g170(.A(new_n341), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n356), .B1(new_n357), .B2(new_n354), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT86), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n348), .A2(new_n350), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT86), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n356), .B(new_n361), .C1(new_n357), .C2(new_n354), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n359), .A2(new_n360), .A3(new_n271), .A4(new_n362), .ZN(new_n363));
  XOR2_X1   g177(.A(G110), .B(G122), .Z(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n353), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT5), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n356), .B1(new_n367), .B2(new_n357), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n360), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n271), .ZN(new_n370));
  XOR2_X1   g184(.A(new_n364), .B(KEYINPUT8), .Z(new_n371));
  NAND3_X1  g185(.A1(new_n359), .A2(new_n360), .A3(new_n362), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n370), .B(new_n371), .C1(new_n372), .C2(new_n271), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n334), .A2(new_n336), .A3(new_n366), .A4(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n353), .A2(new_n363), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n364), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(KEYINPUT6), .A3(new_n366), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT6), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n375), .A2(new_n378), .A3(new_n364), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(new_n333), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n374), .A2(new_n380), .A3(new_n220), .ZN(new_n381));
  OAI21_X1  g195(.A(G210), .B1(G237), .B2(G902), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n381), .A2(KEYINPUT87), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(KEYINPUT87), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n374), .A2(new_n380), .A3(new_n220), .A4(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(G234), .A2(G237), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(G952), .A3(new_n209), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  XOR2_X1   g205(.A(KEYINPUT21), .B(G898), .Z(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n389), .A2(G902), .A3(G953), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n391), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(G214), .B1(G237), .B2(G902), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n388), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G237), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT72), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT72), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G237), .ZN(new_n403));
  AOI21_X1  g217(.A(G953), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G214), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n248), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n406), .B1(G143), .B2(new_n405), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(KEYINPUT17), .A3(G131), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n206), .A2(KEYINPUT91), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT91), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n201), .A2(new_n202), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n203), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n409), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT92), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT92), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n409), .A2(new_n410), .A3(new_n413), .A4(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G131), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n407), .B(new_n418), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n415), .B(new_n417), .C1(KEYINPUT17), .C2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n408), .A2(KEYINPUT18), .A3(G131), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT18), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n407), .B1(new_n422), .B2(new_n418), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n198), .B(KEYINPUT88), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G146), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n204), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n421), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(G113), .B(G122), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT90), .B(G104), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n428), .B(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n420), .A2(new_n427), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n431), .B1(new_n420), .B2(new_n427), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n220), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G475), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n419), .A2(new_n203), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT89), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n438), .B1(new_n198), .B2(KEYINPUT19), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n198), .A2(KEYINPUT19), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n440), .B1(new_n424), .B2(KEYINPUT19), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n439), .B1(new_n441), .B2(new_n438), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(G146), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n427), .B1(new_n437), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n430), .ZN(new_n445));
  AOI21_X1  g259(.A(G475), .B1(new_n432), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n447), .A3(new_n220), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n447), .B1(new_n446), .B2(new_n220), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n436), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G478), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(KEYINPUT15), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n248), .A2(new_n188), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n252), .A2(G128), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n454), .A2(G134), .A3(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(G116), .B(G122), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(G107), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT13), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  OR3_X1    g274(.A1(new_n454), .A2(KEYINPUT93), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n454), .A2(KEYINPUT13), .ZN(new_n462));
  OAI21_X1  g276(.A(KEYINPUT93), .B1(new_n454), .B2(new_n460), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AOI211_X1 g278(.A(new_n456), .B(new_n458), .C1(new_n464), .C2(G134), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n457), .A2(new_n234), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n337), .A2(KEYINPUT14), .A3(G122), .ZN(new_n467));
  INV_X1    g281(.A(new_n457), .ZN(new_n468));
  OAI211_X1 g282(.A(G107), .B(new_n467), .C1(new_n468), .C2(KEYINPUT14), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n454), .A2(new_n455), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(new_n279), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n466), .B(new_n469), .C1(new_n471), .C2(new_n456), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n322), .A2(new_n219), .A3(G953), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n465), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n475), .B1(new_n465), .B2(new_n473), .ZN(new_n478));
  AOI21_X1  g292(.A(G902), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n479), .A2(KEYINPUT94), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n479), .A2(KEYINPUT94), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n453), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OR2_X1    g296(.A1(new_n481), .A2(new_n453), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n451), .A2(new_n484), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n328), .A2(new_n399), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT77), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n261), .A2(KEYINPUT66), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT66), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n251), .A2(new_n489), .A3(new_n256), .A4(new_n260), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n488), .A2(new_n285), .A3(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT30), .ZN(new_n492));
  OR2_X1    g306(.A1(new_n284), .A2(G131), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT67), .ZN(new_n494));
  INV_X1    g308(.A(new_n281), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n279), .A2(G137), .ZN(new_n496));
  OAI21_X1  g310(.A(G131), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n493), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n494), .B1(new_n493), .B2(new_n497), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n276), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n491), .A2(new_n492), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n276), .A2(new_n493), .A3(new_n497), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n285), .A2(new_n251), .A3(new_n256), .A4(new_n260), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT30), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n352), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT71), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n404), .A2(G210), .ZN(new_n509));
  XOR2_X1   g323(.A(KEYINPUT73), .B(KEYINPUT27), .Z(new_n510));
  XNOR2_X1  g324(.A(new_n509), .B(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT26), .B(G101), .ZN(new_n512));
  XOR2_X1   g326(.A(new_n511), .B(new_n512), .Z(new_n513));
  NAND3_X1  g327(.A1(new_n351), .A2(new_n502), .A3(new_n503), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT71), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n506), .A2(new_n515), .A3(new_n352), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n508), .A2(new_n513), .A3(new_n514), .A4(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT31), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n515), .B1(new_n506), .B2(new_n352), .ZN(new_n519));
  AOI211_X1 g333(.A(KEYINPUT71), .B(new_n351), .C1(new_n501), .C2(new_n505), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT31), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n521), .A2(new_n522), .A3(new_n513), .A4(new_n514), .ZN(new_n523));
  INV_X1    g337(.A(new_n514), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(KEYINPUT28), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT28), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n514), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n351), .B1(new_n491), .B2(new_n500), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n525), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT74), .B1(new_n529), .B2(new_n513), .ZN(new_n530));
  INV_X1    g344(.A(new_n525), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n528), .A2(new_n527), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT74), .ZN(new_n534));
  INV_X1    g348(.A(new_n513), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n530), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n518), .A2(new_n523), .A3(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(G472), .A2(G902), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT32), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT75), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n538), .A2(KEYINPUT32), .A3(new_n539), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n540), .A2(KEYINPUT75), .A3(new_n541), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n521), .A2(new_n514), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT29), .B1(new_n548), .B2(new_n535), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n535), .B2(new_n533), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT76), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n352), .A2(new_n504), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n514), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT28), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n551), .B1(new_n531), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n555), .B1(new_n551), .B2(new_n554), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n513), .A2(KEYINPUT29), .ZN(new_n557));
  AOI21_X1  g371(.A(G902), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n550), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(G472), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n487), .B1(new_n547), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(G472), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n562), .B1(new_n550), .B2(new_n558), .ZN(new_n563));
  AOI211_X1 g377(.A(KEYINPUT77), .B(new_n563), .C1(new_n545), .C2(new_n546), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n232), .B(new_n486), .C1(new_n561), .C2(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(G101), .ZN(G3));
  NAND2_X1  g380(.A1(new_n538), .A2(new_n220), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G472), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n568), .A2(new_n540), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n328), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n232), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n381), .B(new_n383), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n397), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT95), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT95), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n573), .A2(new_n576), .A3(new_n397), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(new_n396), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n446), .A2(new_n220), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT20), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n581), .A2(new_n448), .B1(G475), .B2(new_n435), .ZN(new_n582));
  OAI21_X1  g396(.A(KEYINPUT33), .B1(new_n474), .B2(KEYINPUT96), .ZN(new_n583));
  INV_X1    g397(.A(new_n465), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n474), .B1(new_n584), .B2(new_n472), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n583), .B1(new_n585), .B2(new_n476), .ZN(new_n586));
  INV_X1    g400(.A(new_n583), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n477), .A2(new_n478), .A3(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n586), .A2(new_n588), .A3(G478), .A4(new_n220), .ZN(new_n589));
  OR2_X1    g403(.A1(new_n589), .A2(KEYINPUT97), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(KEYINPUT97), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT98), .B1(new_n479), .B2(G478), .ZN(new_n592));
  OR3_X1    g406(.A1(new_n479), .A2(KEYINPUT98), .A3(G478), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n590), .A2(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n582), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n579), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n572), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT34), .B(G104), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(G6));
  AND2_X1   g413(.A1(new_n582), .A2(new_n484), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n579), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n572), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT35), .B(G107), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G9));
  NOR2_X1   g418(.A1(new_n215), .A2(KEYINPUT36), .ZN(new_n605));
  XOR2_X1   g419(.A(new_n605), .B(KEYINPUT99), .Z(new_n606));
  XNOR2_X1  g420(.A(new_n223), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n229), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT100), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT100), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n607), .A2(new_n610), .A3(new_n229), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n227), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n486), .A2(new_n569), .A3(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT37), .B(G110), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G12));
  AND3_X1   g429(.A1(new_n609), .A2(new_n227), .A3(new_n611), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n544), .A2(new_n543), .ZN(new_n617));
  AOI21_X1  g431(.A(KEYINPUT32), .B1(new_n538), .B2(new_n539), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n546), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n560), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(KEYINPUT77), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n547), .A2(new_n487), .A3(new_n560), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n616), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n390), .B(KEYINPUT101), .ZN(new_n625));
  INV_X1    g439(.A(G900), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n625), .B1(new_n626), .B2(new_n395), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n600), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n578), .B1(new_n326), .B2(new_n327), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n624), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G128), .ZN(G30));
  XOR2_X1   g447(.A(KEYINPUT102), .B(KEYINPUT39), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n627), .B(new_n634), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n320), .A2(KEYINPUT84), .A3(new_n323), .ZN(new_n636));
  AOI21_X1  g450(.A(KEYINPUT84), .B1(new_n320), .B2(new_n323), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT40), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n328), .A2(KEYINPUT40), .A3(new_n635), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n387), .B(KEYINPUT38), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n451), .A2(new_n484), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n548), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(new_n535), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n220), .B1(new_n553), .B2(new_n513), .ZN(new_n649));
  OAI21_X1  g463(.A(G472), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n547), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n612), .A2(new_n398), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n642), .A2(new_n646), .A3(new_n651), .A4(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT103), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(new_n254), .ZN(G45));
  NOR3_X1   g470(.A1(new_n582), .A2(new_n594), .A3(new_n627), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n624), .A2(new_n631), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G146), .ZN(G48));
  OR2_X1    g473(.A1(new_n317), .A2(new_n318), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n220), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(G469), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n662), .A2(new_n323), .A3(new_n319), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n232), .B(new_n664), .C1(new_n561), .C2(new_n564), .ZN(new_n665));
  OR2_X1    g479(.A1(new_n665), .A2(new_n596), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT41), .B(G113), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT104), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n666), .B(new_n668), .ZN(G15));
  OR2_X1    g483(.A1(new_n665), .A2(new_n601), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G116), .ZN(G18));
  OAI211_X1 g485(.A(new_n579), .B(new_n612), .C1(new_n561), .C2(new_n564), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n664), .A2(new_n485), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(new_n674), .B(G119), .Z(G21));
  OR2_X1    g489(.A1(new_n568), .A2(KEYINPUT106), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n568), .A2(KEYINPUT106), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n518), .A2(new_n523), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n556), .A2(new_n513), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n539), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OR2_X1    g496(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  AOI22_X1  g497(.A1(new_n676), .A2(new_n677), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n645), .A2(new_n663), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n579), .A2(new_n684), .A3(new_n232), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G122), .ZN(G24));
  NAND2_X1  g501(.A1(new_n684), .A2(new_n612), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n578), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n689), .A2(new_n690), .A3(new_n657), .A4(new_n664), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G125), .ZN(G27));
  NAND2_X1  g506(.A1(new_n622), .A2(new_n623), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n387), .A2(new_n398), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n314), .B(KEYINPUT107), .Z(new_n696));
  NAND2_X1  g510(.A1(new_n305), .A2(new_n308), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n319), .B(new_n696), .C1(new_n313), .C2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n323), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n693), .A2(new_n232), .A3(new_n657), .A4(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT42), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n542), .A2(KEYINPUT108), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n560), .A3(new_n544), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n542), .A2(KEYINPUT108), .ZN(new_n706));
  OAI211_X1 g520(.A(KEYINPUT42), .B(new_n232), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n700), .A2(new_n657), .ZN(new_n708));
  OR3_X1    g522(.A1(new_n707), .A2(KEYINPUT109), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g523(.A(KEYINPUT109), .B1(new_n707), .B2(new_n708), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n703), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT110), .B(G131), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G33));
  AND4_X1   g528(.A1(new_n693), .A2(new_n232), .A3(new_n630), .A4(new_n700), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(new_n279), .ZN(G36));
  NAND2_X1  g530(.A1(new_n568), .A2(new_n540), .ZN(new_n717));
  OAI21_X1  g531(.A(KEYINPUT43), .B1(new_n451), .B2(new_n594), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n590), .A2(new_n591), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n593), .A2(new_n592), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n582), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n612), .A2(new_n717), .A3(new_n718), .A4(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT44), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  INV_X1    g541(.A(new_n323), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT83), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n697), .A2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n730), .A2(new_n731), .A3(new_n309), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n305), .A2(KEYINPUT45), .A3(new_n308), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(G469), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT46), .B1(new_n734), .B2(new_n696), .ZN(new_n735));
  INV_X1    g549(.A(new_n319), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n734), .A2(KEYINPUT46), .A3(new_n696), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n728), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n739), .A2(new_n635), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n726), .A2(new_n694), .A3(new_n727), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G137), .ZN(G39));
  NOR2_X1   g556(.A1(new_n561), .A2(new_n564), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n739), .A2(KEYINPUT47), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT47), .ZN(new_n745));
  INV_X1    g559(.A(new_n738), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n746), .A2(new_n735), .A3(new_n736), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n745), .B1(new_n747), .B2(new_n728), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n657), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n232), .A2(new_n750), .A3(new_n695), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n743), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT111), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT111), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n743), .A2(new_n749), .A3(new_n754), .A4(new_n751), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G140), .ZN(G42));
  NOR2_X1   g571(.A1(G952), .A2(G953), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n759));
  NOR2_X1   g573(.A1(KEYINPUT115), .A2(KEYINPUT50), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n718), .A2(new_n723), .A3(new_n625), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n684), .A2(new_n763), .A3(new_n232), .A4(new_n664), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n397), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n761), .B1(new_n765), .B2(new_n644), .ZN(new_n766));
  NOR4_X1   g580(.A1(new_n764), .A2(new_n397), .A3(new_n643), .A4(new_n760), .ZN(new_n767));
  OAI21_X1  g581(.A(KEYINPUT116), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n676), .A2(new_n677), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n683), .A2(new_n682), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(new_n770), .A3(new_n232), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(new_n762), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n772), .A2(new_n398), .A3(new_n644), .A4(new_n664), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n760), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n765), .A2(new_n644), .A3(new_n761), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT116), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n768), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n651), .A2(new_n231), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n695), .A2(new_n663), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n779), .A2(new_n391), .A3(new_n582), .A4(new_n780), .ZN(new_n781));
  OR3_X1    g595(.A1(new_n781), .A2(KEYINPUT117), .A3(new_n721), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n762), .A2(new_n663), .A3(new_n695), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n689), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(KEYINPUT117), .B1(new_n781), .B2(new_n721), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n662), .A2(new_n319), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n323), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n772), .B(new_n694), .C1(new_n749), .C2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n782), .A2(new_n784), .A3(new_n785), .A4(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n759), .B1(new_n778), .B2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI211_X1 g606(.A(KEYINPUT118), .B(new_n759), .C1(new_n778), .C2(new_n789), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n705), .A2(new_n706), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(new_n231), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n783), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT48), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n779), .A2(new_n391), .A3(new_n780), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n595), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n797), .A2(G952), .A3(new_n209), .A4(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n789), .A2(new_n759), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n774), .A2(new_n775), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n792), .A2(new_n793), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n805));
  OAI22_X1  g619(.A1(new_n601), .A2(new_n665), .B1(new_n672), .B2(new_n673), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n686), .B1(new_n665), .B2(new_n596), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n571), .A2(new_n232), .A3(new_n399), .A4(new_n595), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n565), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT112), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT112), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n565), .A2(new_n812), .A3(new_n809), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n399), .A2(new_n600), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT113), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n613), .B1(new_n816), .B2(new_n572), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n808), .A2(new_n814), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n485), .A2(new_n694), .A3(new_n628), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT114), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n820), .A2(new_n821), .B1(new_n326), .B2(new_n327), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n822), .B(new_n823), .C1(new_n561), .C2(new_n564), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n684), .A2(new_n657), .A3(new_n700), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n616), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n826), .A2(new_n715), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n712), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n819), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n624), .B(new_n631), .C1(new_n630), .C2(new_n657), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n612), .A2(new_n627), .A3(new_n699), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n578), .A2(new_n645), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(new_n832), .A3(new_n651), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n830), .A2(new_n691), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT52), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n830), .A2(new_n836), .A3(new_n691), .A4(new_n833), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT53), .B1(new_n829), .B2(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n806), .A2(new_n807), .A3(new_n817), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n840), .A2(new_n712), .A3(new_n814), .A4(new_n827), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n835), .A2(new_n837), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n805), .B1(new_n839), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n829), .A2(KEYINPUT53), .A3(new_n838), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n843), .B1(new_n841), .B2(new_n842), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n847), .A3(KEYINPUT54), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n804), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n772), .A2(new_n690), .A3(new_n664), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n758), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NOR4_X1   g665(.A1(new_n451), .A2(new_n594), .A3(new_n398), .A4(new_n728), .ZN(new_n852));
  XOR2_X1   g666(.A(new_n786), .B(KEYINPUT49), .Z(new_n853));
  NAND4_X1  g667(.A1(new_n779), .A2(new_n644), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT119), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n804), .ZN(new_n857));
  INV_X1    g671(.A(new_n848), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT54), .B1(new_n846), .B2(new_n847), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n857), .B(new_n850), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n758), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n862), .A2(new_n863), .A3(new_n854), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n856), .A2(new_n864), .ZN(G75));
  NAND2_X1  g679(.A1(new_n377), .A2(new_n379), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n866), .B(new_n333), .Z(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT55), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  OAI211_X1 g683(.A(G210), .B(G902), .C1(new_n839), .C2(new_n844), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT56), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT120), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n870), .A2(new_n874), .A3(new_n871), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n869), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n209), .A2(G952), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n868), .B1(new_n872), .B2(KEYINPUT120), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(G51));
  XOR2_X1   g693(.A(new_n696), .B(KEYINPUT57), .Z(new_n880));
  NAND3_X1  g694(.A1(new_n845), .A2(new_n848), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n660), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n220), .B1(new_n846), .B2(new_n847), .ZN(new_n883));
  INV_X1    g697(.A(new_n734), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n877), .B1(new_n882), .B2(new_n885), .ZN(G54));
  NAND3_X1  g700(.A1(new_n883), .A2(KEYINPUT58), .A3(G475), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n432), .A2(new_n445), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n887), .A2(new_n889), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n890), .A2(new_n891), .A3(new_n877), .ZN(G60));
  NAND2_X1  g706(.A1(G478), .A2(G902), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT121), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT59), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n845), .A2(new_n848), .A3(new_n895), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n586), .A2(new_n588), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n896), .A2(new_n898), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n899), .A2(new_n900), .A3(new_n877), .ZN(G63));
  NAND2_X1  g715(.A1(G217), .A2(G902), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT122), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT60), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(new_n846), .B2(new_n847), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n607), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n877), .B1(KEYINPUT123), .B2(new_n908), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n907), .B(new_n909), .C1(new_n228), .C2(new_n906), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n908), .A2(KEYINPUT123), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT124), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n910), .B(new_n913), .ZN(G66));
  OAI21_X1  g728(.A(G953), .B1(new_n393), .B2(new_n331), .ZN(new_n915));
  INV_X1    g729(.A(new_n819), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n915), .B1(new_n916), .B2(G953), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n866), .B1(G898), .B2(new_n209), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n917), .B(new_n918), .ZN(G69));
  NAND2_X1  g733(.A1(G227), .A2(G900), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(G953), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT125), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n506), .B(new_n442), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n756), .A2(new_n741), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT62), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n830), .A2(new_n691), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n926), .B1(new_n655), .B2(new_n927), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n653), .B(KEYINPUT103), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n929), .A2(KEYINPUT62), .A3(new_n691), .A4(new_n830), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n925), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n600), .A2(new_n595), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n932), .A2(new_n638), .A3(new_n695), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n693), .A2(new_n232), .A3(new_n933), .ZN(new_n934));
  AOI211_X1 g748(.A(G953), .B(new_n924), .C1(new_n931), .C2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n715), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n795), .A2(new_n740), .A3(new_n832), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n756), .A2(new_n936), .A3(new_n741), .A4(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n712), .A2(new_n691), .A3(new_n830), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n209), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n626), .A2(G953), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n942), .A2(new_n923), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n922), .B1(new_n935), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT126), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI211_X1 g760(.A(G953), .B(new_n920), .C1(new_n942), .C2(new_n923), .ZN(new_n947));
  OAI211_X1 g761(.A(KEYINPUT126), .B(new_n922), .C1(new_n935), .C2(new_n943), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(KEYINPUT127), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT127), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n946), .A2(new_n951), .A3(new_n947), .A4(new_n948), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n950), .A2(new_n952), .ZN(G72));
  INV_X1    g767(.A(new_n648), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n931), .A2(new_n934), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n916), .ZN(new_n956));
  NAND2_X1  g770(.A1(G472), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT63), .Z(new_n958));
  AOI21_X1  g772(.A(new_n954), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n647), .A2(new_n535), .ZN(new_n960));
  OR3_X1    g774(.A1(new_n819), .A2(new_n938), .A3(new_n939), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n960), .B1(new_n961), .B2(new_n958), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n954), .A2(new_n958), .A3(new_n960), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n963), .B1(new_n846), .B2(new_n847), .ZN(new_n964));
  NOR4_X1   g778(.A1(new_n959), .A2(new_n877), .A3(new_n962), .A4(new_n964), .ZN(G57));
endmodule


