//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n573, new_n574, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n595, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1179, new_n1180;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g024(.A1(G218), .A2(G221), .A3(G219), .A4(G220), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT65), .Z(new_n454));
  OR2_X1    g029(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT66), .Z(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  NAND2_X1  g032(.A1(new_n452), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n454), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n462), .A2(KEYINPUT67), .A3(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n466), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(KEYINPUT68), .A3(G137), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n474), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n468), .A2(new_n465), .ZN(new_n479));
  INV_X1    g054(.A(G125), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n462), .A2(G2105), .ZN(new_n482));
  AOI22_X1  g057(.A1(new_n481), .A2(G2105), .B1(G101), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G160));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n466), .A2(G2105), .A3(new_n470), .ZN(new_n488));
  INV_X1    g063(.A(G124), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(G136), .B2(new_n472), .ZN(G162));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G126), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n495), .B1(new_n488), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT69), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(new_n495), .C1(new_n488), .C2(new_n496), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT4), .B1(new_n471), .B2(new_n501), .ZN(new_n502));
  OR4_X1    g077(.A1(KEYINPUT4), .A2(new_n479), .A3(new_n501), .A4(G2105), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n498), .A2(new_n500), .B1(new_n502), .B2(new_n503), .ZN(G164));
  NAND2_X1  g079(.A1(G75), .A2(G543), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G62), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G651), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n510), .A2(KEYINPUT70), .A3(G651), .ZN(new_n514));
  OR2_X1    g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n515), .A2(new_n516), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n522), .B1(new_n519), .B2(new_n520), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n521), .A2(G88), .B1(new_n523), .B2(G50), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n513), .A2(new_n514), .A3(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND2_X1  g101(.A1(new_n515), .A2(new_n516), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n523), .A2(G51), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n519), .A2(new_n520), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n527), .A2(new_n530), .A3(G89), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT7), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n534), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n529), .A2(new_n531), .A3(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(G168));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n539));
  AND2_X1   g114(.A1(KEYINPUT6), .A2(G651), .ZN(new_n540));
  NOR2_X1   g115(.A1(KEYINPUT6), .A2(G651), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n507), .A2(new_n506), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  OAI21_X1  g118(.A(G543), .B1(new_n540), .B2(new_n541), .ZN(new_n544));
  XNOR2_X1  g119(.A(KEYINPUT71), .B(G52), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n542), .A2(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g121(.A(G64), .B1(new_n506), .B2(new_n507), .ZN(new_n547));
  NAND2_X1  g122(.A1(G77), .A2(G543), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n518), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n539), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G64), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n551), .B1(new_n515), .B2(new_n516), .ZN(new_n552));
  INV_X1    g127(.A(new_n548), .ZN(new_n553));
  OAI21_X1  g128(.A(G651), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n527), .A2(new_n530), .A3(G90), .ZN(new_n555));
  INV_X1    g130(.A(new_n545), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(new_n523), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n554), .A2(KEYINPUT72), .A3(new_n555), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n550), .A2(new_n558), .ZN(G171));
  INV_X1    g134(.A(KEYINPUT73), .ZN(new_n560));
  INV_X1    g135(.A(G56), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n561), .B1(new_n515), .B2(new_n516), .ZN(new_n562));
  NAND2_X1  g137(.A1(G68), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n560), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g140(.A(KEYINPUT73), .B(new_n563), .C1(new_n508), .C2(new_n561), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n565), .A2(G651), .A3(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n521), .A2(G81), .B1(new_n523), .B2(G43), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G860), .ZN(G153));
  NAND4_X1  g146(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND4_X1  g149(.A1(G319), .A2(G483), .A3(G661), .A4(new_n574), .ZN(G188));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G65), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n508), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n578), .A2(G651), .B1(new_n521), .B2(G91), .ZN(new_n579));
  INV_X1    g154(.A(G53), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT9), .B1(new_n544), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT9), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n523), .A2(new_n582), .A3(G53), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n579), .A2(new_n584), .ZN(G299));
  INV_X1    g160(.A(G171), .ZN(G301));
  INV_X1    g161(.A(G89), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n536), .B1(new_n542), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n528), .B1(new_n506), .B2(new_n507), .ZN(new_n589));
  INV_X1    g164(.A(G51), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n544), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(KEYINPUT74), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT74), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n529), .A2(new_n593), .A3(new_n531), .A4(new_n536), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G286));
  NAND2_X1  g171(.A1(new_n521), .A2(G87), .ZN(new_n597));
  OAI21_X1  g172(.A(G651), .B1(new_n527), .B2(G74), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n523), .A2(G49), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(G288));
  AOI22_X1  g175(.A1(new_n527), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(new_n518), .ZN(new_n602));
  INV_X1    g177(.A(G86), .ZN(new_n603));
  INV_X1    g178(.A(G48), .ZN(new_n604));
  OAI22_X1  g179(.A1(new_n542), .A2(new_n603), .B1(new_n544), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(G305));
  AND2_X1   g182(.A1(new_n527), .A2(G60), .ZN(new_n608));
  AND2_X1   g183(.A1(G72), .A2(G543), .ZN(new_n609));
  OAI21_X1  g184(.A(G651), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT75), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI211_X1 g187(.A(KEYINPUT75), .B(G651), .C1(new_n608), .C2(new_n609), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n521), .A2(G85), .B1(new_n523), .B2(G47), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(G290));
  NAND3_X1  g190(.A1(new_n521), .A2(KEYINPUT10), .A3(G92), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT10), .ZN(new_n617));
  INV_X1    g192(.A(G92), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n542), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(G79), .A2(G543), .ZN(new_n621));
  INV_X1    g196(.A(G66), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n508), .B2(new_n622), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n623), .A2(G651), .B1(G54), .B2(new_n523), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n626), .B1(G868), .B2(G171), .ZN(G284));
  XOR2_X1   g202(.A(G284), .B(KEYINPUT76), .Z(G321));
  NOR2_X1   g203(.A1(G299), .A2(G868), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(G868), .B2(new_n595), .ZN(G297));
  AOI21_X1  g205(.A(new_n629), .B1(G868), .B2(new_n595), .ZN(G280));
  INV_X1    g206(.A(new_n625), .ZN(new_n632));
  INV_X1    g207(.A(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(G860), .ZN(G148));
  INV_X1    g209(.A(KEYINPUT77), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n632), .A2(new_n633), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(G868), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(G868), .B2(new_n570), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n636), .A2(new_n635), .A3(G868), .ZN(new_n639));
  AND2_X1   g214(.A1(new_n638), .A2(new_n639), .ZN(G323));
  XNOR2_X1  g215(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g216(.A1(new_n472), .A2(G135), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n467), .A2(G111), .ZN(new_n643));
  OAI21_X1  g218(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n644));
  INV_X1    g219(.A(new_n488), .ZN(new_n645));
  AND3_X1   g220(.A1(new_n645), .A2(KEYINPUT78), .A3(G123), .ZN(new_n646));
  AOI21_X1  g221(.A(KEYINPUT78), .B1(new_n645), .B2(G123), .ZN(new_n647));
  OAI221_X1 g222(.A(new_n642), .B1(new_n643), .B2(new_n644), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n648), .A2(G2096), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(G2096), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT12), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT13), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2100), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n649), .A2(new_n650), .A3(new_n654), .ZN(G156));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT80), .B(G2438), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2427), .B(G2430), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(KEYINPUT14), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n662), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2451), .B(G2454), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n666), .A2(new_n669), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(G14), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT81), .Z(G401));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2084), .B(G2090), .Z(new_n676));
  XNOR2_X1  g251(.A(G2067), .B(G2678), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT18), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT84), .B(KEYINPUT17), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n674), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n676), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n682), .A2(new_n677), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n679), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n677), .B1(new_n675), .B2(KEYINPUT82), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(KEYINPUT82), .B2(new_n675), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n686), .A2(KEYINPUT83), .A3(new_n682), .ZN(new_n687));
  INV_X1    g262(.A(new_n677), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n688), .B2(new_n681), .ZN(new_n689));
  AOI21_X1  g264(.A(KEYINPUT83), .B1(new_n686), .B2(new_n682), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n684), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(G2100), .Z(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT85), .B(G2096), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(G227));
  XOR2_X1   g270(.A(G1971), .B(G1976), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT19), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1956), .B(G2474), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(G1961), .B(G1966), .Z(new_n700));
  AND2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT20), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n699), .A2(new_n700), .ZN(new_n704));
  NOR3_X1   g279(.A1(new_n697), .A2(new_n701), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n697), .B2(new_n704), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT86), .Z(new_n708));
  XNOR2_X1  g283(.A(G1991), .B(G1996), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(G1981), .B(G1986), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT87), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n710), .B(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(G229));
  INV_X1    g291(.A(G141), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n471), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT100), .ZN(new_n719));
  NAND3_X1  g294(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT26), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n482), .A2(G105), .ZN(new_n722));
  AOI211_X1 g297(.A(new_n721), .B(new_n722), .C1(new_n645), .C2(G129), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n719), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G29), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n726), .B2(G32), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT27), .B(G1996), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n648), .A2(new_n726), .ZN(new_n731));
  INV_X1    g306(.A(G16), .ZN(new_n732));
  NOR2_X1   g307(.A1(G168), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n732), .B2(G21), .ZN(new_n734));
  INV_X1    g309(.A(G1966), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT30), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n737), .A2(G28), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n726), .B1(new_n737), .B2(G28), .ZN(new_n739));
  AND2_X1   g314(.A1(KEYINPUT31), .A2(G11), .ZN(new_n740));
  NOR2_X1   g315(.A1(KEYINPUT31), .A2(G11), .ZN(new_n741));
  OAI22_X1  g316(.A1(new_n738), .A2(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n734), .B2(new_n735), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n730), .A2(new_n731), .A3(new_n736), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT102), .B(KEYINPUT23), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n732), .A2(G20), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G299), .B2(G16), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1956), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n732), .A2(G5), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G171), .B2(new_n732), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n749), .B1(new_n751), .B2(G1961), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n732), .A2(G19), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n570), .B2(new_n732), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1341), .ZN(new_n755));
  OR3_X1    g330(.A1(new_n744), .A2(new_n752), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n726), .A2(G26), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT96), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT28), .ZN(new_n759));
  INV_X1    g334(.A(G128), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n467), .A2(G116), .ZN(new_n761));
  OAI21_X1  g336(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n762));
  OAI22_X1  g337(.A1(new_n488), .A2(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G140), .B2(new_n472), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n759), .B1(new_n764), .B2(new_n726), .ZN(new_n765));
  INV_X1    g340(.A(G2067), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(G34), .ZN(new_n768));
  AOI21_X1  g343(.A(G29), .B1(new_n768), .B2(KEYINPUT24), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(KEYINPUT24), .B2(new_n768), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n484), .B2(new_n726), .ZN(new_n771));
  INV_X1    g346(.A(G2084), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n767), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n771), .A2(new_n772), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n774), .B(new_n775), .C1(new_n728), .C2(new_n729), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n732), .A2(G4), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n632), .B2(new_n732), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT95), .ZN(new_n779));
  INV_X1    g354(.A(G1348), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n751), .A2(G1961), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT101), .Z(new_n783));
  NOR4_X1   g358(.A1(new_n756), .A2(new_n776), .A3(new_n781), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n726), .A2(G33), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n472), .A2(KEYINPUT97), .A3(G139), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT25), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(KEYINPUT97), .B1(new_n472), .B2(G139), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT98), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n468), .A2(new_n465), .A3(G127), .ZN(new_n793));
  NAND2_X1  g368(.A1(G115), .A2(G2104), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n467), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n785), .B1(new_n796), .B2(new_n726), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT99), .ZN(new_n798));
  INV_X1    g373(.A(G2072), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n726), .A2(G35), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G162), .B2(new_n726), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT29), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G2090), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n726), .A2(G27), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G164), .B2(new_n726), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G2078), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n784), .A2(new_n800), .A3(new_n801), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n732), .A2(G6), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n606), .B2(new_n732), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT93), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT32), .B(G1981), .Z(new_n814));
  NAND2_X1  g389(.A1(G166), .A2(G16), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G16), .B2(G22), .ZN(new_n816));
  INV_X1    g391(.A(G1971), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n813), .A2(new_n814), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n817), .B2(new_n816), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n732), .A2(G23), .ZN(new_n820));
  INV_X1    g395(.A(G288), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(new_n732), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT33), .B(G1976), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n813), .B2(new_n814), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n819), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(KEYINPUT34), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT94), .ZN(new_n828));
  NOR2_X1   g403(.A1(G16), .A2(G24), .ZN(new_n829));
  XOR2_X1   g404(.A(G290), .B(KEYINPUT91), .Z(new_n830));
  AOI21_X1  g405(.A(new_n829), .B1(new_n830), .B2(G16), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT92), .Z(new_n832));
  OR2_X1    g407(.A1(new_n832), .A2(G1986), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n826), .A2(KEYINPUT34), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n726), .A2(G25), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT88), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n472), .A2(G131), .ZN(new_n837));
  OR2_X1    g412(.A1(G95), .A2(G2105), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n838), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT89), .Z(new_n840));
  AOI211_X1 g415(.A(new_n837), .B(new_n840), .C1(G119), .C2(new_n645), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n836), .B1(new_n841), .B2(new_n726), .ZN(new_n842));
  XOR2_X1   g417(.A(KEYINPUT35), .B(G1991), .Z(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT90), .Z(new_n844));
  XNOR2_X1  g419(.A(new_n842), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n832), .A2(G1986), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n833), .A2(new_n834), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  OR3_X1    g422(.A1(new_n828), .A2(new_n847), .A3(KEYINPUT36), .ZN(new_n848));
  OAI21_X1  g423(.A(KEYINPUT36), .B1(new_n828), .B2(new_n847), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n810), .B1(new_n848), .B2(new_n849), .ZN(G311));
  INV_X1    g425(.A(G311), .ZN(G150));
  AOI22_X1  g426(.A1(new_n521), .A2(G93), .B1(new_n523), .B2(G55), .ZN(new_n852));
  INV_X1    g427(.A(G67), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(new_n515), .B2(new_n516), .ZN(new_n854));
  NAND2_X1  g429(.A1(G80), .A2(G543), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(G651), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(KEYINPUT103), .B1(new_n852), .B2(new_n857), .ZN(new_n858));
  OAI211_X1 g433(.A(G55), .B(G543), .C1(new_n540), .C2(new_n541), .ZN(new_n859));
  INV_X1    g434(.A(G93), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n859), .B1(new_n542), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(G67), .B1(new_n506), .B2(new_n507), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n518), .B1(new_n862), .B2(new_n855), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT103), .ZN(new_n864));
  NOR3_X1   g439(.A1(new_n861), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n858), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(KEYINPUT105), .B(G860), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT37), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n569), .B1(new_n858), .B2(new_n865), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n861), .A2(new_n863), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n871), .A2(new_n567), .A3(new_n568), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT38), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n632), .A2(G559), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT104), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n867), .B1(new_n876), .B2(new_n877), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n869), .B1(new_n879), .B2(new_n880), .ZN(G145));
  XNOR2_X1  g456(.A(new_n484), .B(G162), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(new_n648), .Z(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n724), .B(new_n764), .ZN(new_n885));
  OR2_X1    g460(.A1(G106), .A2(G2105), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n886), .B(G2104), .C1(G118), .C2(new_n467), .ZN(new_n887));
  INV_X1    g462(.A(G130), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n887), .B1(new_n488), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n889), .B1(G142), .B2(new_n472), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n885), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n885), .A2(new_n891), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n841), .B(new_n652), .ZN(new_n895));
  NOR3_X1   g470(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n895), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n885), .A2(new_n891), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n897), .B1(new_n898), .B2(new_n892), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n796), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n502), .A2(new_n503), .ZN(new_n901));
  INV_X1    g476(.A(new_n497), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n895), .B1(new_n893), .B2(new_n894), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n898), .A2(new_n897), .A3(new_n892), .ZN(new_n906));
  INV_X1    g481(.A(new_n796), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n900), .A2(new_n904), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n904), .B1(new_n900), .B2(new_n908), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n884), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(G37), .ZN(new_n912));
  INV_X1    g487(.A(new_n908), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n907), .B1(new_n905), .B2(new_n906), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n903), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n900), .A2(new_n904), .A3(new_n908), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(new_n883), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n911), .A2(new_n912), .A3(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n918), .B(new_n919), .ZN(G395));
  XNOR2_X1  g495(.A(G166), .B(G290), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n606), .B(new_n821), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n921), .B(new_n922), .ZN(new_n923));
  XOR2_X1   g498(.A(new_n923), .B(KEYINPUT42), .Z(new_n924));
  XOR2_X1   g499(.A(new_n873), .B(new_n636), .Z(new_n925));
  NOR2_X1   g500(.A1(new_n625), .A2(G299), .ZN(new_n926));
  AOI22_X1  g501(.A1(new_n620), .A2(new_n624), .B1(new_n579), .B2(new_n584), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n930), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n925), .A2(new_n932), .ZN(new_n933));
  OR2_X1    g508(.A1(new_n933), .A2(KEYINPUT108), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(KEYINPUT108), .ZN(new_n935));
  INV_X1    g510(.A(new_n928), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n934), .B(new_n935), .C1(new_n925), .C2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT109), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n924), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n940), .A2(new_n924), .ZN(new_n942));
  OAI21_X1  g517(.A(G868), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n943), .B1(G868), .B2(new_n866), .ZN(G295));
  OAI21_X1  g519(.A(new_n943), .B1(G868), .B2(new_n866), .ZN(G331));
  AOI22_X1  g520(.A1(new_n558), .A2(new_n550), .B1(new_n592), .B2(new_n594), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n550), .A2(new_n537), .A3(new_n558), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n864), .B1(new_n861), .B2(new_n863), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n527), .A2(new_n530), .A3(G93), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n857), .A2(KEYINPUT103), .A3(new_n859), .A4(new_n949), .ZN(new_n950));
  AOI22_X1  g525(.A1(new_n948), .A2(new_n950), .B1(new_n567), .B2(new_n568), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n871), .A2(new_n567), .A3(new_n568), .ZN(new_n952));
  OAI22_X1  g527(.A1(new_n946), .A2(new_n947), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(G171), .A2(new_n595), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n550), .A2(new_n537), .A3(new_n558), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n954), .A2(new_n870), .A3(new_n872), .A4(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n953), .A2(new_n956), .A3(new_n928), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n957), .B(KEYINPUT112), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n959), .B1(new_n953), .B2(new_n956), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n954), .A2(new_n955), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT110), .B1(new_n961), .B2(new_n873), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n932), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n932), .B(KEYINPUT111), .C1(new_n960), .C2(new_n962), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n958), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n923), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n912), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI211_X1 g544(.A(new_n923), .B(new_n958), .C1(new_n965), .C2(new_n966), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT43), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT113), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n974));
  OAI211_X1 g549(.A(KEYINPUT113), .B(KEYINPUT43), .C1(new_n969), .C2(new_n970), .ZN(new_n975));
  XOR2_X1   g550(.A(new_n957), .B(KEYINPUT112), .Z(new_n976));
  NAND2_X1  g551(.A1(new_n953), .A2(new_n956), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT110), .ZN(new_n978));
  INV_X1    g553(.A(new_n962), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT111), .B1(new_n980), .B2(new_n932), .ZN(new_n981));
  INV_X1    g556(.A(new_n966), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n968), .B(new_n976), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n936), .A2(new_n929), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n985), .B(new_n977), .C1(new_n936), .C2(new_n931), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n986), .B1(new_n980), .B2(new_n936), .ZN(new_n987));
  AOI21_X1  g562(.A(G37), .B1(new_n987), .B2(new_n923), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n983), .A2(new_n984), .A3(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n973), .A2(new_n974), .A3(new_n975), .A4(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n976), .B1(new_n981), .B2(new_n982), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n923), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n992), .A2(new_n984), .A3(new_n912), .A4(new_n983), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n983), .A2(new_n994), .A3(new_n988), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT43), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n994), .B1(new_n983), .B2(new_n988), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n993), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT44), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n990), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT115), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT115), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n990), .A2(new_n999), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(G397));
  INV_X1    g579(.A(G8), .ZN(new_n1005));
  NOR2_X1   g580(.A1(G168), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n477), .A2(G40), .A3(new_n483), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n1008));
  AOI21_X1  g583(.A(G1384), .B1(new_n901), .B2(new_n902), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n1010), .A2(new_n772), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1384), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n903), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1007), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n498), .A2(new_n500), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n901), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1018), .A2(KEYINPUT45), .A3(new_n1013), .ZN(new_n1019));
  AOI21_X1  g594(.A(G1966), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1006), .B1(new_n1012), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(G8), .B1(new_n1012), .B2(new_n1020), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1006), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT123), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1024), .A2(KEYINPUT51), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n1026));
  AOI211_X1 g601(.A(KEYINPUT123), .B(new_n1026), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1021), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT62), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1007), .B1(KEYINPUT45), .B2(new_n1009), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1015), .B1(G164), .B2(G1384), .ZN(new_n1031));
  AOI21_X1  g606(.A(G1971), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G2090), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1010), .A2(new_n1034), .A3(new_n1011), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT117), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(G303), .A2(G8), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n1038), .B(KEYINPUT55), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1033), .A2(KEYINPUT117), .A3(new_n1035), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1037), .A2(G8), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n602), .B1(KEYINPUT118), .B2(new_n605), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1043), .B1(KEYINPUT118), .B2(new_n605), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G1981), .ZN(new_n1045));
  INV_X1    g620(.A(G1981), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n606), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(KEYINPUT119), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT119), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1044), .A2(new_n1049), .A3(G1981), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT49), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1014), .A2(new_n1007), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(new_n1005), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT49), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1048), .A2(new_n1055), .A3(new_n1050), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1052), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1976), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT52), .B1(G288), .B2(new_n1058), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1054), .B(new_n1059), .C1(new_n1058), .C2(G288), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1054), .B1(new_n1058), .B2(G288), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT52), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1057), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1007), .B1(new_n1014), .B2(KEYINPUT50), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1018), .A2(new_n1008), .A3(new_n1013), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1067), .A2(G2090), .ZN(new_n1068));
  OAI21_X1  g643(.A(G8), .B1(new_n1068), .B2(new_n1032), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n1039), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1042), .A2(new_n1064), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G2078), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1030), .A2(new_n1072), .A3(new_n1031), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1075));
  INV_X1    g650(.A(G1961), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1073), .A2(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1074), .A2(G2078), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1016), .A2(new_n1019), .A3(new_n1078), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n1080), .A2(G301), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1071), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT62), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1083), .B(new_n1021), .C1(new_n1025), .C2(new_n1027), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1029), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT63), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n1063), .A2(G286), .A3(new_n1022), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1041), .A2(G8), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1039), .B1(new_n1088), .B2(new_n1036), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1086), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1022), .A2(G286), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1070), .A2(new_n1091), .A3(new_n1086), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1063), .B1(new_n1092), .B2(new_n1042), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1057), .A2(new_n1058), .A3(new_n821), .ZN(new_n1094));
  AOI211_X1 g669(.A(new_n1005), .B(new_n1053), .C1(new_n1094), .C2(new_n1047), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n1090), .A2(new_n1093), .A3(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n1097));
  XNOR2_X1  g672(.A(G299), .B(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT56), .B(G2072), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1030), .A2(new_n1031), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(G1956), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT120), .B1(new_n1067), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n1104));
  AOI211_X1 g679(.A(new_n1104), .B(G1956), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1099), .B(new_n1101), .C1(new_n1103), .C2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1053), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1107), .A2(G2067), .ZN(new_n1108));
  AOI21_X1  g683(.A(G1348), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1110), .A2(new_n625), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1106), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1101), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n1098), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(G1996), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1030), .A2(new_n1116), .A3(new_n1031), .ZN(new_n1117));
  XNOR2_X1  g692(.A(KEYINPUT58), .B(G1341), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1117), .B1(new_n1053), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT59), .B1(new_n1119), .B2(new_n570), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n625), .A2(KEYINPUT60), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1120), .B1(new_n1110), .B2(new_n1121), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1108), .A2(new_n1109), .A3(new_n632), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT60), .B1(new_n1111), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1119), .A2(KEYINPUT59), .A3(new_n570), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1122), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT61), .B1(new_n1114), .B2(new_n1106), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n1129));
  OR2_X1    g704(.A1(new_n1106), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1106), .A2(new_n1129), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1130), .A2(KEYINPUT61), .A3(new_n1131), .A4(new_n1114), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1115), .B1(new_n1128), .B2(new_n1132), .ZN(new_n1133));
  XOR2_X1   g708(.A(G171), .B(KEYINPUT54), .Z(new_n1134));
  OAI211_X1 g709(.A(new_n1016), .B(new_n1078), .C1(new_n1015), .C2(new_n1014), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1134), .B1(new_n1077), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1136), .B1(new_n1080), .B2(new_n1134), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1071), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n1028), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1085), .B(new_n1096), .C1(new_n1133), .C2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n764), .B(G2067), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1141), .B1(new_n725), .B2(new_n1116), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1007), .A2(new_n1009), .A3(KEYINPUT45), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT116), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1143), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1145), .B1(new_n1146), .B2(G1996), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1143), .A2(KEYINPUT116), .A3(new_n1116), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1144), .B1(new_n1150), .B2(new_n724), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n841), .A2(new_n843), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n841), .A2(new_n843), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1151), .B1(new_n1143), .B2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(G290), .B(G1986), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1143), .A2(new_n1157), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1140), .A2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1144), .B(new_n1152), .C1(new_n1150), .C2(new_n724), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n764), .A2(new_n766), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1146), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  XOR2_X1   g738(.A(new_n1163), .B(KEYINPUT124), .Z(new_n1164));
  XNOR2_X1  g739(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1149), .A2(KEYINPUT46), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1166), .B(KEYINPUT125), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1146), .B1(new_n725), .B2(new_n1141), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1168), .B1(new_n1149), .B2(KEYINPUT46), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1165), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1167), .A2(new_n1169), .A3(new_n1165), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1146), .A2(G1986), .A3(G290), .ZN(new_n1172));
  XOR2_X1   g747(.A(new_n1172), .B(KEYINPUT48), .Z(new_n1173));
  NAND2_X1  g748(.A1(new_n1156), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1164), .A2(new_n1170), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1160), .A2(new_n1176), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g752(.A1(G229), .A2(new_n460), .A3(G401), .A4(G227), .ZN(new_n1179));
  NAND3_X1  g753(.A1(new_n973), .A2(new_n975), .A3(new_n989), .ZN(new_n1180));
  NAND3_X1  g754(.A1(new_n918), .A2(new_n1179), .A3(new_n1180), .ZN(G225));
  INV_X1    g755(.A(G225), .ZN(G308));
endmodule


