//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 1 1 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 0 1 1 0 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT71), .ZN(new_n206));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(G211gat), .A2(G218gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n207), .B1(KEYINPUT22), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G211gat), .ZN(new_n211));
  INV_X1    g010(.A(G218gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n210), .A2(new_n208), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n208), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n215), .B(new_n207), .C1(KEYINPUT22), .C2(new_n209), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n219), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n220));
  OR2_X1    g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AND3_X1   g022(.A1(new_n220), .A2(new_n223), .A3(KEYINPUT66), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT66), .B1(new_n220), .B2(new_n223), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT28), .ZN(new_n227));
  INV_X1    g026(.A(G183gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT27), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT27), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G183gat), .ZN(new_n231));
  INV_X1    g030(.A(G190gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n229), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n227), .B1(new_n233), .B2(KEYINPUT65), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT64), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT27), .B(G183gat), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n235), .B1(new_n236), .B2(new_n232), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n234), .B1(new_n237), .B2(KEYINPUT65), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT65), .B1(new_n233), .B2(KEYINPUT64), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(new_n227), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n226), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G183gat), .A2(G190gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n242), .A2(KEYINPUT24), .ZN(new_n243));
  AND2_X1   g042(.A1(G169gat), .A2(G176gat), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT23), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n219), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n228), .A2(new_n232), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(KEYINPUT24), .A3(new_n242), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n245), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT25), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n245), .A2(new_n249), .A3(KEYINPUT25), .A4(new_n251), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n256), .ZN(new_n257));
  AND2_X1   g056(.A1(G226gat), .A2(G233gat), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n257), .A2(KEYINPUT70), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT70), .B1(new_n257), .B2(new_n258), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT29), .B1(new_n241), .B2(new_n256), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n262), .A2(new_n258), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n218), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n257), .A2(new_n258), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n265), .B(new_n217), .C1(new_n258), .C2(new_n262), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n206), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n257), .A2(KEYINPUT70), .A3(new_n258), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n263), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n206), .B(new_n266), .C1(new_n271), .C2(new_n217), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n205), .B1(new_n267), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G120gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(G113gat), .ZN(new_n276));
  INV_X1    g075(.A(G113gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(G120gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT1), .ZN(new_n280));
  INV_X1    g079(.A(G134gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(G127gat), .ZN(new_n282));
  INV_X1    g081(.A(G127gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G134gat), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n279), .A2(new_n280), .A3(new_n282), .A4(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n282), .A2(new_n284), .ZN(new_n286));
  XNOR2_X1  g085(.A(G113gat), .B(G120gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n286), .B1(new_n287), .B2(KEYINPUT1), .ZN(new_n288));
  AND2_X1   g087(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n241), .A2(new_n289), .A3(new_n256), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n289), .B1(new_n241), .B2(new_n256), .ZN(new_n291));
  INV_X1    g090(.A(G227gat), .ZN(new_n292));
  INV_X1    g091(.A(G233gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(KEYINPUT68), .A2(KEYINPUT34), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NOR4_X1   g095(.A1(new_n290), .A2(new_n291), .A3(new_n294), .A4(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n291), .ZN(new_n298));
  INV_X1    g097(.A(new_n294), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n241), .A2(new_n289), .A3(new_n256), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(KEYINPUT68), .A2(KEYINPUT34), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n297), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G15gat), .B(G43gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n306), .B(KEYINPUT67), .ZN(new_n307));
  INV_X1    g106(.A(G71gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n309), .B(G99gat), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n294), .B1(new_n290), .B2(new_n291), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT33), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(KEYINPUT32), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n311), .B(KEYINPUT32), .C1(new_n310), .C2(new_n312), .ZN(new_n316));
  AND3_X1   g115(.A1(new_n305), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n304), .ZN(new_n318));
  INV_X1    g117(.A(new_n297), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n315), .A2(new_n316), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n204), .B(new_n266), .C1(new_n271), .C2(new_n217), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT30), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n264), .A2(KEYINPUT30), .A3(new_n204), .A4(new_n266), .ZN(new_n325));
  AND2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G78gat), .B(G106gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(KEYINPUT79), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT31), .B(G50gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT81), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT29), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT3), .B1(new_n217), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT72), .ZN(new_n335));
  INV_X1    g134(.A(G148gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G141gat), .ZN(new_n337));
  INV_X1    g136(.A(G141gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(G148gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G155gat), .B(G162gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(G155gat), .A2(G162gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT2), .ZN(new_n343));
  AND4_X1   g142(.A1(new_n335), .A2(new_n340), .A3(new_n341), .A4(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT72), .B1(new_n337), .B2(new_n339), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n341), .B1(new_n345), .B2(new_n343), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  OR2_X1    g146(.A1(new_n334), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n338), .A2(G148gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n336), .A2(G141gat), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n335), .B(new_n343), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n341), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n345), .A2(new_n341), .A3(new_n343), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n333), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n356), .A2(KEYINPUT80), .A3(new_n333), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n359), .A2(new_n218), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n348), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(G228gat), .A2(G233gat), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n363), .B1(new_n334), .B2(new_n347), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n217), .B1(new_n356), .B2(new_n333), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(G22gat), .B1(new_n365), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n363), .B1(new_n348), .B2(new_n361), .ZN(new_n371));
  INV_X1    g170(.A(G22gat), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n371), .A2(new_n372), .A3(new_n368), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n332), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n365), .A2(new_n369), .A3(G22gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n330), .B(new_n331), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n372), .B1(new_n371), .B2(new_n368), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT35), .B1(new_n374), .B2(new_n378), .ZN(new_n379));
  AND4_X1   g178(.A1(new_n274), .A2(new_n321), .A3(new_n326), .A4(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G1gat), .B(G29gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(KEYINPUT0), .ZN(new_n382));
  XOR2_X1   g181(.A(G57gat), .B(G85gat), .Z(new_n383));
  XNOR2_X1  g182(.A(new_n382), .B(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT75), .ZN(new_n385));
  XOR2_X1   g184(.A(KEYINPUT74), .B(KEYINPUT4), .Z(new_n386));
  NAND4_X1  g185(.A1(new_n347), .A2(new_n385), .A3(new_n289), .A4(new_n386), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n353), .A2(new_n285), .A3(new_n355), .A4(new_n288), .ZN(new_n388));
  INV_X1    g187(.A(new_n386), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT75), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT4), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n391), .B1(new_n347), .B2(new_n289), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n387), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT76), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT76), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n395), .B(new_n387), .C1(new_n390), .C2(new_n392), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT3), .B1(new_n344), .B2(new_n346), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n285), .A2(new_n288), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(new_n398), .A3(new_n356), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT73), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT73), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n397), .A2(new_n401), .A3(new_n398), .A4(new_n356), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(G225gat), .A2(G233gat), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n405), .A2(KEYINPUT5), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n394), .A2(new_n396), .A3(new_n403), .A4(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT77), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI22_X1  g208(.A1(new_n393), .A2(KEYINPUT76), .B1(new_n400), .B2(new_n402), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n410), .A2(KEYINPUT77), .A3(new_n396), .A4(new_n406), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n388), .A2(new_n386), .ZN(new_n413));
  INV_X1    g212(.A(new_n388), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n405), .B1(new_n414), .B2(KEYINPUT4), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n403), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n347), .A2(new_n289), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n405), .B1(new_n417), .B2(new_n414), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT5), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n384), .B1(new_n412), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n413), .B(new_n404), .C1(new_n391), .C2(new_n388), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n424), .B1(new_n400), .B2(new_n402), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n384), .B1(new_n425), .B2(new_n419), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n426), .B1(new_n409), .B2(new_n411), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT78), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI22_X1  g229(.A1(new_n409), .A2(new_n411), .B1(new_n416), .B2(new_n420), .ZN(new_n431));
  OAI22_X1  g230(.A1(new_n431), .A2(new_n384), .B1(new_n427), .B2(KEYINPUT78), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n423), .A2(new_n430), .B1(new_n432), .B2(new_n429), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT84), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n380), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n426), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT78), .B1(new_n412), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n429), .B1(new_n422), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT78), .ZN(new_n439));
  AOI211_X1 g238(.A(new_n439), .B(new_n426), .C1(new_n409), .C2(new_n411), .ZN(new_n440));
  OAI22_X1  g239(.A1(new_n440), .A2(KEYINPUT6), .B1(new_n431), .B2(new_n384), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n321), .A2(new_n326), .A3(new_n274), .A4(new_n379), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT84), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n435), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n266), .B1(new_n271), .B2(new_n217), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT71), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n204), .B1(new_n447), .B2(new_n272), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n324), .A2(new_n325), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n438), .A2(new_n450), .A3(new_n441), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n374), .A2(new_n378), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT69), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n317), .A2(new_n320), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n320), .A2(new_n453), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n452), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT35), .B1(new_n451), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT37), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n459), .B1(new_n447), .B2(new_n272), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n205), .B1(new_n446), .B2(KEYINPUT37), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT38), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT83), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI211_X1 g263(.A(KEYINPUT83), .B(KEYINPUT38), .C1(new_n460), .C2(new_n461), .ZN(new_n465));
  INV_X1    g264(.A(new_n322), .ZN(new_n466));
  INV_X1    g265(.A(new_n461), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n263), .B1(new_n258), .B2(new_n257), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n459), .B1(new_n468), .B2(new_n218), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n217), .B1(new_n261), .B2(new_n263), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT38), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n466), .B1(new_n467), .B2(new_n471), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n464), .A2(new_n442), .A3(new_n465), .A4(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n452), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n450), .A2(new_n422), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n394), .A2(new_n396), .A3(new_n403), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n405), .ZN(new_n477));
  OR2_X1    g276(.A1(new_n477), .A2(KEYINPUT39), .ZN(new_n478));
  OR2_X1    g277(.A1(new_n417), .A2(new_n414), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n477), .B(KEYINPUT39), .C1(new_n405), .C2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n480), .A3(new_n384), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT82), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n481), .B1(new_n482), .B2(KEYINPUT40), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(KEYINPUT40), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n478), .A2(new_n480), .A3(new_n384), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n474), .B1(new_n475), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n473), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n315), .A2(new_n316), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n319), .A2(new_n318), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n305), .A2(new_n315), .A3(new_n316), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(KEYINPUT69), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n493), .A2(KEYINPUT36), .A3(new_n455), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT36), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n321), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n497), .B1(new_n474), .B2(new_n451), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n445), .A2(new_n458), .B1(new_n488), .B2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G15gat), .B(G22gat), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT16), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n500), .B1(new_n501), .B2(G1gat), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n502), .B1(G1gat), .B2(new_n500), .ZN(new_n503));
  OR2_X1    g302(.A1(new_n503), .A2(G8gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(G8gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(G29gat), .A2(G36gat), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NOR3_X1   g308(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(G43gat), .B(G50gat), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(KEYINPUT15), .A3(new_n512), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n512), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n514), .B1(KEYINPUT15), .B2(new_n512), .ZN(new_n515));
  OR2_X1    g314(.A1(new_n510), .A2(KEYINPUT86), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n510), .A2(KEYINPUT86), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n509), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n513), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT17), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT17), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n521), .B(new_n513), .C1(new_n515), .C2(new_n518), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n506), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  OR2_X1    g322(.A1(new_n515), .A2(new_n518), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n524), .A2(new_n513), .B1(new_n504), .B2(new_n505), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT18), .ZN(new_n526));
  NAND2_X1  g325(.A1(G229gat), .A2(G233gat), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NOR4_X1   g327(.A1(new_n523), .A2(new_n525), .A3(new_n526), .A4(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n527), .B(KEYINPUT13), .Z(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n506), .ZN(new_n532));
  INV_X1    g331(.A(new_n519), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n525), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n531), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT87), .B1(new_n529), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n532), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n539), .A2(new_n535), .A3(new_n527), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n526), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n506), .B(new_n519), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n530), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n539), .A2(new_n535), .A3(KEYINPUT18), .A4(new_n527), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT87), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n537), .A2(new_n541), .A3(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G113gat), .B(G141gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(G197gat), .ZN(new_n549));
  XOR2_X1   g348(.A(KEYINPUT11), .B(G169gat), .Z(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(KEYINPUT12), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n552), .B(KEYINPUT85), .Z(new_n553));
  AND3_X1   g352(.A1(new_n540), .A2(KEYINPUT88), .A3(new_n526), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT88), .B1(new_n540), .B2(new_n526), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AND3_X1   g355(.A1(new_n543), .A2(new_n544), .A3(new_n552), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n547), .A2(new_n553), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n499), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(KEYINPUT91), .B(G64gat), .ZN(new_n560));
  INV_X1    g359(.A(G57gat), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT92), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n561), .A2(G64gat), .ZN(new_n564));
  OR3_X1    g363(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G71gat), .A2(G78gat), .ZN(new_n566));
  INV_X1    g365(.A(G78gat), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n308), .A2(new_n567), .A3(KEYINPUT9), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n562), .A2(new_n563), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n561), .A2(G64gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n566), .ZN(new_n572));
  OAI22_X1  g371(.A1(new_n564), .A2(new_n571), .B1(new_n572), .B2(KEYINPUT9), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n566), .B(KEYINPUT89), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n308), .A2(new_n567), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT90), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n573), .A2(new_n574), .A3(KEYINPUT90), .A4(new_n575), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n570), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(KEYINPUT93), .B(KEYINPUT21), .Z(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n583), .B(new_n584), .Z(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(G127gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n583), .B(new_n584), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n283), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT21), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n532), .B1(new_n581), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT94), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n586), .A2(new_n588), .A3(new_n592), .ZN(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(G155gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(G183gat), .B(G211gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n594), .A2(new_n595), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n599), .B1(new_n594), .B2(new_n595), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G190gat), .B(G218gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(G134gat), .B(G162gat), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n603), .B(new_n604), .Z(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(KEYINPUT95), .A2(G85gat), .A3(G92gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT7), .ZN(new_n608));
  INV_X1    g407(.A(G99gat), .ZN(new_n609));
  INV_X1    g408(.A(G106gat), .ZN(new_n610));
  OAI21_X1  g409(.A(KEYINPUT8), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT96), .B(G92gat), .ZN(new_n612));
  INV_X1    g411(.A(G85gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n608), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(G99gat), .B(G106gat), .Z(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT97), .ZN(new_n618));
  INV_X1    g417(.A(new_n616), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n619), .A2(new_n608), .A3(new_n611), .A4(new_n614), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n617), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n620), .A2(new_n618), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(new_n519), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G232gat), .A2(G233gat), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT41), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(KEYINPUT98), .B1(new_n625), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT98), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n624), .B(new_n630), .C1(new_n627), .C2(new_n626), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n621), .A2(new_n622), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n538), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n626), .A2(new_n627), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n632), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n635), .B1(new_n632), .B2(new_n634), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n606), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n632), .A2(new_n634), .ZN(new_n640));
  INV_X1    g439(.A(new_n635), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n642), .A2(new_n636), .A3(new_n605), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n602), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n570), .A2(new_n580), .A3(new_n620), .A4(new_n617), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT10), .ZN(new_n647));
  INV_X1    g446(.A(new_n581), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n646), .B(new_n647), .C1(new_n648), .C2(new_n623), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n570), .A2(new_n580), .A3(KEYINPUT10), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n623), .ZN(new_n651));
  AOI22_X1  g450(.A1(new_n649), .A2(new_n651), .B1(G230gat), .B2(G233gat), .ZN(new_n652));
  NAND2_X1  g451(.A1(G230gat), .A2(G233gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n633), .A2(new_n581), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n653), .B1(new_n654), .B2(new_n646), .ZN(new_n655));
  XOR2_X1   g454(.A(G120gat), .B(G148gat), .Z(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT99), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n657), .B(KEYINPUT100), .Z(new_n658));
  XNOR2_X1  g457(.A(G176gat), .B(G204gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  OR3_X1    g459(.A1(new_n652), .A2(new_n655), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n660), .B1(new_n652), .B2(new_n655), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n645), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n559), .A2(new_n442), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g465(.A1(new_n559), .A2(new_n664), .ZN(new_n667));
  INV_X1    g466(.A(new_n450), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT16), .B(G8gat), .Z(new_n669));
  AND3_X1   g468(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(G8gat), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n671), .B1(new_n667), .B2(new_n668), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT42), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n673), .B1(KEYINPUT42), .B2(new_n670), .ZN(G1325gat));
  AOI21_X1  g473(.A(G15gat), .B1(new_n667), .B2(new_n321), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n494), .A2(KEYINPUT101), .A3(new_n496), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT101), .B1(new_n494), .B2(new_n496), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(G15gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT102), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n675), .B1(new_n667), .B2(new_n680), .ZN(G1326gat));
  XNOR2_X1  g480(.A(KEYINPUT43), .B(G22gat), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n474), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT103), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n684), .A2(KEYINPUT103), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n683), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n687), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n689), .A2(new_n685), .A3(new_n682), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(G1327gat));
  NAND2_X1  g490(.A1(new_n488), .A2(new_n498), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n458), .A2(new_n444), .A3(new_n435), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n644), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n602), .A2(new_n558), .A3(new_n663), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(G29gat), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n696), .A2(new_n697), .A3(new_n442), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT45), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(new_n499), .B2(new_n644), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n692), .A2(new_n693), .ZN(new_n703));
  INV_X1    g502(.A(new_n644), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(KEYINPUT44), .A3(new_n704), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n702), .A2(new_n442), .A3(new_n705), .A4(new_n695), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(G29gat), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n696), .A2(KEYINPUT45), .A3(new_n697), .A4(new_n442), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n700), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT104), .ZN(G1328gat));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n712));
  AOI211_X1 g511(.A(G36gat), .B(new_n450), .C1(new_n712), .C2(KEYINPUT46), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n712), .A2(KEYINPUT46), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n714), .B(new_n716), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n702), .A2(new_n668), .A3(new_n705), .A4(new_n695), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(G36gat), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n711), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n714), .B(new_n715), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n722), .A2(KEYINPUT106), .A3(new_n719), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(G1329gat));
  INV_X1    g523(.A(G43gat), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n696), .A2(new_n725), .A3(new_n321), .ZN(new_n726));
  AND4_X1   g525(.A1(new_n497), .A2(new_n702), .A3(new_n695), .A4(new_n705), .ZN(new_n727));
  OAI211_X1 g526(.A(KEYINPUT47), .B(new_n726), .C1(new_n727), .C2(new_n725), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n702), .A2(new_n678), .A3(new_n705), .A4(new_n695), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(G43gat), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT47), .B1(new_n730), .B2(new_n726), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(KEYINPUT107), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n733));
  AOI211_X1 g532(.A(new_n733), .B(KEYINPUT47), .C1(new_n730), .C2(new_n726), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n728), .B1(new_n732), .B2(new_n734), .ZN(G1330gat));
  INV_X1    g534(.A(G50gat), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n702), .A2(new_n474), .A3(new_n705), .A4(new_n695), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n736), .B1(new_n737), .B2(KEYINPUT108), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(KEYINPUT108), .B2(new_n737), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n696), .A2(new_n736), .A3(new_n474), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n739), .A2(KEYINPUT48), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n737), .A2(G50gat), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n740), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT48), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n741), .A2(new_n745), .ZN(G1331gat));
  INV_X1    g545(.A(new_n558), .ZN(new_n747));
  INV_X1    g546(.A(new_n663), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n645), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n703), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(new_n433), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(new_n561), .ZN(G1332gat));
  INV_X1    g551(.A(KEYINPUT109), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n750), .B(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n668), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n755), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n756));
  XOR2_X1   g555(.A(KEYINPUT49), .B(G64gat), .Z(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(new_n755), .B2(new_n757), .ZN(G1333gat));
  NAND3_X1  g557(.A1(new_n754), .A2(G71gat), .A3(new_n678), .ZN(new_n759));
  INV_X1    g558(.A(new_n321), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n308), .B1(new_n750), .B2(new_n760), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n759), .A2(KEYINPUT50), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT50), .B1(new_n759), .B2(new_n761), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(G1334gat));
  NAND2_X1  g563(.A1(new_n754), .A2(new_n474), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g565(.A1(new_n602), .A2(new_n747), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n451), .A2(new_n474), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n494), .A2(new_n496), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n473), .B2(new_n487), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n458), .A2(new_n444), .A3(new_n435), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n704), .B(new_n767), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n694), .A2(KEYINPUT51), .A3(new_n767), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n748), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n777), .A2(new_n613), .A3(new_n442), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n602), .A2(new_n747), .A3(new_n748), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n702), .A2(new_n705), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT110), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT110), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n702), .A2(new_n782), .A3(new_n705), .A4(new_n779), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n781), .A2(new_n442), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n778), .B1(new_n784), .B2(new_n613), .ZN(G1336gat));
  NOR2_X1   g584(.A1(new_n450), .A2(G92gat), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n777), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT112), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n777), .A2(new_n789), .A3(new_n786), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n702), .A2(new_n668), .A3(new_n705), .A4(new_n779), .ZN(new_n791));
  INV_X1    g590(.A(new_n612), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT52), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n788), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n775), .A2(new_n795), .A3(new_n776), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n773), .A2(KEYINPUT111), .A3(new_n774), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n786), .A2(new_n663), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n796), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n781), .A2(new_n668), .A3(new_n783), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n800), .B1(new_n792), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n794), .B1(new_n802), .B2(new_n803), .ZN(G1337gat));
  NAND3_X1  g603(.A1(new_n777), .A2(new_n609), .A3(new_n321), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n781), .A2(new_n678), .A3(new_n783), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n805), .B1(new_n806), .B2(new_n609), .ZN(G1338gat));
  NAND2_X1  g606(.A1(new_n775), .A2(new_n776), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n748), .A2(new_n452), .A3(G106gat), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT53), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(G106gat), .B1(new_n780), .B2(new_n452), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n796), .A2(new_n797), .A3(new_n809), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n781), .A2(new_n474), .A3(new_n783), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n813), .B1(G106gat), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n812), .B1(new_n815), .B2(new_n816), .ZN(G1339gat));
  NAND4_X1  g616(.A1(new_n602), .A2(new_n558), .A3(new_n644), .A4(new_n748), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n652), .A2(new_n655), .A3(new_n660), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n649), .A2(new_n651), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n653), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n653), .B1(new_n650), .B2(new_n623), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n823), .B1(new_n649), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n820), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n660), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n827), .B1(new_n652), .B2(new_n823), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n819), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n821), .A2(new_n823), .A3(new_n653), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n649), .A2(new_n824), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT54), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n830), .B(new_n660), .C1(new_n832), .C2(new_n652), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n820), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n829), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n556), .A2(new_n557), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n542), .A2(new_n530), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n527), .B1(new_n539), .B2(new_n535), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n551), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n644), .A2(new_n835), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n663), .A2(new_n836), .A3(new_n839), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n842), .B1(new_n835), .B2(new_n558), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT113), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n704), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n842), .B(KEYINPUT113), .C1(new_n835), .C2(new_n558), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n841), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n818), .B1(new_n847), .B2(new_n602), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n493), .A2(new_n455), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n848), .A2(new_n442), .A3(new_n452), .A4(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT115), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n668), .B1(new_n850), .B2(new_n851), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(KEYINPUT116), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n856), .B1(new_n852), .B2(new_n853), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n277), .B(new_n747), .C1(new_n855), .C2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n602), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n860), .A2(new_n644), .A3(new_n846), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n859), .B1(new_n861), .B2(new_n841), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n474), .B1(new_n862), .B2(new_n818), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n863), .A2(new_n442), .A3(new_n450), .A4(new_n321), .ZN(new_n864));
  OAI21_X1  g663(.A(G113gat), .B1(new_n864), .B2(new_n558), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT114), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n865), .B(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n858), .A2(new_n867), .ZN(G1340gat));
  OAI211_X1 g667(.A(new_n275), .B(new_n663), .C1(new_n855), .C2(new_n857), .ZN(new_n869));
  OAI21_X1  g668(.A(G120gat), .B1(new_n864), .B2(new_n748), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(G1341gat));
  OAI21_X1  g670(.A(G127gat), .B1(new_n864), .B2(new_n859), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n602), .A2(new_n283), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n854), .B2(new_n873), .ZN(G1342gat));
  NOR2_X1   g673(.A1(new_n644), .A2(G134gat), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  OR3_X1    g675(.A1(new_n854), .A2(KEYINPUT56), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(G134gat), .B1(new_n864), .B2(new_n644), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT56), .B1(new_n854), .B2(new_n876), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(G1343gat));
  NAND2_X1  g679(.A1(new_n442), .A2(new_n450), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(new_n497), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  OR3_X1    g682(.A1(new_n644), .A2(new_n835), .A3(new_n840), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n843), .A2(new_n644), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n602), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(new_n818), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n888), .A2(new_n889), .A3(new_n452), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT57), .B1(new_n848), .B2(new_n474), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n452), .B1(new_n862), .B2(new_n818), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT117), .B1(new_n894), .B2(KEYINPUT57), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n883), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n338), .B1(new_n896), .B2(new_n747), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n898));
  INV_X1    g697(.A(new_n678), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n894), .A2(new_n442), .A3(new_n450), .A4(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n558), .A2(G141gat), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n898), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT58), .B1(new_n897), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n848), .A2(new_n474), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n905), .A2(new_n892), .A3(new_n889), .ZN(new_n906));
  INV_X1    g705(.A(new_n890), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n891), .A2(new_n892), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n747), .B(new_n882), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(G141gat), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT58), .ZN(new_n912));
  INV_X1    g711(.A(new_n903), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n904), .A2(new_n914), .ZN(G1344gat));
  INV_X1    g714(.A(new_n900), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n336), .A3(new_n663), .ZN(new_n917));
  AOI211_X1 g716(.A(KEYINPUT59), .B(new_n336), .C1(new_n896), .C2(new_n663), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n452), .A2(new_n889), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n848), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n889), .B1(new_n888), .B2(new_n452), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n883), .A2(new_n748), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n336), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT59), .ZN(new_n925));
  OR3_X1    g724(.A1(new_n924), .A2(KEYINPUT119), .A3(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(KEYINPUT119), .B1(new_n924), .B2(new_n925), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n917), .B1(new_n918), .B2(new_n928), .ZN(G1345gat));
  INV_X1    g728(.A(KEYINPUT120), .ZN(new_n930));
  INV_X1    g729(.A(G155gat), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n931), .B1(new_n896), .B2(new_n602), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n900), .A2(G155gat), .A3(new_n859), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n602), .B(new_n882), .C1(new_n908), .C2(new_n909), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G155gat), .ZN(new_n936));
  INV_X1    g735(.A(new_n933), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(KEYINPUT120), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n934), .A2(new_n938), .ZN(G1346gat));
  AOI21_X1  g738(.A(G162gat), .B1(new_n916), .B2(new_n704), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n704), .A2(G162gat), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n896), .B2(new_n941), .ZN(G1347gat));
  INV_X1    g741(.A(new_n457), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n943), .A2(new_n668), .A3(KEYINPUT121), .ZN(new_n944));
  AOI21_X1  g743(.A(KEYINPUT121), .B1(new_n943), .B2(new_n668), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n944), .A2(new_n945), .A3(new_n442), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n848), .A2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(G169gat), .B1(new_n948), .B2(new_n747), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n442), .A2(new_n760), .A3(new_n450), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n863), .A2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n747), .A2(G169gat), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(G1348gat));
  OAI21_X1  g753(.A(G176gat), .B1(new_n951), .B2(new_n748), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n748), .A2(G176gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n947), .B2(new_n956), .ZN(G1349gat));
  OAI21_X1  g756(.A(G183gat), .B1(new_n951), .B2(new_n859), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n948), .A2(new_n236), .A3(new_n602), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g760(.A1(new_n948), .A2(new_n232), .A3(new_n704), .ZN(new_n962));
  OAI21_X1  g761(.A(G190gat), .B1(new_n951), .B2(new_n644), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n963), .A2(KEYINPUT61), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n963), .A2(KEYINPUT61), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(G1351gat));
  NAND2_X1  g765(.A1(new_n433), .A2(new_n668), .ZN(new_n967));
  OR3_X1    g766(.A1(new_n678), .A2(KEYINPUT122), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(KEYINPUT122), .B1(new_n678), .B2(new_n967), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n922), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g770(.A(G197gat), .B1(new_n971), .B2(new_n558), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n678), .A2(new_n442), .A3(new_n450), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n894), .A2(new_n973), .ZN(new_n974));
  OR3_X1    g773(.A1(new_n974), .A2(G197gat), .A3(new_n558), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n976), .B(KEYINPUT123), .ZN(G1352gat));
  NOR3_X1   g776(.A1(new_n974), .A2(G204gat), .A3(new_n748), .ZN(new_n978));
  XNOR2_X1  g777(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n978), .B(new_n979), .ZN(new_n980));
  OAI21_X1  g779(.A(G204gat), .B1(new_n971), .B2(new_n748), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(G1353gat));
  NAND3_X1  g781(.A1(new_n922), .A2(new_n602), .A3(new_n970), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(G211gat), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT63), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n983), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n986), .A2(KEYINPUT125), .A3(new_n987), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n894), .A2(new_n211), .A3(new_n602), .A4(new_n973), .ZN(new_n989));
  OAI211_X1 g788(.A(new_n988), .B(new_n989), .C1(KEYINPUT125), .C2(new_n986), .ZN(G1354gat));
  NOR2_X1   g789(.A1(new_n971), .A2(KEYINPUT127), .ZN(new_n991));
  NOR3_X1   g790(.A1(new_n991), .A2(new_n212), .A3(new_n644), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n971), .A2(KEYINPUT127), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n212), .B1(new_n974), .B2(new_n644), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT126), .ZN(new_n995));
  OR2_X1    g794(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n994), .A2(new_n995), .ZN(new_n997));
  AOI22_X1  g796(.A1(new_n992), .A2(new_n993), .B1(new_n996), .B2(new_n997), .ZN(G1355gat));
endmodule


