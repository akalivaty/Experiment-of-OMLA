

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U552 ( .A(n604), .B(KEYINPUT95), .ZN(n638) );
  NOR2_X1 U553 ( .A1(n544), .A2(G2105), .ZN(n992) );
  NOR2_X4 U554 ( .A1(G2104), .A2(G2105), .ZN(n547) );
  XNOR2_X1 U555 ( .A(n688), .B(n687), .ZN(n689) );
  INV_X1 U556 ( .A(KEYINPUT101), .ZN(n687) );
  INV_X1 U557 ( .A(KEYINPUT66), .ZN(n592) );
  XNOR2_X2 U558 ( .A(n549), .B(KEYINPUT64), .ZN(n710) );
  NAND2_X1 U559 ( .A1(n766), .A2(n765), .ZN(n768) );
  NOR2_X2 U560 ( .A1(n599), .A2(n598), .ZN(n769) );
  NAND2_X1 U561 ( .A1(n698), .A2(KEYINPUT33), .ZN(n519) );
  INV_X1 U562 ( .A(KEYINPUT30), .ZN(n656) );
  XNOR2_X1 U563 ( .A(n686), .B(KEYINPUT100), .ZN(n701) );
  NOR2_X1 U564 ( .A1(G164), .A2(G1384), .ZN(n721) );
  INV_X1 U565 ( .A(G2105), .ZN(n548) );
  NOR2_X1 U566 ( .A1(G651), .A2(n528), .ZN(n802) );
  INV_X1 U567 ( .A(KEYINPUT40), .ZN(n767) );
  BUF_X1 U568 ( .A(n769), .Z(G160) );
  XOR2_X1 U569 ( .A(G543), .B(KEYINPUT0), .Z(n528) );
  NAND2_X1 U570 ( .A1(G49), .A2(n802), .ZN(n520) );
  XNOR2_X1 U571 ( .A(n520), .B(KEYINPUT80), .ZN(n526) );
  INV_X1 U572 ( .A(G651), .ZN(n527) );
  NOR2_X1 U573 ( .A1(G543), .A2(n527), .ZN(n521) );
  XOR2_X1 U574 ( .A(KEYINPUT1), .B(n521), .Z(n803) );
  NAND2_X1 U575 ( .A1(G87), .A2(n528), .ZN(n523) );
  NAND2_X1 U576 ( .A1(G74), .A2(G651), .ZN(n522) );
  NAND2_X1 U577 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U578 ( .A1(n803), .A2(n524), .ZN(n525) );
  NAND2_X1 U579 ( .A1(n526), .A2(n525), .ZN(G288) );
  NOR2_X1 U580 ( .A1(G651), .A2(G543), .ZN(n798) );
  NAND2_X1 U581 ( .A1(G88), .A2(n798), .ZN(n530) );
  NOR2_X1 U582 ( .A1(n528), .A2(n527), .ZN(n796) );
  NAND2_X1 U583 ( .A1(G75), .A2(n796), .ZN(n529) );
  NAND2_X1 U584 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U585 ( .A(KEYINPUT82), .B(n531), .ZN(n535) );
  NAND2_X1 U586 ( .A1(G50), .A2(n802), .ZN(n533) );
  NAND2_X1 U587 ( .A1(G62), .A2(n803), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U589 ( .A1(n535), .A2(n534), .ZN(G166) );
  INV_X1 U590 ( .A(G166), .ZN(G303) );
  NAND2_X1 U591 ( .A1(G53), .A2(n802), .ZN(n537) );
  NAND2_X1 U592 ( .A1(G65), .A2(n803), .ZN(n536) );
  NAND2_X1 U593 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U594 ( .A(KEYINPUT70), .B(n538), .Z(n542) );
  NAND2_X1 U595 ( .A1(G91), .A2(n798), .ZN(n540) );
  NAND2_X1 U596 ( .A1(G78), .A2(n796), .ZN(n539) );
  AND2_X1 U597 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n542), .A2(n541), .ZN(G299) );
  INV_X1 U599 ( .A(G2104), .ZN(n544) );
  NOR2_X2 U600 ( .A1(n544), .A2(n548), .ZN(n989) );
  NAND2_X1 U601 ( .A1(n989), .A2(G114), .ZN(n543) );
  XNOR2_X1 U602 ( .A(n543), .B(KEYINPUT84), .ZN(n546) );
  NAND2_X1 U603 ( .A1(G102), .A2(n992), .ZN(n545) );
  NAND2_X1 U604 ( .A1(n546), .A2(n545), .ZN(n553) );
  XOR2_X2 U605 ( .A(KEYINPUT17), .B(n547), .Z(n993) );
  NAND2_X1 U606 ( .A1(G138), .A2(n993), .ZN(n551) );
  NOR2_X1 U607 ( .A1(n548), .A2(G2104), .ZN(n549) );
  NAND2_X1 U608 ( .A1(G126), .A2(n710), .ZN(n550) );
  NAND2_X1 U609 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U610 ( .A1(n553), .A2(n552), .ZN(G164) );
  NAND2_X1 U611 ( .A1(G52), .A2(n802), .ZN(n555) );
  NAND2_X1 U612 ( .A1(G64), .A2(n803), .ZN(n554) );
  NAND2_X1 U613 ( .A1(n555), .A2(n554), .ZN(n561) );
  NAND2_X1 U614 ( .A1(G90), .A2(n798), .ZN(n557) );
  NAND2_X1 U615 ( .A1(G77), .A2(n796), .ZN(n556) );
  NAND2_X1 U616 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U617 ( .A(KEYINPUT68), .B(n558), .Z(n559) );
  XNOR2_X1 U618 ( .A(KEYINPUT9), .B(n559), .ZN(n560) );
  NOR2_X1 U619 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U620 ( .A(KEYINPUT69), .B(n562), .ZN(G301) );
  INV_X1 U621 ( .A(G301), .ZN(G171) );
  NAND2_X1 U622 ( .A1(G89), .A2(n798), .ZN(n563) );
  XOR2_X1 U623 ( .A(KEYINPUT4), .B(n563), .Z(n564) );
  XNOR2_X1 U624 ( .A(n564), .B(KEYINPUT73), .ZN(n566) );
  NAND2_X1 U625 ( .A1(G76), .A2(n796), .ZN(n565) );
  NAND2_X1 U626 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U627 ( .A(n567), .B(KEYINPUT5), .ZN(n572) );
  NAND2_X1 U628 ( .A1(G51), .A2(n802), .ZN(n569) );
  NAND2_X1 U629 ( .A1(G63), .A2(n803), .ZN(n568) );
  NAND2_X1 U630 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U631 ( .A(KEYINPUT6), .B(n570), .Z(n571) );
  NAND2_X1 U632 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U633 ( .A(n573), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U634 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U635 ( .A1(G73), .A2(n796), .ZN(n574) );
  XNOR2_X1 U636 ( .A(n574), .B(KEYINPUT2), .ZN(n581) );
  NAND2_X1 U637 ( .A1(G86), .A2(n798), .ZN(n576) );
  NAND2_X1 U638 ( .A1(G48), .A2(n802), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n576), .A2(n575), .ZN(n579) );
  NAND2_X1 U640 ( .A1(G61), .A2(n803), .ZN(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT81), .B(n577), .ZN(n578) );
  NOR2_X1 U642 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n581), .A2(n580), .ZN(G305) );
  NAND2_X1 U644 ( .A1(G47), .A2(n802), .ZN(n583) );
  NAND2_X1 U645 ( .A1(G60), .A2(n803), .ZN(n582) );
  NAND2_X1 U646 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U647 ( .A1(G85), .A2(n798), .ZN(n585) );
  NAND2_X1 U648 ( .A1(G72), .A2(n796), .ZN(n584) );
  NAND2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U650 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U651 ( .A(n588), .B(KEYINPUT67), .ZN(G290) );
  NOR2_X1 U652 ( .A1(G1976), .A2(G288), .ZN(n691) );
  NOR2_X1 U653 ( .A1(G1971), .A2(G303), .ZN(n589) );
  NOR2_X1 U654 ( .A1(n691), .A2(n589), .ZN(n873) );
  INV_X1 U655 ( .A(n721), .ZN(n600) );
  NAND2_X1 U656 ( .A1(n993), .A2(G137), .ZN(n591) );
  NAND2_X1 U657 ( .A1(G113), .A2(n989), .ZN(n590) );
  NAND2_X1 U658 ( .A1(n591), .A2(n590), .ZN(n593) );
  XNOR2_X1 U659 ( .A(n593), .B(n592), .ZN(n596) );
  NAND2_X1 U660 ( .A1(n710), .A2(G125), .ZN(n594) );
  XOR2_X1 U661 ( .A(KEYINPUT65), .B(n594), .Z(n595) );
  NAND2_X1 U662 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U663 ( .A1(G101), .A2(n992), .ZN(n597) );
  XNOR2_X1 U664 ( .A(KEYINPUT23), .B(n597), .ZN(n598) );
  NAND2_X1 U665 ( .A1(n769), .A2(G40), .ZN(n720) );
  NOR2_X2 U666 ( .A1(n600), .A2(n720), .ZN(n644) );
  XNOR2_X1 U667 ( .A(n644), .B(KEYINPUT93), .ZN(n646) );
  INV_X1 U668 ( .A(n646), .ZN(n629) );
  NAND2_X1 U669 ( .A1(n629), .A2(G2072), .ZN(n601) );
  XNOR2_X1 U670 ( .A(n601), .B(KEYINPUT27), .ZN(n603) );
  AND2_X1 U671 ( .A1(G1956), .A2(n646), .ZN(n602) );
  NOR2_X1 U672 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X2 U673 ( .A1(G299), .A2(n638), .ZN(n606) );
  INV_X1 U674 ( .A(KEYINPUT96), .ZN(n605) );
  XNOR2_X1 U675 ( .A(n606), .B(n605), .ZN(n637) );
  NAND2_X1 U676 ( .A1(G92), .A2(n798), .ZN(n608) );
  NAND2_X1 U677 ( .A1(G79), .A2(n796), .ZN(n607) );
  NAND2_X1 U678 ( .A1(n608), .A2(n607), .ZN(n612) );
  NAND2_X1 U679 ( .A1(G54), .A2(n802), .ZN(n610) );
  NAND2_X1 U680 ( .A1(G66), .A2(n803), .ZN(n609) );
  NAND2_X1 U681 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U683 ( .A(KEYINPUT15), .B(n613), .ZN(n1015) );
  INV_X1 U684 ( .A(n1015), .ZN(n869) );
  NAND2_X1 U685 ( .A1(n798), .A2(G81), .ZN(n614) );
  XNOR2_X1 U686 ( .A(n614), .B(KEYINPUT12), .ZN(n616) );
  NAND2_X1 U687 ( .A1(G68), .A2(n796), .ZN(n615) );
  NAND2_X1 U688 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U689 ( .A(n617), .B(KEYINPUT13), .ZN(n619) );
  NAND2_X1 U690 ( .A1(G43), .A2(n802), .ZN(n618) );
  NAND2_X1 U691 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U692 ( .A1(n803), .A2(G56), .ZN(n620) );
  XOR2_X1 U693 ( .A(KEYINPUT14), .B(n620), .Z(n621) );
  NOR2_X1 U694 ( .A1(n622), .A2(n621), .ZN(n623) );
  XOR2_X1 U695 ( .A(KEYINPUT72), .B(n623), .Z(n880) );
  INV_X1 U696 ( .A(n644), .ZN(n671) );
  INV_X1 U697 ( .A(G1996), .ZN(n978) );
  NOR2_X1 U698 ( .A1(n671), .A2(n978), .ZN(n624) );
  XOR2_X1 U699 ( .A(n624), .B(KEYINPUT26), .Z(n626) );
  NAND2_X1 U700 ( .A1(n671), .A2(G1341), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U702 ( .A1(n880), .A2(n627), .ZN(n628) );
  OR2_X1 U703 ( .A1(n869), .A2(n628), .ZN(n635) );
  NAND2_X1 U704 ( .A1(n869), .A2(n628), .ZN(n633) );
  NAND2_X1 U705 ( .A1(G2067), .A2(n629), .ZN(n631) );
  NAND2_X1 U706 ( .A1(G1348), .A2(n671), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U708 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U709 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U710 ( .A1(n637), .A2(n636), .ZN(n641) );
  NAND2_X1 U711 ( .A1(G299), .A2(n638), .ZN(n639) );
  XNOR2_X1 U712 ( .A(n639), .B(KEYINPUT28), .ZN(n640) );
  NAND2_X1 U713 ( .A1(n641), .A2(n640), .ZN(n643) );
  XNOR2_X1 U714 ( .A(KEYINPUT29), .B(KEYINPUT97), .ZN(n642) );
  XNOR2_X1 U715 ( .A(n643), .B(n642), .ZN(n668) );
  NOR2_X1 U716 ( .A1(n644), .A2(G1961), .ZN(n645) );
  XNOR2_X1 U717 ( .A(n645), .B(KEYINPUT92), .ZN(n648) );
  XOR2_X1 U718 ( .A(G2078), .B(KEYINPUT25), .Z(n848) );
  NOR2_X1 U719 ( .A1(n646), .A2(n848), .ZN(n647) );
  NOR2_X1 U720 ( .A1(n648), .A2(n647), .ZN(n649) );
  XOR2_X1 U721 ( .A(KEYINPUT94), .B(n649), .Z(n659) );
  NAND2_X1 U722 ( .A1(n659), .A2(G171), .ZN(n666) );
  NOR2_X1 U723 ( .A1(G2084), .A2(n671), .ZN(n653) );
  AND2_X1 U724 ( .A1(G8), .A2(n653), .ZN(n650) );
  NAND2_X1 U725 ( .A1(G8), .A2(n671), .ZN(n706) );
  NOR2_X1 U726 ( .A1(G1966), .A2(n706), .ZN(n654) );
  OR2_X1 U727 ( .A1(n650), .A2(n654), .ZN(n663) );
  INV_X1 U728 ( .A(n663), .ZN(n651) );
  AND2_X1 U729 ( .A1(n666), .A2(n651), .ZN(n652) );
  NAND2_X1 U730 ( .A1(n668), .A2(n652), .ZN(n665) );
  NOR2_X1 U731 ( .A1(n654), .A2(n653), .ZN(n655) );
  AND2_X1 U732 ( .A1(n655), .A2(G8), .ZN(n657) );
  XNOR2_X1 U733 ( .A(n657), .B(n656), .ZN(n658) );
  NOR2_X1 U734 ( .A1(G168), .A2(n658), .ZN(n661) );
  NOR2_X1 U735 ( .A1(G171), .A2(n659), .ZN(n660) );
  NOR2_X1 U736 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U737 ( .A(KEYINPUT31), .B(n662), .Z(n669) );
  OR2_X1 U738 ( .A1(n663), .A2(n669), .ZN(n664) );
  AND2_X1 U739 ( .A1(n665), .A2(n664), .ZN(n685) );
  AND2_X1 U740 ( .A1(n666), .A2(G286), .ZN(n667) );
  NAND2_X1 U741 ( .A1(n668), .A2(n667), .ZN(n681) );
  INV_X1 U742 ( .A(G286), .ZN(n670) );
  OR2_X1 U743 ( .A1(n670), .A2(n669), .ZN(n679) );
  INV_X1 U744 ( .A(G8), .ZN(n677) );
  NOR2_X1 U745 ( .A1(G1971), .A2(n706), .ZN(n673) );
  NOR2_X1 U746 ( .A1(G2090), .A2(n671), .ZN(n672) );
  NOR2_X1 U747 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U748 ( .A1(n674), .A2(G303), .ZN(n675) );
  XNOR2_X1 U749 ( .A(n675), .B(KEYINPUT98), .ZN(n676) );
  OR2_X1 U750 ( .A1(n677), .A2(n676), .ZN(n678) );
  AND2_X1 U751 ( .A1(n679), .A2(n678), .ZN(n680) );
  AND2_X1 U752 ( .A1(n681), .A2(n680), .ZN(n683) );
  XOR2_X1 U753 ( .A(KEYINPUT99), .B(KEYINPUT32), .Z(n682) );
  XNOR2_X1 U754 ( .A(n683), .B(n682), .ZN(n684) );
  NAND2_X1 U755 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U756 ( .A1(n873), .A2(n701), .ZN(n688) );
  NAND2_X1 U757 ( .A1(G1976), .A2(G288), .ZN(n872) );
  NAND2_X1 U758 ( .A1(n689), .A2(n872), .ZN(n690) );
  XNOR2_X1 U759 ( .A(n690), .B(KEYINPUT102), .ZN(n696) );
  XOR2_X1 U760 ( .A(G1981), .B(G305), .Z(n887) );
  INV_X1 U761 ( .A(n887), .ZN(n694) );
  NAND2_X1 U762 ( .A1(n691), .A2(KEYINPUT33), .ZN(n692) );
  NOR2_X1 U763 ( .A1(n692), .A2(n706), .ZN(n693) );
  OR2_X1 U764 ( .A1(n694), .A2(n693), .ZN(n697) );
  OR2_X1 U765 ( .A1(n706), .A2(n697), .ZN(n695) );
  OR2_X2 U766 ( .A1(n696), .A2(n695), .ZN(n753) );
  INV_X1 U767 ( .A(n697), .ZN(n698) );
  NOR2_X1 U768 ( .A1(G2090), .A2(G303), .ZN(n699) );
  NAND2_X1 U769 ( .A1(G8), .A2(n699), .ZN(n700) );
  NAND2_X1 U770 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U771 ( .A1(n702), .A2(n706), .ZN(n703) );
  XNOR2_X1 U772 ( .A(n703), .B(KEYINPUT103), .ZN(n708) );
  NOR2_X1 U773 ( .A1(G1981), .A2(G305), .ZN(n704) );
  XOR2_X1 U774 ( .A(n704), .B(KEYINPUT24), .Z(n705) );
  NOR2_X1 U775 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U776 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U777 ( .A1(n519), .A2(n709), .ZN(n751) );
  NAND2_X1 U778 ( .A1(n710), .A2(G129), .ZN(n711) );
  XNOR2_X1 U779 ( .A(n711), .B(KEYINPUT90), .ZN(n718) );
  NAND2_X1 U780 ( .A1(G117), .A2(n989), .ZN(n713) );
  NAND2_X1 U781 ( .A1(G141), .A2(n993), .ZN(n712) );
  NAND2_X1 U782 ( .A1(n713), .A2(n712), .ZN(n716) );
  NAND2_X1 U783 ( .A1(n992), .A2(G105), .ZN(n714) );
  XOR2_X1 U784 ( .A(KEYINPUT38), .B(n714), .Z(n715) );
  NOR2_X1 U785 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U786 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U787 ( .A(KEYINPUT91), .B(n719), .Z(n1002) );
  NOR2_X1 U788 ( .A1(G1996), .A2(n1002), .ZN(n937) );
  NOR2_X1 U789 ( .A1(n721), .A2(n720), .ZN(n756) );
  NAND2_X1 U790 ( .A1(G1996), .A2(n1002), .ZN(n729) );
  XOR2_X1 U791 ( .A(G1991), .B(KEYINPUT89), .Z(n852) );
  NAND2_X1 U792 ( .A1(G107), .A2(n989), .ZN(n723) );
  NAND2_X1 U793 ( .A1(G95), .A2(n992), .ZN(n722) );
  NAND2_X1 U794 ( .A1(n723), .A2(n722), .ZN(n727) );
  NAND2_X1 U795 ( .A1(G131), .A2(n993), .ZN(n725) );
  NAND2_X1 U796 ( .A1(G119), .A2(n710), .ZN(n724) );
  NAND2_X1 U797 ( .A1(n725), .A2(n724), .ZN(n726) );
  OR2_X1 U798 ( .A1(n727), .A2(n726), .ZN(n988) );
  NAND2_X1 U799 ( .A1(n852), .A2(n988), .ZN(n728) );
  NAND2_X1 U800 ( .A1(n729), .A2(n728), .ZN(n943) );
  NAND2_X1 U801 ( .A1(n756), .A2(n943), .ZN(n759) );
  INV_X1 U802 ( .A(n759), .ZN(n732) );
  NOR2_X1 U803 ( .A1(G1986), .A2(G290), .ZN(n730) );
  NOR2_X1 U804 ( .A1(n852), .A2(n988), .ZN(n939) );
  NOR2_X1 U805 ( .A1(n730), .A2(n939), .ZN(n731) );
  NOR2_X1 U806 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U807 ( .A1(n937), .A2(n733), .ZN(n734) );
  XNOR2_X1 U808 ( .A(n734), .B(KEYINPUT39), .ZN(n746) );
  XNOR2_X1 U809 ( .A(G2067), .B(KEYINPUT37), .ZN(n747) );
  NAND2_X1 U810 ( .A1(G116), .A2(n989), .ZN(n736) );
  NAND2_X1 U811 ( .A1(G128), .A2(n710), .ZN(n735) );
  NAND2_X1 U812 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U813 ( .A(n737), .B(KEYINPUT35), .ZN(n742) );
  NAND2_X1 U814 ( .A1(G104), .A2(n992), .ZN(n739) );
  NAND2_X1 U815 ( .A1(G140), .A2(n993), .ZN(n738) );
  NAND2_X1 U816 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U817 ( .A(KEYINPUT34), .B(n740), .Z(n741) );
  NAND2_X1 U818 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U819 ( .A(n743), .B(KEYINPUT36), .Z(n1011) );
  OR2_X1 U820 ( .A1(n747), .A2(n1011), .ZN(n744) );
  XNOR2_X1 U821 ( .A(n744), .B(KEYINPUT87), .ZN(n947) );
  NAND2_X1 U822 ( .A1(n947), .A2(n756), .ZN(n745) );
  XNOR2_X1 U823 ( .A(n745), .B(KEYINPUT88), .ZN(n760) );
  NAND2_X1 U824 ( .A1(n746), .A2(n760), .ZN(n748) );
  NAND2_X1 U825 ( .A1(n1011), .A2(n747), .ZN(n952) );
  NAND2_X1 U826 ( .A1(n748), .A2(n952), .ZN(n749) );
  XNOR2_X1 U827 ( .A(KEYINPUT104), .B(n749), .ZN(n750) );
  NAND2_X1 U828 ( .A1(n750), .A2(n756), .ZN(n754) );
  AND2_X1 U829 ( .A1(n751), .A2(n754), .ZN(n752) );
  NAND2_X1 U830 ( .A1(n753), .A2(n752), .ZN(n766) );
  INV_X1 U831 ( .A(n754), .ZN(n764) );
  XOR2_X1 U832 ( .A(G1986), .B(KEYINPUT85), .Z(n755) );
  XNOR2_X1 U833 ( .A(G290), .B(n755), .ZN(n882) );
  NAND2_X1 U834 ( .A1(n882), .A2(n756), .ZN(n757) );
  XNOR2_X1 U835 ( .A(KEYINPUT86), .B(n757), .ZN(n758) );
  NAND2_X1 U836 ( .A1(n759), .A2(n758), .ZN(n762) );
  INV_X1 U837 ( .A(n760), .ZN(n761) );
  NOR2_X1 U838 ( .A1(n762), .A2(n761), .ZN(n763) );
  OR2_X1 U839 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U840 ( .A(n768), .B(n767), .ZN(G329) );
  AND2_X1 U841 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U842 ( .A1(G111), .A2(n989), .ZN(n771) );
  NAND2_X1 U843 ( .A1(G99), .A2(n992), .ZN(n770) );
  NAND2_X1 U844 ( .A1(n771), .A2(n770), .ZN(n777) );
  NAND2_X1 U845 ( .A1(n710), .A2(G123), .ZN(n772) );
  XNOR2_X1 U846 ( .A(n772), .B(KEYINPUT18), .ZN(n773) );
  XNOR2_X1 U847 ( .A(n773), .B(KEYINPUT74), .ZN(n775) );
  NAND2_X1 U848 ( .A1(G135), .A2(n993), .ZN(n774) );
  NAND2_X1 U849 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U850 ( .A1(n777), .A2(n776), .ZN(n985) );
  XNOR2_X1 U851 ( .A(n985), .B(G2096), .ZN(n778) );
  XNOR2_X1 U852 ( .A(n778), .B(KEYINPUT75), .ZN(n779) );
  OR2_X1 U853 ( .A1(G2100), .A2(n779), .ZN(G156) );
  INV_X1 U854 ( .A(G860), .ZN(n787) );
  OR2_X1 U855 ( .A1(n787), .A2(n880), .ZN(G153) );
  INV_X1 U856 ( .A(G57), .ZN(G237) );
  INV_X1 U857 ( .A(G132), .ZN(G219) );
  INV_X1 U858 ( .A(G82), .ZN(G220) );
  XOR2_X1 U859 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n781) );
  NAND2_X1 U860 ( .A1(G7), .A2(G661), .ZN(n780) );
  XOR2_X1 U861 ( .A(n781), .B(n780), .Z(n834) );
  NAND2_X1 U862 ( .A1(n834), .A2(G567), .ZN(n782) );
  XOR2_X1 U863 ( .A(KEYINPUT11), .B(n782), .Z(G234) );
  NAND2_X1 U864 ( .A1(G868), .A2(G301), .ZN(n784) );
  INV_X1 U865 ( .A(G868), .ZN(n819) );
  NAND2_X1 U866 ( .A1(n1015), .A2(n819), .ZN(n783) );
  NAND2_X1 U867 ( .A1(n784), .A2(n783), .ZN(G284) );
  NOR2_X1 U868 ( .A1(G286), .A2(n819), .ZN(n786) );
  NOR2_X1 U869 ( .A1(G868), .A2(G299), .ZN(n785) );
  NOR2_X1 U870 ( .A1(n786), .A2(n785), .ZN(G297) );
  NAND2_X1 U871 ( .A1(n787), .A2(G559), .ZN(n788) );
  NAND2_X1 U872 ( .A1(n788), .A2(n869), .ZN(n789) );
  XNOR2_X1 U873 ( .A(n789), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U874 ( .A1(n880), .A2(G868), .ZN(n792) );
  NAND2_X1 U875 ( .A1(G868), .A2(n869), .ZN(n790) );
  NOR2_X1 U876 ( .A1(G559), .A2(n790), .ZN(n791) );
  NOR2_X1 U877 ( .A1(n792), .A2(n791), .ZN(G282) );
  NAND2_X1 U878 ( .A1(G559), .A2(n869), .ZN(n793) );
  XNOR2_X1 U879 ( .A(n793), .B(KEYINPUT76), .ZN(n816) );
  XNOR2_X1 U880 ( .A(n880), .B(n816), .ZN(n794) );
  NOR2_X1 U881 ( .A1(G860), .A2(n794), .ZN(n795) );
  XNOR2_X1 U882 ( .A(n795), .B(KEYINPUT77), .ZN(n808) );
  NAND2_X1 U883 ( .A1(n796), .A2(G80), .ZN(n797) );
  XNOR2_X1 U884 ( .A(n797), .B(KEYINPUT78), .ZN(n800) );
  NAND2_X1 U885 ( .A1(G93), .A2(n798), .ZN(n799) );
  NAND2_X1 U886 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U887 ( .A(KEYINPUT79), .B(n801), .ZN(n807) );
  NAND2_X1 U888 ( .A1(G55), .A2(n802), .ZN(n805) );
  NAND2_X1 U889 ( .A1(G67), .A2(n803), .ZN(n804) );
  AND2_X1 U890 ( .A1(n805), .A2(n804), .ZN(n806) );
  NAND2_X1 U891 ( .A1(n807), .A2(n806), .ZN(n818) );
  XNOR2_X1 U892 ( .A(n808), .B(n818), .ZN(G145) );
  XOR2_X1 U893 ( .A(G290), .B(G305), .Z(n809) );
  XNOR2_X1 U894 ( .A(G288), .B(n809), .ZN(n810) );
  XOR2_X1 U895 ( .A(n810), .B(KEYINPUT19), .Z(n812) );
  XOR2_X1 U896 ( .A(n818), .B(KEYINPUT83), .Z(n811) );
  XNOR2_X1 U897 ( .A(n812), .B(n811), .ZN(n813) );
  XNOR2_X1 U898 ( .A(G299), .B(n813), .ZN(n815) );
  XOR2_X1 U899 ( .A(G303), .B(n880), .Z(n814) );
  XNOR2_X1 U900 ( .A(n815), .B(n814), .ZN(n1014) );
  XNOR2_X1 U901 ( .A(n816), .B(n1014), .ZN(n817) );
  NAND2_X1 U902 ( .A1(n817), .A2(G868), .ZN(n821) );
  NAND2_X1 U903 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U904 ( .A1(n821), .A2(n820), .ZN(G295) );
  NAND2_X1 U905 ( .A1(G2078), .A2(G2084), .ZN(n822) );
  XOR2_X1 U906 ( .A(KEYINPUT20), .B(n822), .Z(n823) );
  NAND2_X1 U907 ( .A1(G2090), .A2(n823), .ZN(n824) );
  XNOR2_X1 U908 ( .A(KEYINPUT21), .B(n824), .ZN(n825) );
  NAND2_X1 U909 ( .A1(n825), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U910 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U911 ( .A1(G220), .A2(G219), .ZN(n826) );
  XOR2_X1 U912 ( .A(KEYINPUT22), .B(n826), .Z(n827) );
  NOR2_X1 U913 ( .A1(G218), .A2(n827), .ZN(n828) );
  NAND2_X1 U914 ( .A1(G96), .A2(n828), .ZN(n961) );
  NAND2_X1 U915 ( .A1(n961), .A2(G2106), .ZN(n832) );
  NAND2_X1 U916 ( .A1(G120), .A2(G69), .ZN(n829) );
  NOR2_X1 U917 ( .A1(G237), .A2(n829), .ZN(n830) );
  NAND2_X1 U918 ( .A1(G108), .A2(n830), .ZN(n962) );
  NAND2_X1 U919 ( .A1(n962), .A2(G567), .ZN(n831) );
  NAND2_X1 U920 ( .A1(n832), .A2(n831), .ZN(n963) );
  NAND2_X1 U921 ( .A1(G483), .A2(G661), .ZN(n833) );
  NOR2_X1 U922 ( .A1(n963), .A2(n833), .ZN(n838) );
  NAND2_X1 U923 ( .A1(n838), .A2(G36), .ZN(G176) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n834), .ZN(G217) );
  INV_X1 U925 ( .A(n834), .ZN(G223) );
  AND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U927 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n836) );
  XOR2_X1 U929 ( .A(KEYINPUT107), .B(n836), .Z(n837) );
  NAND2_X1 U930 ( .A1(n838), .A2(n837), .ZN(G188) );
  XOR2_X1 U931 ( .A(G69), .B(KEYINPUT108), .Z(G235) );
  NAND2_X1 U933 ( .A1(G112), .A2(n989), .ZN(n840) );
  NAND2_X1 U934 ( .A1(G100), .A2(n992), .ZN(n839) );
  NAND2_X1 U935 ( .A1(n840), .A2(n839), .ZN(n846) );
  NAND2_X1 U936 ( .A1(n710), .A2(G124), .ZN(n841) );
  XNOR2_X1 U937 ( .A(n841), .B(KEYINPUT44), .ZN(n844) );
  NAND2_X1 U938 ( .A1(G136), .A2(n993), .ZN(n842) );
  XOR2_X1 U939 ( .A(KEYINPUT111), .B(n842), .Z(n843) );
  NAND2_X1 U940 ( .A1(n844), .A2(n843), .ZN(n845) );
  NOR2_X1 U941 ( .A1(n846), .A2(n845), .ZN(G162) );
  XOR2_X1 U942 ( .A(G2090), .B(G35), .Z(n862) );
  XOR2_X1 U943 ( .A(G2072), .B(G33), .Z(n847) );
  NAND2_X1 U944 ( .A1(n847), .A2(G28), .ZN(n858) );
  XNOR2_X1 U945 ( .A(G27), .B(n848), .ZN(n849) );
  XNOR2_X1 U946 ( .A(n849), .B(KEYINPUT117), .ZN(n856) );
  XOR2_X1 U947 ( .A(G2067), .B(G26), .Z(n851) );
  XOR2_X1 U948 ( .A(G1996), .B(G32), .Z(n850) );
  NAND2_X1 U949 ( .A1(n851), .A2(n850), .ZN(n854) );
  XNOR2_X1 U950 ( .A(G25), .B(n852), .ZN(n853) );
  NOR2_X1 U951 ( .A1(n854), .A2(n853), .ZN(n855) );
  NAND2_X1 U952 ( .A1(n856), .A2(n855), .ZN(n857) );
  NOR2_X1 U953 ( .A1(n858), .A2(n857), .ZN(n859) );
  XOR2_X1 U954 ( .A(KEYINPUT53), .B(n859), .Z(n860) );
  XNOR2_X1 U955 ( .A(n860), .B(KEYINPUT118), .ZN(n861) );
  NAND2_X1 U956 ( .A1(n862), .A2(n861), .ZN(n865) );
  XNOR2_X1 U957 ( .A(KEYINPUT54), .B(G2084), .ZN(n863) );
  XNOR2_X1 U958 ( .A(G34), .B(n863), .ZN(n864) );
  NOR2_X1 U959 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U960 ( .A(KEYINPUT55), .B(n866), .ZN(n867) );
  XNOR2_X1 U961 ( .A(KEYINPUT119), .B(n867), .ZN(n868) );
  NOR2_X1 U962 ( .A1(G29), .A2(n868), .ZN(n923) );
  INV_X1 U963 ( .A(G16), .ZN(n919) );
  XOR2_X1 U964 ( .A(n919), .B(KEYINPUT56), .Z(n895) );
  XOR2_X1 U965 ( .A(n869), .B(G1348), .Z(n871) );
  XOR2_X1 U966 ( .A(G171), .B(G1961), .Z(n870) );
  NOR2_X1 U967 ( .A1(n871), .A2(n870), .ZN(n893) );
  XOR2_X1 U968 ( .A(G299), .B(G1956), .Z(n878) );
  INV_X1 U969 ( .A(G1971), .ZN(n974) );
  NOR2_X1 U970 ( .A1(G166), .A2(n974), .ZN(n875) );
  NAND2_X1 U971 ( .A1(n873), .A2(n872), .ZN(n874) );
  NOR2_X1 U972 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U973 ( .A(KEYINPUT122), .B(n876), .ZN(n877) );
  NAND2_X1 U974 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U975 ( .A(KEYINPUT123), .B(n879), .ZN(n884) );
  XNOR2_X1 U976 ( .A(G1341), .B(n880), .ZN(n881) );
  NOR2_X1 U977 ( .A1(n882), .A2(n881), .ZN(n883) );
  NAND2_X1 U978 ( .A1(n884), .A2(n883), .ZN(n891) );
  XOR2_X1 U979 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n889) );
  XNOR2_X1 U980 ( .A(G1966), .B(G168), .ZN(n885) );
  XNOR2_X1 U981 ( .A(n885), .B(KEYINPUT120), .ZN(n886) );
  NAND2_X1 U982 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U983 ( .A(n889), .B(n888), .Z(n890) );
  NOR2_X1 U984 ( .A1(n891), .A2(n890), .ZN(n892) );
  NAND2_X1 U985 ( .A1(n893), .A2(n892), .ZN(n894) );
  NAND2_X1 U986 ( .A1(n895), .A2(n894), .ZN(n921) );
  XOR2_X1 U987 ( .A(G1348), .B(KEYINPUT59), .Z(n896) );
  XNOR2_X1 U988 ( .A(G4), .B(n896), .ZN(n904) );
  XNOR2_X1 U989 ( .A(G1981), .B(G6), .ZN(n898) );
  XNOR2_X1 U990 ( .A(G19), .B(G1341), .ZN(n897) );
  NOR2_X1 U991 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U992 ( .A(KEYINPUT124), .B(n899), .Z(n901) );
  XNOR2_X1 U993 ( .A(G1956), .B(G20), .ZN(n900) );
  NOR2_X1 U994 ( .A1(n901), .A2(n900), .ZN(n902) );
  XNOR2_X1 U995 ( .A(n902), .B(KEYINPUT125), .ZN(n903) );
  NOR2_X1 U996 ( .A1(n904), .A2(n903), .ZN(n905) );
  XNOR2_X1 U997 ( .A(KEYINPUT60), .B(n905), .ZN(n909) );
  XNOR2_X1 U998 ( .A(G1966), .B(G21), .ZN(n907) );
  XNOR2_X1 U999 ( .A(G5), .B(G1961), .ZN(n906) );
  NOR2_X1 U1000 ( .A1(n907), .A2(n906), .ZN(n908) );
  NAND2_X1 U1001 ( .A1(n909), .A2(n908), .ZN(n916) );
  XNOR2_X1 U1002 ( .A(G1976), .B(G23), .ZN(n911) );
  XOR2_X1 U1003 ( .A(n974), .B(G22), .Z(n910) );
  NOR2_X1 U1004 ( .A1(n911), .A2(n910), .ZN(n913) );
  XOR2_X1 U1005 ( .A(G1986), .B(G24), .Z(n912) );
  NAND2_X1 U1006 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1007 ( .A(KEYINPUT58), .B(n914), .ZN(n915) );
  NOR2_X1 U1008 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1009 ( .A(KEYINPUT61), .B(n917), .ZN(n918) );
  NAND2_X1 U1010 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1011 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1012 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1013 ( .A1(G11), .A2(n924), .ZN(n925) );
  XNOR2_X1 U1014 ( .A(n925), .B(KEYINPUT126), .ZN(n959) );
  INV_X1 U1015 ( .A(G29), .ZN(n957) );
  NAND2_X1 U1016 ( .A1(G103), .A2(n992), .ZN(n927) );
  NAND2_X1 U1017 ( .A1(G139), .A2(n993), .ZN(n926) );
  NAND2_X1 U1018 ( .A1(n927), .A2(n926), .ZN(n932) );
  NAND2_X1 U1019 ( .A1(G115), .A2(n989), .ZN(n929) );
  NAND2_X1 U1020 ( .A1(G127), .A2(n710), .ZN(n928) );
  NAND2_X1 U1021 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1022 ( .A(KEYINPUT47), .B(n930), .Z(n931) );
  NOR2_X1 U1023 ( .A1(n932), .A2(n931), .ZN(n986) );
  XOR2_X1 U1024 ( .A(G2072), .B(n986), .Z(n934) );
  XOR2_X1 U1025 ( .A(G164), .B(G2078), .Z(n933) );
  NOR2_X1 U1026 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1027 ( .A(KEYINPUT50), .B(n935), .Z(n950) );
  XOR2_X1 U1028 ( .A(G2090), .B(G162), .Z(n936) );
  NOR2_X1 U1029 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1030 ( .A(KEYINPUT51), .B(n938), .Z(n945) );
  XNOR2_X1 U1031 ( .A(G160), .B(G2084), .ZN(n941) );
  NOR2_X1 U1032 ( .A1(n939), .A2(n985), .ZN(n940) );
  NAND2_X1 U1033 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1034 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1035 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1036 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1037 ( .A(KEYINPUT115), .B(n948), .ZN(n949) );
  NOR2_X1 U1038 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1039 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1040 ( .A(n953), .B(KEYINPUT52), .ZN(n954) );
  XNOR2_X1 U1041 ( .A(n954), .B(KEYINPUT116), .ZN(n955) );
  NOR2_X1 U1042 ( .A1(KEYINPUT55), .A2(n955), .ZN(n956) );
  NOR2_X1 U1043 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1044 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1045 ( .A(KEYINPUT62), .B(n960), .ZN(G311) );
  XNOR2_X1 U1046 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1047 ( .A(G120), .ZN(G236) );
  INV_X1 U1048 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1049 ( .A1(n962), .A2(n961), .ZN(G325) );
  INV_X1 U1050 ( .A(G325), .ZN(G261) );
  INV_X1 U1051 ( .A(n963), .ZN(G319) );
  XOR2_X1 U1052 ( .A(G2678), .B(KEYINPUT43), .Z(n965) );
  XNOR2_X1 U1053 ( .A(G2072), .B(G2090), .ZN(n964) );
  XNOR2_X1 U1054 ( .A(n965), .B(n964), .ZN(n969) );
  XOR2_X1 U1055 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n967) );
  XNOR2_X1 U1056 ( .A(G2067), .B(KEYINPUT110), .ZN(n966) );
  XNOR2_X1 U1057 ( .A(n967), .B(n966), .ZN(n968) );
  XOR2_X1 U1058 ( .A(n969), .B(n968), .Z(n971) );
  XNOR2_X1 U1059 ( .A(G2096), .B(G2100), .ZN(n970) );
  XNOR2_X1 U1060 ( .A(n971), .B(n970), .ZN(n973) );
  XOR2_X1 U1061 ( .A(G2078), .B(G2084), .Z(n972) );
  XNOR2_X1 U1062 ( .A(n973), .B(n972), .ZN(G227) );
  XOR2_X1 U1063 ( .A(G1961), .B(G1956), .Z(n976) );
  XOR2_X1 U1064 ( .A(G1986), .B(n974), .Z(n975) );
  XNOR2_X1 U1065 ( .A(n976), .B(n975), .ZN(n977) );
  XOR2_X1 U1066 ( .A(n977), .B(KEYINPUT41), .Z(n980) );
  XOR2_X1 U1067 ( .A(n978), .B(G1966), .Z(n979) );
  XNOR2_X1 U1068 ( .A(n980), .B(n979), .ZN(n984) );
  XOR2_X1 U1069 ( .A(G2474), .B(G1976), .Z(n982) );
  XNOR2_X1 U1070 ( .A(G1991), .B(G1981), .ZN(n981) );
  XNOR2_X1 U1071 ( .A(n982), .B(n981), .ZN(n983) );
  XNOR2_X1 U1072 ( .A(n984), .B(n983), .ZN(G229) );
  XOR2_X1 U1073 ( .A(n986), .B(n985), .Z(n987) );
  XNOR2_X1 U1074 ( .A(n988), .B(n987), .ZN(n1001) );
  NAND2_X1 U1075 ( .A1(G118), .A2(n989), .ZN(n991) );
  NAND2_X1 U1076 ( .A1(G130), .A2(n710), .ZN(n990) );
  NAND2_X1 U1077 ( .A1(n991), .A2(n990), .ZN(n999) );
  NAND2_X1 U1078 ( .A1(G106), .A2(n992), .ZN(n995) );
  NAND2_X1 U1079 ( .A1(G142), .A2(n993), .ZN(n994) );
  NAND2_X1 U1080 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1081 ( .A(KEYINPUT112), .B(n996), .Z(n997) );
  XNOR2_X1 U1082 ( .A(KEYINPUT45), .B(n997), .ZN(n998) );
  NOR2_X1 U1083 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1084 ( .A(n1001), .B(n1000), .ZN(n1004) );
  XNOR2_X1 U1085 ( .A(n1002), .B(G162), .ZN(n1003) );
  XNOR2_X1 U1086 ( .A(n1004), .B(n1003), .ZN(n1008) );
  XOR2_X1 U1087 ( .A(KEYINPUT46), .B(KEYINPUT113), .Z(n1006) );
  XNOR2_X1 U1088 ( .A(KEYINPUT114), .B(KEYINPUT48), .ZN(n1005) );
  XNOR2_X1 U1089 ( .A(n1006), .B(n1005), .ZN(n1007) );
  XOR2_X1 U1090 ( .A(n1008), .B(n1007), .Z(n1010) );
  XNOR2_X1 U1091 ( .A(G164), .B(G160), .ZN(n1009) );
  XNOR2_X1 U1092 ( .A(n1010), .B(n1009), .ZN(n1012) );
  XNOR2_X1 U1093 ( .A(n1012), .B(n1011), .ZN(n1013) );
  NOR2_X1 U1094 ( .A1(G37), .A2(n1013), .ZN(G395) );
  XOR2_X1 U1095 ( .A(n1014), .B(G286), .Z(n1017) );
  XOR2_X1 U1096 ( .A(n1015), .B(G171), .Z(n1016) );
  XNOR2_X1 U1097 ( .A(n1017), .B(n1016), .ZN(n1018) );
  NOR2_X1 U1098 ( .A1(G37), .A2(n1018), .ZN(G397) );
  XNOR2_X1 U1099 ( .A(G1348), .B(G2446), .ZN(n1028) );
  XOR2_X1 U1100 ( .A(G2435), .B(G2454), .Z(n1020) );
  XNOR2_X1 U1101 ( .A(G1341), .B(G2430), .ZN(n1019) );
  XNOR2_X1 U1102 ( .A(n1020), .B(n1019), .ZN(n1024) );
  XOR2_X1 U1103 ( .A(G2443), .B(G2451), .Z(n1022) );
  XNOR2_X1 U1104 ( .A(KEYINPUT105), .B(G2427), .ZN(n1021) );
  XNOR2_X1 U1105 ( .A(n1022), .B(n1021), .ZN(n1023) );
  XOR2_X1 U1106 ( .A(n1024), .B(n1023), .Z(n1026) );
  XNOR2_X1 U1107 ( .A(KEYINPUT106), .B(G2438), .ZN(n1025) );
  XNOR2_X1 U1108 ( .A(n1026), .B(n1025), .ZN(n1027) );
  XNOR2_X1 U1109 ( .A(n1028), .B(n1027), .ZN(n1029) );
  NAND2_X1 U1110 ( .A1(n1029), .A2(G14), .ZN(n1035) );
  NAND2_X1 U1111 ( .A1(G319), .A2(n1035), .ZN(n1032) );
  NOR2_X1 U1112 ( .A1(G227), .A2(G229), .ZN(n1030) );
  XNOR2_X1 U1113 ( .A(KEYINPUT49), .B(n1030), .ZN(n1031) );
  NOR2_X1 U1114 ( .A1(n1032), .A2(n1031), .ZN(n1034) );
  NOR2_X1 U1115 ( .A1(G395), .A2(G397), .ZN(n1033) );
  NAND2_X1 U1116 ( .A1(n1034), .A2(n1033), .ZN(G225) );
  INV_X1 U1117 ( .A(G225), .ZN(G308) );
  INV_X1 U1118 ( .A(G108), .ZN(G238) );
  INV_X1 U1119 ( .A(n1035), .ZN(G401) );
endmodule

