

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U557 ( .A1(n698), .A2(n764), .ZN(n738) );
  AND2_X1 U558 ( .A1(n539), .A2(G2104), .ZN(n893) );
  XOR2_X1 U559 ( .A(n718), .B(KEYINPUT28), .Z(n523) );
  XNOR2_X1 U560 ( .A(n721), .B(n720), .ZN(n726) );
  NOR2_X1 U561 ( .A1(G651), .A2(n650), .ZN(n649) );
  NOR2_X1 U562 ( .A1(n816), .A2(n815), .ZN(n524) );
  NAND2_X1 U563 ( .A1(n819), .A2(n818), .ZN(n525) );
  XOR2_X1 U564 ( .A(n760), .B(KEYINPUT64), .Z(n526) );
  NOR2_X1 U565 ( .A1(n698), .A2(n764), .ZN(n722) );
  INV_X1 U566 ( .A(KEYINPUT29), .ZN(n720) );
  NOR2_X1 U567 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U568 ( .A1(G8), .A2(n738), .ZN(n810) );
  NOR2_X1 U569 ( .A1(n539), .A2(G2104), .ZN(n540) );
  INV_X1 U570 ( .A(KEYINPUT93), .ZN(n541) );
  XNOR2_X1 U571 ( .A(n540), .B(KEYINPUT66), .ZN(n688) );
  XNOR2_X1 U572 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U573 ( .A(KEYINPUT1), .B(n528), .Z(n654) );
  XOR2_X1 U574 ( .A(G543), .B(KEYINPUT0), .Z(n527) );
  XNOR2_X1 U575 ( .A(KEYINPUT68), .B(n527), .ZN(n650) );
  NAND2_X1 U576 ( .A1(n649), .A2(G52), .ZN(n530) );
  XNOR2_X1 U577 ( .A(KEYINPUT69), .B(G651), .ZN(n531) );
  NOR2_X1 U578 ( .A1(G543), .A2(n531), .ZN(n528) );
  NAND2_X1 U579 ( .A1(G64), .A2(n654), .ZN(n529) );
  NAND2_X1 U580 ( .A1(n530), .A2(n529), .ZN(n537) );
  NOR2_X1 U581 ( .A1(G543), .A2(G651), .ZN(n640) );
  NAND2_X1 U582 ( .A1(G90), .A2(n640), .ZN(n533) );
  NOR2_X1 U583 ( .A1(n650), .A2(n531), .ZN(n643) );
  NAND2_X1 U584 ( .A1(G77), .A2(n643), .ZN(n532) );
  NAND2_X1 U585 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U586 ( .A(KEYINPUT72), .B(n534), .Z(n535) );
  XNOR2_X1 U587 ( .A(KEYINPUT9), .B(n535), .ZN(n536) );
  NOR2_X1 U588 ( .A1(n537), .A2(n536), .ZN(G171) );
  AND2_X1 U589 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U590 ( .A(G57), .ZN(G237) );
  INV_X1 U591 ( .A(G2105), .ZN(n539) );
  NAND2_X1 U592 ( .A1(G102), .A2(n893), .ZN(n538) );
  XNOR2_X1 U593 ( .A(n538), .B(KEYINPUT94), .ZN(n544) );
  NAND2_X1 U594 ( .A1(n688), .A2(G126), .ZN(n542) );
  NAND2_X1 U595 ( .A1(n544), .A2(n543), .ZN(n549) );
  NOR2_X1 U596 ( .A1(G2105), .A2(G2104), .ZN(n545) );
  XOR2_X1 U597 ( .A(KEYINPUT17), .B(n545), .Z(n607) );
  NAND2_X1 U598 ( .A1(n607), .A2(G138), .ZN(n547) );
  AND2_X1 U599 ( .A1(G2105), .A2(G2104), .ZN(n901) );
  NAND2_X1 U600 ( .A1(n901), .A2(G114), .ZN(n546) );
  NAND2_X1 U601 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U602 ( .A1(n549), .A2(n548), .ZN(n696) );
  BUF_X1 U603 ( .A(n696), .Z(G164) );
  NAND2_X1 U604 ( .A1(n640), .A2(G89), .ZN(n550) );
  XNOR2_X1 U605 ( .A(n550), .B(KEYINPUT4), .ZN(n552) );
  NAND2_X1 U606 ( .A1(G76), .A2(n643), .ZN(n551) );
  NAND2_X1 U607 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U608 ( .A(n553), .B(KEYINPUT5), .ZN(n560) );
  XNOR2_X1 U609 ( .A(KEYINPUT6), .B(KEYINPUT77), .ZN(n558) );
  NAND2_X1 U610 ( .A1(n649), .A2(G51), .ZN(n554) );
  XNOR2_X1 U611 ( .A(n554), .B(KEYINPUT76), .ZN(n556) );
  NAND2_X1 U612 ( .A1(G63), .A2(n654), .ZN(n555) );
  NAND2_X1 U613 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U614 ( .A(n558), .B(n557), .ZN(n559) );
  NAND2_X1 U615 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U616 ( .A(KEYINPUT7), .B(n561), .ZN(G168) );
  XOR2_X1 U617 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U618 ( .A1(G7), .A2(G661), .ZN(n562) );
  XNOR2_X1 U619 ( .A(n562), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U620 ( .A(G223), .ZN(n841) );
  NAND2_X1 U621 ( .A1(n841), .A2(G567), .ZN(n563) );
  XOR2_X1 U622 ( .A(KEYINPUT11), .B(n563), .Z(G234) );
  NAND2_X1 U623 ( .A1(n640), .A2(G81), .ZN(n564) );
  XNOR2_X1 U624 ( .A(n564), .B(KEYINPUT12), .ZN(n566) );
  NAND2_X1 U625 ( .A1(G68), .A2(n643), .ZN(n565) );
  NAND2_X1 U626 ( .A1(n566), .A2(n565), .ZN(n568) );
  XOR2_X1 U627 ( .A(KEYINPUT74), .B(KEYINPUT13), .Z(n567) );
  XNOR2_X1 U628 ( .A(n568), .B(n567), .ZN(n571) );
  NAND2_X1 U629 ( .A1(G56), .A2(n654), .ZN(n569) );
  XOR2_X1 U630 ( .A(KEYINPUT14), .B(n569), .Z(n570) );
  NOR2_X1 U631 ( .A1(n571), .A2(n570), .ZN(n573) );
  NAND2_X1 U632 ( .A1(n649), .A2(G43), .ZN(n572) );
  NAND2_X1 U633 ( .A1(n573), .A2(n572), .ZN(n981) );
  INV_X1 U634 ( .A(G860), .ZN(n594) );
  OR2_X1 U635 ( .A1(n981), .A2(n594), .ZN(G153) );
  XNOR2_X1 U636 ( .A(G171), .B(KEYINPUT75), .ZN(G301) );
  NAND2_X1 U637 ( .A1(G868), .A2(G301), .ZN(n582) );
  NAND2_X1 U638 ( .A1(n649), .A2(G54), .ZN(n575) );
  NAND2_X1 U639 ( .A1(G66), .A2(n654), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n579) );
  NAND2_X1 U641 ( .A1(G92), .A2(n640), .ZN(n577) );
  NAND2_X1 U642 ( .A1(G79), .A2(n643), .ZN(n576) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(KEYINPUT15), .ZN(n988) );
  INV_X1 U646 ( .A(G868), .ZN(n668) );
  NAND2_X1 U647 ( .A1(n988), .A2(n668), .ZN(n581) );
  NAND2_X1 U648 ( .A1(n582), .A2(n581), .ZN(G284) );
  NAND2_X1 U649 ( .A1(G65), .A2(n654), .ZN(n584) );
  NAND2_X1 U650 ( .A1(G78), .A2(n643), .ZN(n583) );
  NAND2_X1 U651 ( .A1(n584), .A2(n583), .ZN(n587) );
  NAND2_X1 U652 ( .A1(G91), .A2(n640), .ZN(n585) );
  XNOR2_X1 U653 ( .A(KEYINPUT73), .B(n585), .ZN(n586) );
  NOR2_X1 U654 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U655 ( .A1(n649), .A2(G53), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n589), .A2(n588), .ZN(G299) );
  NOR2_X1 U657 ( .A1(G286), .A2(n668), .ZN(n590) );
  XNOR2_X1 U658 ( .A(n590), .B(KEYINPUT78), .ZN(n592) );
  NOR2_X1 U659 ( .A1(G299), .A2(G868), .ZN(n591) );
  NOR2_X1 U660 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U661 ( .A(KEYINPUT79), .B(n593), .Z(G297) );
  NAND2_X1 U662 ( .A1(n594), .A2(G559), .ZN(n595) );
  INV_X1 U663 ( .A(n988), .ZN(n615) );
  NAND2_X1 U664 ( .A1(n595), .A2(n615), .ZN(n596) );
  XNOR2_X1 U665 ( .A(n596), .B(KEYINPUT80), .ZN(n597) );
  XNOR2_X1 U666 ( .A(KEYINPUT16), .B(n597), .ZN(G148) );
  NOR2_X1 U667 ( .A1(G868), .A2(n981), .ZN(n598) );
  XOR2_X1 U668 ( .A(KEYINPUT81), .B(n598), .Z(n601) );
  NAND2_X1 U669 ( .A1(G868), .A2(n615), .ZN(n599) );
  NOR2_X1 U670 ( .A1(G559), .A2(n599), .ZN(n600) );
  NOR2_X1 U671 ( .A1(n601), .A2(n600), .ZN(G282) );
  NAND2_X1 U672 ( .A1(G99), .A2(n893), .ZN(n603) );
  NAND2_X1 U673 ( .A1(G111), .A2(n901), .ZN(n602) );
  NAND2_X1 U674 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U675 ( .A(KEYINPUT83), .B(n604), .ZN(n612) );
  INV_X1 U676 ( .A(n688), .ZN(n605) );
  INV_X1 U677 ( .A(n605), .ZN(n898) );
  NAND2_X1 U678 ( .A1(G123), .A2(n898), .ZN(n606) );
  XNOR2_X1 U679 ( .A(n606), .B(KEYINPUT18), .ZN(n609) );
  BUF_X1 U680 ( .A(n607), .Z(n894) );
  NAND2_X1 U681 ( .A1(G135), .A2(n894), .ZN(n608) );
  NAND2_X1 U682 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U683 ( .A(KEYINPUT82), .B(n610), .Z(n611) );
  NAND2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n935) );
  XNOR2_X1 U685 ( .A(G2096), .B(n935), .ZN(n613) );
  NOR2_X1 U686 ( .A1(G2100), .A2(n613), .ZN(n614) );
  XOR2_X1 U687 ( .A(KEYINPUT84), .B(n614), .Z(G156) );
  NAND2_X1 U688 ( .A1(n615), .A2(G559), .ZN(n666) );
  XNOR2_X1 U689 ( .A(n981), .B(n666), .ZN(n616) );
  NOR2_X1 U690 ( .A1(n616), .A2(G860), .ZN(n623) );
  NAND2_X1 U691 ( .A1(G93), .A2(n640), .ZN(n618) );
  NAND2_X1 U692 ( .A1(G80), .A2(n643), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U694 ( .A1(n649), .A2(G55), .ZN(n620) );
  NAND2_X1 U695 ( .A1(G67), .A2(n654), .ZN(n619) );
  NAND2_X1 U696 ( .A1(n620), .A2(n619), .ZN(n621) );
  OR2_X1 U697 ( .A1(n622), .A2(n621), .ZN(n669) );
  XOR2_X1 U698 ( .A(n623), .B(n669), .Z(G145) );
  NAND2_X1 U699 ( .A1(G50), .A2(n649), .ZN(n624) );
  XOR2_X1 U700 ( .A(KEYINPUT86), .B(n624), .Z(n629) );
  NAND2_X1 U701 ( .A1(G88), .A2(n640), .ZN(n626) );
  NAND2_X1 U702 ( .A1(G75), .A2(n643), .ZN(n625) );
  NAND2_X1 U703 ( .A1(n626), .A2(n625), .ZN(n627) );
  XOR2_X1 U704 ( .A(KEYINPUT87), .B(n627), .Z(n628) );
  NOR2_X1 U705 ( .A1(n629), .A2(n628), .ZN(n631) );
  NAND2_X1 U706 ( .A1(G62), .A2(n654), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n631), .A2(n630), .ZN(G303) );
  INV_X1 U708 ( .A(G303), .ZN(G166) );
  NAND2_X1 U709 ( .A1(G60), .A2(n654), .ZN(n632) );
  XNOR2_X1 U710 ( .A(n632), .B(KEYINPUT70), .ZN(n634) );
  NAND2_X1 U711 ( .A1(G85), .A2(n640), .ZN(n633) );
  NAND2_X1 U712 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U713 ( .A1(n649), .A2(G47), .ZN(n636) );
  NAND2_X1 U714 ( .A1(G72), .A2(n643), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U716 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U717 ( .A(KEYINPUT71), .B(n639), .ZN(G290) );
  NAND2_X1 U718 ( .A1(G86), .A2(n640), .ZN(n642) );
  NAND2_X1 U719 ( .A1(G48), .A2(n649), .ZN(n641) );
  NAND2_X1 U720 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U721 ( .A1(n643), .A2(G73), .ZN(n644) );
  XOR2_X1 U722 ( .A(KEYINPUT2), .B(n644), .Z(n645) );
  NOR2_X1 U723 ( .A1(n646), .A2(n645), .ZN(n648) );
  NAND2_X1 U724 ( .A1(G61), .A2(n654), .ZN(n647) );
  NAND2_X1 U725 ( .A1(n648), .A2(n647), .ZN(G305) );
  NAND2_X1 U726 ( .A1(G49), .A2(n649), .ZN(n652) );
  NAND2_X1 U727 ( .A1(G87), .A2(n650), .ZN(n651) );
  NAND2_X1 U728 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U729 ( .A1(n654), .A2(n653), .ZN(n657) );
  NAND2_X1 U730 ( .A1(G74), .A2(G651), .ZN(n655) );
  XOR2_X1 U731 ( .A(KEYINPUT85), .B(n655), .Z(n656) );
  NAND2_X1 U732 ( .A1(n657), .A2(n656), .ZN(G288) );
  INV_X1 U733 ( .A(G299), .ZN(n716) );
  XNOR2_X1 U734 ( .A(n716), .B(G290), .ZN(n658) );
  XOR2_X1 U735 ( .A(n669), .B(n658), .Z(n663) );
  XNOR2_X1 U736 ( .A(KEYINPUT89), .B(KEYINPUT19), .ZN(n660) );
  XNOR2_X1 U737 ( .A(G288), .B(KEYINPUT88), .ZN(n659) );
  XNOR2_X1 U738 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U739 ( .A(G305), .B(n661), .ZN(n662) );
  XNOR2_X1 U740 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U741 ( .A(G166), .B(n664), .ZN(n665) );
  XNOR2_X1 U742 ( .A(n665), .B(n981), .ZN(n911) );
  XOR2_X1 U743 ( .A(n911), .B(n666), .Z(n667) );
  NOR2_X1 U744 ( .A1(n668), .A2(n667), .ZN(n671) );
  NOR2_X1 U745 ( .A1(G868), .A2(n669), .ZN(n670) );
  NOR2_X1 U746 ( .A1(n671), .A2(n670), .ZN(G295) );
  NAND2_X1 U747 ( .A1(G2078), .A2(G2084), .ZN(n673) );
  XOR2_X1 U748 ( .A(KEYINPUT20), .B(KEYINPUT90), .Z(n672) );
  XNOR2_X1 U749 ( .A(n673), .B(n672), .ZN(n674) );
  NAND2_X1 U750 ( .A1(G2090), .A2(n674), .ZN(n675) );
  XNOR2_X1 U751 ( .A(KEYINPUT21), .B(n675), .ZN(n676) );
  NAND2_X1 U752 ( .A1(n676), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U753 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U754 ( .A1(G120), .A2(G69), .ZN(n677) );
  NOR2_X1 U755 ( .A1(G237), .A2(n677), .ZN(n678) );
  NAND2_X1 U756 ( .A1(G108), .A2(n678), .ZN(n847) );
  NAND2_X1 U757 ( .A1(n847), .A2(G567), .ZN(n685) );
  XOR2_X1 U758 ( .A(KEYINPUT22), .B(KEYINPUT91), .Z(n680) );
  NAND2_X1 U759 ( .A1(G132), .A2(G82), .ZN(n679) );
  XNOR2_X1 U760 ( .A(n680), .B(n679), .ZN(n681) );
  NOR2_X1 U761 ( .A1(n681), .A2(G218), .ZN(n682) );
  NAND2_X1 U762 ( .A1(G96), .A2(n682), .ZN(n846) );
  NAND2_X1 U763 ( .A1(G2106), .A2(n846), .ZN(n683) );
  XNOR2_X1 U764 ( .A(KEYINPUT92), .B(n683), .ZN(n684) );
  NAND2_X1 U765 ( .A1(n685), .A2(n684), .ZN(n848) );
  NAND2_X1 U766 ( .A1(G483), .A2(G661), .ZN(n686) );
  NOR2_X1 U767 ( .A1(n848), .A2(n686), .ZN(n845) );
  NAND2_X1 U768 ( .A1(n845), .A2(G36), .ZN(G176) );
  NAND2_X1 U769 ( .A1(G101), .A2(n893), .ZN(n687) );
  XOR2_X1 U770 ( .A(KEYINPUT23), .B(n687), .Z(n691) );
  NAND2_X1 U771 ( .A1(n688), .A2(G125), .ZN(n689) );
  XOR2_X1 U772 ( .A(KEYINPUT67), .B(n689), .Z(n690) );
  NAND2_X1 U773 ( .A1(n691), .A2(n690), .ZN(n695) );
  NAND2_X1 U774 ( .A1(G113), .A2(n901), .ZN(n693) );
  NAND2_X1 U775 ( .A1(G137), .A2(n894), .ZN(n692) );
  NAND2_X1 U776 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U777 ( .A1(n695), .A2(n694), .ZN(G160) );
  NOR2_X1 U778 ( .A1(n696), .A2(G1384), .ZN(n697) );
  XOR2_X1 U779 ( .A(KEYINPUT65), .B(n697), .Z(n765) );
  INV_X1 U780 ( .A(n765), .ZN(n698) );
  NAND2_X1 U781 ( .A1(G160), .A2(G40), .ZN(n764) );
  NAND2_X1 U782 ( .A1(n722), .A2(G2072), .ZN(n699) );
  XNOR2_X1 U783 ( .A(n699), .B(KEYINPUT27), .ZN(n701) );
  INV_X1 U784 ( .A(G1956), .ZN(n1008) );
  NOR2_X1 U785 ( .A1(n1008), .A2(n722), .ZN(n700) );
  NOR2_X1 U786 ( .A1(n701), .A2(n700), .ZN(n717) );
  NAND2_X1 U787 ( .A1(n716), .A2(n717), .ZN(n715) );
  INV_X1 U788 ( .A(G1996), .ZN(n963) );
  NOR2_X1 U789 ( .A1(n738), .A2(n963), .ZN(n702) );
  XNOR2_X1 U790 ( .A(n702), .B(KEYINPUT26), .ZN(n706) );
  NAND2_X1 U791 ( .A1(n738), .A2(G1341), .ZN(n704) );
  INV_X1 U792 ( .A(n981), .ZN(n703) );
  NAND2_X1 U793 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U794 ( .A1(n706), .A2(n705), .ZN(n710) );
  NAND2_X1 U795 ( .A1(G1348), .A2(n738), .ZN(n708) );
  NAND2_X1 U796 ( .A1(G2067), .A2(n722), .ZN(n707) );
  NAND2_X1 U797 ( .A1(n708), .A2(n707), .ZN(n711) );
  NOR2_X1 U798 ( .A1(n988), .A2(n711), .ZN(n709) );
  OR2_X1 U799 ( .A1(n710), .A2(n709), .ZN(n713) );
  NAND2_X1 U800 ( .A1(n988), .A2(n711), .ZN(n712) );
  NAND2_X1 U801 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U802 ( .A1(n715), .A2(n714), .ZN(n719) );
  NOR2_X1 U803 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U804 ( .A1(n719), .A2(n523), .ZN(n721) );
  XOR2_X1 U805 ( .A(G1961), .B(KEYINPUT100), .Z(n1007) );
  NAND2_X1 U806 ( .A1(n1007), .A2(n738), .ZN(n724) );
  XNOR2_X1 U807 ( .A(KEYINPUT25), .B(G2078), .ZN(n961) );
  NAND2_X1 U808 ( .A1(n722), .A2(n961), .ZN(n723) );
  NAND2_X1 U809 ( .A1(n724), .A2(n723), .ZN(n730) );
  NAND2_X1 U810 ( .A1(n730), .A2(G171), .ZN(n725) );
  NAND2_X1 U811 ( .A1(n726), .A2(n725), .ZN(n736) );
  INV_X1 U812 ( .A(KEYINPUT31), .ZN(n734) );
  NOR2_X1 U813 ( .A1(G1966), .A2(n810), .ZN(n748) );
  NOR2_X1 U814 ( .A1(G2084), .A2(n738), .ZN(n747) );
  NOR2_X1 U815 ( .A1(n748), .A2(n747), .ZN(n727) );
  NAND2_X1 U816 ( .A1(G8), .A2(n727), .ZN(n728) );
  XNOR2_X1 U817 ( .A(KEYINPUT30), .B(n728), .ZN(n729) );
  NOR2_X1 U818 ( .A1(n729), .A2(G168), .ZN(n732) );
  NOR2_X1 U819 ( .A1(G171), .A2(n730), .ZN(n731) );
  XNOR2_X1 U820 ( .A(n734), .B(n733), .ZN(n735) );
  NAND2_X1 U821 ( .A1(n736), .A2(n735), .ZN(n751) );
  AND2_X1 U822 ( .A1(G286), .A2(G8), .ZN(n737) );
  NAND2_X1 U823 ( .A1(n751), .A2(n737), .ZN(n745) );
  INV_X1 U824 ( .A(G8), .ZN(n743) );
  NOR2_X1 U825 ( .A1(G1971), .A2(n810), .ZN(n740) );
  NOR2_X1 U826 ( .A1(G2090), .A2(n738), .ZN(n739) );
  NOR2_X1 U827 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U828 ( .A1(n741), .A2(G303), .ZN(n742) );
  OR2_X1 U829 ( .A1(n743), .A2(n742), .ZN(n744) );
  AND2_X1 U830 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U831 ( .A(n746), .B(KEYINPUT32), .ZN(n754) );
  AND2_X1 U832 ( .A1(G8), .A2(n747), .ZN(n749) );
  NOR2_X1 U833 ( .A1(n749), .A2(n748), .ZN(n750) );
  AND2_X1 U834 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U835 ( .A(KEYINPUT101), .B(n752), .ZN(n753) );
  NAND2_X1 U836 ( .A1(n754), .A2(n753), .ZN(n763) );
  NOR2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n984) );
  NOR2_X1 U838 ( .A1(G1971), .A2(G303), .ZN(n755) );
  NOR2_X1 U839 ( .A1(n984), .A2(n755), .ZN(n756) );
  NAND2_X1 U840 ( .A1(n763), .A2(n756), .ZN(n757) );
  XOR2_X1 U841 ( .A(n757), .B(KEYINPUT102), .Z(n758) );
  NOR2_X1 U842 ( .A1(n810), .A2(n758), .ZN(n759) );
  NAND2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n986) );
  NAND2_X1 U844 ( .A1(n759), .A2(n986), .ZN(n760) );
  INV_X1 U845 ( .A(KEYINPUT103), .ZN(n806) );
  NOR2_X1 U846 ( .A1(n810), .A2(n806), .ZN(n816) );
  NOR2_X1 U847 ( .A1(G2090), .A2(G303), .ZN(n761) );
  NAND2_X1 U848 ( .A1(G8), .A2(n761), .ZN(n762) );
  NAND2_X1 U849 ( .A1(n763), .A2(n762), .ZN(n798) );
  NOR2_X1 U850 ( .A1(n765), .A2(n764), .ZN(n836) );
  NAND2_X1 U851 ( .A1(G104), .A2(n893), .ZN(n767) );
  NAND2_X1 U852 ( .A1(G140), .A2(n894), .ZN(n766) );
  NAND2_X1 U853 ( .A1(n767), .A2(n766), .ZN(n769) );
  XOR2_X1 U854 ( .A(KEYINPUT34), .B(KEYINPUT95), .Z(n768) );
  XNOR2_X1 U855 ( .A(n769), .B(n768), .ZN(n774) );
  NAND2_X1 U856 ( .A1(n901), .A2(G116), .ZN(n771) );
  NAND2_X1 U857 ( .A1(G128), .A2(n898), .ZN(n770) );
  NAND2_X1 U858 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U859 ( .A(KEYINPUT35), .B(n772), .Z(n773) );
  NOR2_X1 U860 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U861 ( .A(KEYINPUT36), .B(n775), .ZN(n890) );
  XNOR2_X1 U862 ( .A(G2067), .B(KEYINPUT37), .ZN(n834) );
  NOR2_X1 U863 ( .A1(n890), .A2(n834), .ZN(n938) );
  NAND2_X1 U864 ( .A1(n836), .A2(n938), .ZN(n776) );
  XNOR2_X1 U865 ( .A(KEYINPUT96), .B(n776), .ZN(n832) );
  NAND2_X1 U866 ( .A1(G95), .A2(n893), .ZN(n778) );
  NAND2_X1 U867 ( .A1(G131), .A2(n894), .ZN(n777) );
  NAND2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n783) );
  NAND2_X1 U869 ( .A1(n901), .A2(G107), .ZN(n780) );
  NAND2_X1 U870 ( .A1(G119), .A2(n898), .ZN(n779) );
  NAND2_X1 U871 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U872 ( .A(KEYINPUT97), .B(n781), .Z(n782) );
  NOR2_X1 U873 ( .A1(n783), .A2(n782), .ZN(n885) );
  INV_X1 U874 ( .A(G1991), .ZN(n825) );
  NOR2_X1 U875 ( .A1(n885), .A2(n825), .ZN(n793) );
  XOR2_X1 U876 ( .A(KEYINPUT38), .B(KEYINPUT98), .Z(n785) );
  NAND2_X1 U877 ( .A1(G105), .A2(n893), .ZN(n784) );
  XNOR2_X1 U878 ( .A(n785), .B(n784), .ZN(n789) );
  NAND2_X1 U879 ( .A1(n901), .A2(G117), .ZN(n787) );
  NAND2_X1 U880 ( .A1(G129), .A2(n898), .ZN(n786) );
  NAND2_X1 U881 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U882 ( .A1(n789), .A2(n788), .ZN(n791) );
  NAND2_X1 U883 ( .A1(n894), .A2(G141), .ZN(n790) );
  NAND2_X1 U884 ( .A1(n791), .A2(n790), .ZN(n889) );
  AND2_X1 U885 ( .A1(G1996), .A2(n889), .ZN(n792) );
  NOR2_X1 U886 ( .A1(n793), .A2(n792), .ZN(n936) );
  INV_X1 U887 ( .A(n836), .ZN(n794) );
  NOR2_X1 U888 ( .A1(n936), .A2(n794), .ZN(n828) );
  INV_X1 U889 ( .A(n828), .ZN(n795) );
  NAND2_X1 U890 ( .A1(n832), .A2(n795), .ZN(n796) );
  XNOR2_X1 U891 ( .A(KEYINPUT99), .B(n796), .ZN(n811) );
  AND2_X1 U892 ( .A1(n810), .A2(n811), .ZN(n797) );
  NAND2_X1 U893 ( .A1(n798), .A2(n797), .ZN(n804) );
  INV_X1 U894 ( .A(n811), .ZN(n802) );
  NOR2_X1 U895 ( .A1(G1981), .A2(G305), .ZN(n799) );
  XOR2_X1 U896 ( .A(n799), .B(KEYINPUT24), .Z(n800) );
  OR2_X1 U897 ( .A1(n810), .A2(n800), .ZN(n801) );
  OR2_X1 U898 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U899 ( .A1(n804), .A2(n803), .ZN(n817) );
  NAND2_X1 U900 ( .A1(n984), .A2(KEYINPUT33), .ZN(n805) );
  NAND2_X1 U901 ( .A1(n806), .A2(n805), .ZN(n808) );
  NAND2_X1 U902 ( .A1(n984), .A2(KEYINPUT103), .ZN(n807) );
  NAND2_X1 U903 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n813) );
  XOR2_X1 U905 ( .A(G1981), .B(G305), .Z(n1000) );
  NAND2_X1 U906 ( .A1(n1000), .A2(n811), .ZN(n812) );
  NOR2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n814) );
  OR2_X1 U908 ( .A1(n817), .A2(n814), .ZN(n819) );
  INV_X1 U909 ( .A(n819), .ZN(n815) );
  NAND2_X1 U910 ( .A1(n526), .A2(n524), .ZN(n820) );
  OR2_X1 U911 ( .A1(KEYINPUT33), .A2(n817), .ZN(n818) );
  NAND2_X1 U912 ( .A1(n820), .A2(n525), .ZN(n821) );
  XNOR2_X1 U913 ( .A(n821), .B(KEYINPUT104), .ZN(n823) );
  XNOR2_X1 U914 ( .A(G1986), .B(G290), .ZN(n998) );
  NAND2_X1 U915 ( .A1(n998), .A2(n836), .ZN(n822) );
  NAND2_X1 U916 ( .A1(n823), .A2(n822), .ZN(n839) );
  NOR2_X1 U917 ( .A1(G1996), .A2(n889), .ZN(n824) );
  XOR2_X1 U918 ( .A(KEYINPUT105), .B(n824), .Z(n947) );
  NOR2_X1 U919 ( .A1(G1986), .A2(G290), .ZN(n826) );
  AND2_X1 U920 ( .A1(n825), .A2(n885), .ZN(n934) );
  NOR2_X1 U921 ( .A1(n826), .A2(n934), .ZN(n827) );
  NOR2_X1 U922 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U923 ( .A(n829), .B(KEYINPUT106), .ZN(n830) );
  NOR2_X1 U924 ( .A1(n947), .A2(n830), .ZN(n831) );
  XNOR2_X1 U925 ( .A(n831), .B(KEYINPUT39), .ZN(n833) );
  NAND2_X1 U926 ( .A1(n833), .A2(n832), .ZN(n835) );
  NAND2_X1 U927 ( .A1(n890), .A2(n834), .ZN(n931) );
  NAND2_X1 U928 ( .A1(n835), .A2(n931), .ZN(n837) );
  NAND2_X1 U929 ( .A1(n837), .A2(n836), .ZN(n838) );
  NAND2_X1 U930 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U931 ( .A(KEYINPUT40), .B(n840), .ZN(G329) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n841), .ZN(G217) );
  NAND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n842) );
  XOR2_X1 U934 ( .A(KEYINPUT108), .B(n842), .Z(n843) );
  NAND2_X1 U935 ( .A1(G661), .A2(n843), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U937 ( .A1(n845), .A2(n844), .ZN(G188) );
  XNOR2_X1 U938 ( .A(G69), .B(KEYINPUT109), .ZN(G235) );
  INV_X1 U940 ( .A(G132), .ZN(G219) );
  INV_X1 U941 ( .A(G120), .ZN(G236) );
  INV_X1 U942 ( .A(G96), .ZN(G221) );
  INV_X1 U943 ( .A(G82), .ZN(G220) );
  NOR2_X1 U944 ( .A1(n847), .A2(n846), .ZN(G325) );
  INV_X1 U945 ( .A(G325), .ZN(G261) );
  INV_X1 U946 ( .A(n848), .ZN(G319) );
  XOR2_X1 U947 ( .A(G2100), .B(G2096), .Z(n850) );
  XNOR2_X1 U948 ( .A(KEYINPUT42), .B(G2678), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U950 ( .A(KEYINPUT43), .B(G2090), .Z(n852) );
  XNOR2_X1 U951 ( .A(G2067), .B(G2072), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U953 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U954 ( .A(G2078), .B(G2084), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(G227) );
  XOR2_X1 U956 ( .A(KEYINPUT41), .B(G1981), .Z(n858) );
  XNOR2_X1 U957 ( .A(G1996), .B(G1991), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U959 ( .A(n859), .B(KEYINPUT111), .Z(n861) );
  XNOR2_X1 U960 ( .A(G1971), .B(G1976), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U962 ( .A(G1956), .B(G1961), .Z(n863) );
  XNOR2_X1 U963 ( .A(G1986), .B(G1966), .ZN(n862) );
  XNOR2_X1 U964 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U965 ( .A(n865), .B(n864), .Z(n867) );
  XNOR2_X1 U966 ( .A(KEYINPUT110), .B(G2474), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n867), .B(n866), .ZN(G229) );
  NAND2_X1 U968 ( .A1(n898), .A2(G124), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n868), .B(KEYINPUT44), .ZN(n875) );
  NAND2_X1 U970 ( .A1(G100), .A2(n893), .ZN(n870) );
  NAND2_X1 U971 ( .A1(G112), .A2(n901), .ZN(n869) );
  NAND2_X1 U972 ( .A1(n870), .A2(n869), .ZN(n873) );
  NAND2_X1 U973 ( .A1(n894), .A2(G136), .ZN(n871) );
  XOR2_X1 U974 ( .A(KEYINPUT112), .B(n871), .Z(n872) );
  NOR2_X1 U975 ( .A1(n873), .A2(n872), .ZN(n874) );
  NAND2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U977 ( .A(KEYINPUT113), .B(n876), .ZN(G162) );
  XOR2_X1 U978 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n887) );
  NAND2_X1 U979 ( .A1(G103), .A2(n893), .ZN(n878) );
  NAND2_X1 U980 ( .A1(G139), .A2(n894), .ZN(n877) );
  NAND2_X1 U981 ( .A1(n878), .A2(n877), .ZN(n883) );
  NAND2_X1 U982 ( .A1(n901), .A2(G115), .ZN(n880) );
  NAND2_X1 U983 ( .A1(G127), .A2(n898), .ZN(n879) );
  NAND2_X1 U984 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U985 ( .A(KEYINPUT47), .B(n881), .Z(n882) );
  NOR2_X1 U986 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U987 ( .A(KEYINPUT115), .B(n884), .Z(n941) );
  XNOR2_X1 U988 ( .A(n885), .B(n941), .ZN(n886) );
  XNOR2_X1 U989 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U990 ( .A(G162), .B(n888), .ZN(n892) );
  XOR2_X1 U991 ( .A(n890), .B(n889), .Z(n891) );
  XNOR2_X1 U992 ( .A(n892), .B(n891), .ZN(n906) );
  NAND2_X1 U993 ( .A1(G106), .A2(n893), .ZN(n896) );
  NAND2_X1 U994 ( .A1(G142), .A2(n894), .ZN(n895) );
  NAND2_X1 U995 ( .A1(n896), .A2(n895), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n897), .B(KEYINPUT45), .ZN(n900) );
  NAND2_X1 U997 ( .A1(G130), .A2(n898), .ZN(n899) );
  NAND2_X1 U998 ( .A1(n900), .A2(n899), .ZN(n904) );
  NAND2_X1 U999 ( .A1(n901), .A2(G118), .ZN(n902) );
  XOR2_X1 U1000 ( .A(KEYINPUT114), .B(n902), .Z(n903) );
  NOR2_X1 U1001 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U1002 ( .A(n906), .B(n905), .Z(n908) );
  XNOR2_X1 U1003 ( .A(G164), .B(G160), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1005 ( .A(n909), .B(n935), .Z(n910) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n910), .ZN(G395) );
  XNOR2_X1 U1007 ( .A(G286), .B(n988), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1009 ( .A(G171), .B(n913), .Z(n914) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n914), .ZN(G397) );
  XOR2_X1 U1011 ( .A(G2454), .B(G2430), .Z(n916) );
  XNOR2_X1 U1012 ( .A(G2451), .B(G2446), .ZN(n915) );
  XNOR2_X1 U1013 ( .A(n916), .B(n915), .ZN(n923) );
  XOR2_X1 U1014 ( .A(G2443), .B(G2427), .Z(n918) );
  XNOR2_X1 U1015 ( .A(G2438), .B(KEYINPUT107), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(n918), .B(n917), .ZN(n919) );
  XOR2_X1 U1017 ( .A(n919), .B(G2435), .Z(n921) );
  XNOR2_X1 U1018 ( .A(G1341), .B(G1348), .ZN(n920) );
  XNOR2_X1 U1019 ( .A(n921), .B(n920), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(n923), .B(n922), .ZN(n924) );
  NAND2_X1 U1021 ( .A1(n924), .A2(G14), .ZN(n930) );
  NAND2_X1 U1022 ( .A1(G319), .A2(n930), .ZN(n927) );
  NOR2_X1 U1023 ( .A1(G227), .A2(G229), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(KEYINPUT49), .B(n925), .ZN(n926) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n929) );
  NOR2_X1 U1026 ( .A1(G395), .A2(G397), .ZN(n928) );
  NAND2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(G225) );
  INV_X1 U1028 ( .A(G225), .ZN(G308) );
  INV_X1 U1029 ( .A(G108), .ZN(G238) );
  INV_X1 U1030 ( .A(n930), .ZN(G401) );
  XNOR2_X1 U1031 ( .A(G2084), .B(G160), .ZN(n932) );
  NAND2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(n940) );
  NAND2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n952) );
  XOR2_X1 U1037 ( .A(G2072), .B(n941), .Z(n943) );
  XOR2_X1 U1038 ( .A(G164), .B(G2078), .Z(n942) );
  NOR2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1040 ( .A(n944), .B(KEYINPUT116), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(n945), .B(KEYINPUT50), .ZN(n950) );
  XOR2_X1 U1042 ( .A(G2090), .B(G162), .Z(n946) );
  NOR2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1044 ( .A(KEYINPUT51), .B(n948), .Z(n949) );
  NAND2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(KEYINPUT52), .B(n953), .ZN(n955) );
  INV_X1 U1048 ( .A(KEYINPUT55), .ZN(n954) );
  NAND2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1050 ( .A1(n956), .A2(G29), .ZN(n1039) );
  XOR2_X1 U1051 ( .A(G2090), .B(G35), .Z(n960) );
  XOR2_X1 U1052 ( .A(G2084), .B(G34), .Z(n957) );
  XNOR2_X1 U1053 ( .A(KEYINPUT120), .B(n957), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(n958), .B(KEYINPUT54), .ZN(n959) );
  NAND2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n977) );
  XNOR2_X1 U1056 ( .A(n961), .B(G27), .ZN(n973) );
  XNOR2_X1 U1057 ( .A(KEYINPUT117), .B(G2067), .ZN(n962) );
  XNOR2_X1 U1058 ( .A(n962), .B(G26), .ZN(n968) );
  XNOR2_X1 U1059 ( .A(G32), .B(n963), .ZN(n964) );
  NAND2_X1 U1060 ( .A1(n964), .A2(G28), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(G25), .B(G1991), .ZN(n965) );
  NOR2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(KEYINPUT118), .B(G2072), .ZN(n969) );
  XNOR2_X1 U1065 ( .A(G33), .B(n969), .ZN(n970) );
  NOR2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(n974), .B(KEYINPUT119), .ZN(n975) );
  XNOR2_X1 U1069 ( .A(n975), .B(KEYINPUT53), .ZN(n976) );
  NOR2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1071 ( .A(KEYINPUT55), .B(n978), .Z(n979) );
  NOR2_X1 U1072 ( .A1(G29), .A2(n979), .ZN(n1035) );
  INV_X1 U1073 ( .A(G16), .ZN(n1031) );
  XNOR2_X1 U1074 ( .A(KEYINPUT56), .B(KEYINPUT121), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(n1031), .B(n980), .ZN(n1006) );
  XOR2_X1 U1076 ( .A(G171), .B(G1961), .Z(n983) );
  XNOR2_X1 U1077 ( .A(n981), .B(G1341), .ZN(n982) );
  NOR2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n996) );
  XOR2_X1 U1079 ( .A(n984), .B(KEYINPUT122), .Z(n985) );
  NAND2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1081 ( .A(n987), .B(KEYINPUT123), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(n988), .B(G1348), .ZN(n990) );
  XNOR2_X1 U1083 ( .A(G299), .B(G1956), .ZN(n989) );
  NOR2_X1 U1084 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n994) );
  XNOR2_X1 U1086 ( .A(G1971), .B(G303), .ZN(n993) );
  NOR2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1090 ( .A(KEYINPUT124), .B(n999), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(G1966), .B(G168), .ZN(n1001) );
  NAND2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(KEYINPUT57), .B(n1002), .ZN(n1003) );
  NAND2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1033) );
  XNOR2_X1 U1096 ( .A(n1007), .B(G5), .ZN(n1020) );
  XNOR2_X1 U1097 ( .A(G20), .B(n1008), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(G1341), .B(G19), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(G1981), .B(G6), .ZN(n1009) );
  NOR2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1015) );
  XOR2_X1 U1102 ( .A(KEYINPUT59), .B(G1348), .Z(n1013) );
  XNOR2_X1 U1103 ( .A(G4), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1105 ( .A(KEYINPUT60), .B(n1016), .Z(n1018) );
  XNOR2_X1 U1106 ( .A(G1966), .B(G21), .ZN(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1028) );
  XNOR2_X1 U1109 ( .A(G1986), .B(G24), .ZN(n1022) );
  XNOR2_X1 U1110 ( .A(G23), .B(G1976), .ZN(n1021) );
  NOR2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1025) );
  XNOR2_X1 U1112 ( .A(G1971), .B(KEYINPUT125), .ZN(n1023) );
  XNOR2_X1 U1113 ( .A(n1023), .B(G22), .ZN(n1024) );
  NAND2_X1 U1114 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1115 ( .A(KEYINPUT58), .B(n1026), .ZN(n1027) );
  NOR2_X1 U1116 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1117 ( .A(KEYINPUT61), .B(n1029), .ZN(n1030) );
  NAND2_X1 U1118 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1119 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NOR2_X1 U1120 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1121 ( .A1(G11), .A2(n1036), .ZN(n1037) );
  XOR2_X1 U1122 ( .A(KEYINPUT126), .B(n1037), .Z(n1038) );
  NAND2_X1 U1123 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  XNOR2_X1 U1124 ( .A(n1040), .B(KEYINPUT127), .ZN(n1041) );
  XNOR2_X1 U1125 ( .A(KEYINPUT62), .B(n1041), .ZN(G311) );
  INV_X1 U1126 ( .A(G311), .ZN(G150) );
endmodule

