//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 1 0 0 1 0 0 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1221, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1280, new_n1281;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  NAND2_X1  g0011(.A1(G116), .A2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G77), .ZN(new_n213));
  INV_X1    g0013(.A(G244), .ZN(new_n214));
  INV_X1    g0014(.A(G87), .ZN(new_n215));
  INV_X1    g0015(.A(G250), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  INV_X1    g0018(.A(G226), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n202), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI211_X1 g0022(.A(new_n217), .B(new_n222), .C1(G97), .C2(G257), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(G1), .B2(G20), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT1), .Z(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(new_n201), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n211), .B(new_n225), .C1(new_n228), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT64), .B(G264), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT65), .ZN(new_n243));
  INV_X1    g0043(.A(G107), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  NAND2_X1  g0051(.A1(new_n220), .A2(G20), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n227), .A2(G33), .A3(G77), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  AND3_X1   g0054(.A1(new_n227), .A2(new_n254), .A3(KEYINPUT69), .ZN(new_n255));
  AOI21_X1  g0055(.A(KEYINPUT69), .B1(new_n227), .B2(new_n254), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n252), .B(new_n253), .C1(new_n257), .C2(new_n202), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n226), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT68), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n259), .A2(KEYINPUT68), .A3(new_n226), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n258), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT11), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G13), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(G1), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G20), .A3(new_n220), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n270), .B(KEYINPUT12), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(G20), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT70), .ZN(new_n274));
  INV_X1    g0074(.A(G1), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n274), .B1(new_n275), .B2(G20), .ZN(new_n276));
  NOR3_X1   g0076(.A1(new_n227), .A2(KEYINPUT70), .A3(G1), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NOR3_X1   g0078(.A1(new_n264), .A2(new_n273), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G68), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n258), .A2(KEYINPUT11), .A3(new_n264), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n267), .A2(new_n271), .A3(new_n280), .A4(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(new_n282), .B(KEYINPUT74), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT13), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n275), .B1(G41), .B2(G45), .ZN(new_n285));
  INV_X1    g0085(.A(G274), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n219), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G232), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G1698), .ZN(new_n291));
  AND2_X1   g0091(.A1(KEYINPUT3), .A2(G33), .ZN(new_n292));
  NOR2_X1   g0092(.A1(KEYINPUT3), .A2(G33), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n289), .B(new_n291), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G97), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G33), .A2(G41), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n297), .A2(G1), .A3(G13), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n287), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  AND3_X1   g0100(.A1(new_n298), .A2(G238), .A3(new_n285), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n284), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n298), .B1(new_n294), .B2(new_n295), .ZN(new_n304));
  NOR4_X1   g0104(.A1(new_n304), .A2(KEYINPUT13), .A3(new_n301), .A4(new_n287), .ZN(new_n305));
  OAI21_X1  g0105(.A(G169), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT14), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n307), .A2(KEYINPUT75), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  OAI221_X1 g0109(.A(G169), .B1(KEYINPUT75), .B2(new_n307), .C1(new_n303), .C2(new_n305), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n303), .A2(new_n305), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G179), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n309), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT76), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT76), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n309), .A2(new_n310), .A3(new_n312), .A4(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n283), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n311), .A2(G190), .ZN(new_n318));
  INV_X1    g0118(.A(G200), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT73), .B1(new_n311), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT73), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n321), .B(G200), .C1(new_n303), .C2(new_n305), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  AND3_X1   g0123(.A1(new_n283), .A2(new_n318), .A3(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n317), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT3), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n254), .ZN(new_n327));
  NAND2_X1  g0127(.A1(KEYINPUT3), .A2(G33), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(G222), .A2(G1698), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n288), .A2(G223), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(G77), .B2(new_n329), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n333), .B(KEYINPUT67), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n287), .B1(new_n334), .B2(new_n299), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n298), .A2(new_n285), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  OR2_X1    g0137(.A1(KEYINPUT66), .A2(G226), .ZN(new_n338));
  NAND2_X1  g0138(.A1(KEYINPUT66), .A2(G226), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n335), .A2(G190), .A3(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(G50), .B1(new_n276), .B2(new_n277), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n342), .B(KEYINPUT71), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n264), .A2(new_n273), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n273), .A2(new_n202), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n203), .A2(G20), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT8), .B(G58), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n227), .A2(G33), .ZN(new_n349));
  INV_X1    g0149(.A(G150), .ZN(new_n350));
  OAI221_X1 g0150(.A(new_n347), .B1(new_n348), .B2(new_n349), .C1(new_n257), .C2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n264), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n345), .A2(new_n346), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT9), .ZN(new_n354));
  OR2_X1    g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n341), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT10), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n319), .B1(new_n335), .B2(new_n340), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n353), .A2(new_n354), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n356), .A2(new_n357), .A3(new_n359), .A4(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n341), .A2(new_n355), .A3(new_n360), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT10), .B1(new_n362), .B2(new_n358), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n325), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n335), .A2(new_n340), .ZN(new_n366));
  INV_X1    g0166(.A(G169), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G179), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n335), .A2(new_n369), .A3(new_n340), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n370), .A3(new_n353), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT72), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n368), .A2(KEYINPUT72), .A3(new_n370), .A4(new_n353), .ZN(new_n374));
  INV_X1    g0174(.A(new_n257), .ZN(new_n375));
  XOR2_X1   g0175(.A(KEYINPUT8), .B(G58), .Z(new_n376));
  AOI22_X1  g0176(.A1(new_n375), .A2(new_n376), .B1(G20), .B2(G77), .ZN(new_n377));
  XOR2_X1   g0177(.A(KEYINPUT15), .B(G87), .Z(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n377), .B1(new_n349), .B2(new_n379), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n380), .A2(new_n264), .B1(G77), .B2(new_n279), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(G77), .B2(new_n272), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G238), .A2(G1698), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n329), .B(new_n383), .C1(new_n290), .C2(G1698), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n384), .B(new_n299), .C1(G107), .C2(new_n329), .ZN(new_n385));
  INV_X1    g0185(.A(new_n287), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n385), .B(new_n386), .C1(new_n214), .C2(new_n336), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G169), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n369), .B2(new_n387), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n382), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n387), .A2(G200), .ZN(new_n391));
  INV_X1    g0191(.A(G190), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n391), .B1(new_n392), .B2(new_n387), .ZN(new_n393));
  OR2_X1    g0193(.A1(new_n382), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n373), .A2(new_n374), .A3(new_n390), .A4(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n327), .A2(new_n227), .A3(new_n328), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n327), .A2(KEYINPUT7), .A3(new_n227), .A4(new_n328), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n220), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(G159), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n257), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G58), .A2(G68), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n227), .B1(new_n229), .B2(new_n403), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n400), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(KEYINPUT16), .B1(new_n405), .B2(KEYINPUT77), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT77), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT16), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n292), .A2(new_n293), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT7), .B1(new_n409), .B2(new_n227), .ZN(new_n410));
  INV_X1    g0210(.A(new_n399), .ZN(new_n411));
  OAI21_X1  g0211(.A(G68), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n404), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n407), .B(new_n408), .C1(new_n414), .C2(new_n402), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n406), .A2(new_n415), .A3(new_n264), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT78), .B1(new_n278), .B2(new_n348), .ZN(new_n417));
  AND3_X1   g0217(.A1(new_n259), .A2(KEYINPUT68), .A3(new_n226), .ZN(new_n418));
  AOI21_X1  g0218(.A(KEYINPUT68), .B1(new_n259), .B2(new_n226), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT78), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n376), .B(new_n421), .C1(new_n277), .C2(new_n276), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n417), .A2(new_n272), .A3(new_n420), .A4(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n273), .A2(new_n348), .ZN(new_n424));
  AND3_X1   g0224(.A1(new_n423), .A2(KEYINPUT79), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(KEYINPUT79), .B1(new_n423), .B2(new_n424), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n219), .A2(G1698), .ZN(new_n428));
  OAI221_X1 g0228(.A(new_n428), .B1(G223), .B2(G1698), .C1(new_n292), .C2(new_n293), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G33), .A2(G87), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n298), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n336), .A2(new_n290), .ZN(new_n432));
  NOR3_X1   g0232(.A1(new_n431), .A2(new_n287), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n392), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n433), .B2(G200), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n416), .A2(new_n427), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT17), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n416), .A2(new_n427), .A3(KEYINPUT17), .A4(new_n435), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n416), .A2(new_n427), .ZN(new_n440));
  NOR4_X1   g0240(.A1(new_n431), .A2(new_n369), .A3(new_n432), .A4(new_n287), .ZN(new_n441));
  INV_X1    g0241(.A(new_n433), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n441), .B1(new_n442), .B2(G169), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT18), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT18), .ZN(new_n446));
  AOI211_X1 g0246(.A(new_n446), .B(new_n443), .C1(new_n416), .C2(new_n427), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n438), .B(new_n439), .C1(new_n445), .C2(new_n447), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n365), .A2(new_n395), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT21), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n269), .A2(G20), .A3(new_n246), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n275), .A2(G33), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n262), .A2(new_n272), .A3(new_n263), .A4(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n451), .B1(new_n453), .B2(new_n246), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n259), .A2(new_n226), .B1(G20), .B2(new_n246), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G283), .ZN(new_n456));
  INV_X1    g0256(.A(G97), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n456), .B(new_n227), .C1(G33), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(KEYINPUT83), .A2(KEYINPUT20), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT83), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT20), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n459), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n455), .A2(new_n461), .A3(new_n458), .A4(new_n462), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n454), .A2(new_n466), .ZN(new_n467));
  AND2_X1   g0267(.A1(KEYINPUT82), .A2(G303), .ZN(new_n468));
  NOR2_X1   g0268(.A1(KEYINPUT82), .A2(G303), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n327), .B(new_n328), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n288), .A2(G257), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G264), .A2(G1698), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n471), .B(new_n472), .C1(new_n292), .C2(new_n293), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n470), .A2(new_n473), .A3(new_n299), .ZN(new_n474));
  INV_X1    g0274(.A(G45), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(G1), .ZN(new_n476));
  AND2_X1   g0276(.A1(KEYINPUT5), .A2(G41), .ZN(new_n477));
  NOR2_X1   g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n479), .A2(G270), .A3(new_n298), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n476), .B(G274), .C1(new_n478), .C2(new_n477), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n474), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G169), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n450), .B1(new_n467), .B2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n420), .A2(G116), .A3(new_n272), .A4(new_n452), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n485), .A2(new_n451), .A3(new_n465), .A4(new_n464), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n486), .A2(KEYINPUT21), .A3(G169), .A4(new_n482), .ZN(new_n487));
  AND4_X1   g0287(.A1(G179), .A2(new_n474), .A3(new_n480), .A4(new_n481), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n484), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT84), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n482), .A2(G200), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n491), .B1(new_n492), .B2(new_n486), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n482), .A2(G200), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n467), .A2(KEYINPUT84), .A3(new_n494), .ZN(new_n495));
  OR2_X1    g0295(.A1(new_n482), .A2(new_n392), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n493), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT85), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT85), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n493), .A2(new_n495), .A3(new_n499), .A4(new_n496), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n490), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n215), .A2(new_n457), .A3(new_n244), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n295), .A2(new_n227), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT19), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n227), .B(G68), .C1(new_n292), .C2(new_n293), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT19), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n506), .B1(new_n349), .B2(new_n457), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n504), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n508), .A2(new_n264), .B1(new_n273), .B2(new_n379), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n420), .A2(new_n272), .A3(new_n378), .A4(new_n452), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n221), .A2(new_n288), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n214), .A2(G1698), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n512), .B(new_n513), .C1(new_n292), .C2(new_n293), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G116), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n298), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n275), .A2(G45), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n298), .A2(G250), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n476), .A2(G274), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n369), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n367), .B1(new_n516), .B2(new_n520), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n511), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n520), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n514), .A2(new_n515), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n525), .B(G190), .C1(new_n526), .C2(new_n298), .ZN(new_n527));
  OAI21_X1  g0327(.A(G200), .B1(new_n516), .B2(new_n520), .ZN(new_n528));
  INV_X1    g0328(.A(new_n453), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G87), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n527), .A2(new_n528), .A3(new_n530), .A4(new_n509), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n524), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT4), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n534), .A2(G1698), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n535), .B(G244), .C1(new_n293), .C2(new_n292), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n214), .B1(new_n327), .B2(new_n328), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n536), .B(new_n456), .C1(new_n537), .C2(KEYINPUT4), .ZN(new_n538));
  OAI21_X1  g0338(.A(G250), .B1(new_n292), .B2(new_n293), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n288), .B1(new_n539), .B2(KEYINPUT4), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n299), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n479), .A2(G257), .A3(new_n298), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n481), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT81), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n542), .A2(KEYINPUT81), .A3(new_n481), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n541), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(G200), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n257), .A2(new_n213), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(G107), .B1(new_n410), .B2(new_n411), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT6), .ZN(new_n552));
  AND2_X1   g0352(.A1(G97), .A2(G107), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n552), .B1(new_n553), .B2(new_n205), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n244), .A2(KEYINPUT6), .A3(G97), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n227), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n550), .A2(new_n551), .A3(new_n557), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n558), .A2(new_n264), .B1(G97), .B2(new_n529), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n273), .A2(new_n457), .ZN(new_n560));
  XNOR2_X1  g0360(.A(new_n560), .B(KEYINPUT80), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n541), .A2(new_n545), .A3(G190), .A4(new_n546), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n548), .A2(new_n559), .A3(new_n561), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n547), .A2(new_n367), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n529), .A2(G97), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n244), .B1(new_n398), .B2(new_n399), .ZN(new_n566));
  NOR3_X1   g0366(.A1(new_n566), .A2(new_n549), .A3(new_n556), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n561), .B(new_n565), .C1(new_n567), .C2(new_n420), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n541), .A2(new_n545), .A3(new_n369), .A4(new_n546), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n564), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n227), .A2(G33), .A3(G116), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n227), .A2(G107), .ZN(new_n572));
  XNOR2_X1  g0372(.A(new_n572), .B(KEYINPUT23), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT22), .ZN(new_n574));
  AOI21_X1  g0374(.A(G20), .B1(new_n327), .B2(new_n328), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n574), .B1(new_n575), .B2(G87), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n227), .B(G87), .C1(new_n292), .C2(new_n293), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n577), .A2(KEYINPUT22), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n571), .B(new_n573), .C1(new_n576), .C2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT24), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g0381(.A(new_n577), .B(KEYINPUT22), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n582), .A2(KEYINPUT24), .A3(new_n571), .A4(new_n573), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n581), .A2(new_n583), .A3(new_n264), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n529), .A2(G107), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n216), .A2(new_n288), .ZN(new_n586));
  INV_X1    g0386(.A(G257), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(G1698), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n586), .B(new_n588), .C1(new_n292), .C2(new_n293), .ZN(new_n589));
  NAND2_X1  g0389(.A1(G33), .A2(G294), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n298), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n479), .A2(G264), .A3(new_n298), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n592), .A2(new_n392), .A3(new_n481), .A4(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n593), .ZN(new_n595));
  INV_X1    g0395(.A(new_n481), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n595), .A2(new_n591), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n594), .B1(new_n597), .B2(G200), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT86), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n273), .B(new_n244), .C1(new_n599), .C2(KEYINPUT25), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(KEYINPUT25), .ZN(new_n601));
  XNOR2_X1  g0401(.A(new_n600), .B(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n584), .A2(new_n585), .A3(new_n598), .A4(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n563), .A2(new_n570), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n584), .A2(new_n585), .A3(new_n602), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n597), .A2(G169), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(new_n369), .B2(new_n597), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  AND4_X1   g0409(.A1(new_n449), .A2(new_n501), .A3(new_n533), .A4(new_n609), .ZN(G372));
  AND3_X1   g0410(.A1(new_n524), .A2(new_n531), .A3(KEYINPUT87), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT87), .B1(new_n524), .B2(new_n531), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n604), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n490), .A2(KEYINPUT88), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT88), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n484), .A2(new_n616), .A3(new_n487), .A4(new_n489), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n614), .B1(new_n618), .B2(new_n608), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n564), .A2(new_n568), .A3(new_n569), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT26), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n620), .B(new_n621), .C1(new_n612), .C2(new_n611), .ZN(new_n622));
  OAI21_X1  g0422(.A(KEYINPUT26), .B1(new_n570), .B2(new_n532), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n622), .A2(new_n524), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n449), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g0426(.A(new_n626), .B(KEYINPUT89), .Z(new_n627));
  NAND2_X1  g0427(.A1(new_n373), .A2(new_n374), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n440), .A2(new_n444), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n446), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n440), .A2(KEYINPUT18), .A3(new_n444), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n324), .ZN(new_n633));
  INV_X1    g0433(.A(new_n390), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n633), .B1(new_n317), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n438), .A2(new_n439), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n628), .B1(new_n637), .B2(new_n364), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n627), .A2(new_n638), .ZN(G369));
  NOR2_X1   g0439(.A1(new_n268), .A2(G20), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n269), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n642), .A2(KEYINPUT90), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(KEYINPUT90), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n643), .A2(G213), .A3(new_n644), .A4(new_n645), .ZN(new_n646));
  XNOR2_X1  g0446(.A(KEYINPUT91), .B(G343), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n486), .ZN(new_n650));
  MUX2_X1   g0450(.A(new_n618), .B(new_n501), .S(new_n650), .Z(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(G330), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n605), .A2(new_n607), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n605), .A2(new_n649), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(new_n654), .A3(new_n603), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(KEYINPUT92), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT92), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n653), .A2(new_n654), .A3(new_n657), .A4(new_n603), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n649), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n653), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n652), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n653), .A2(new_n649), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n490), .A2(new_n660), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n665), .B1(new_n656), .B2(new_n658), .ZN(new_n666));
  OR3_X1    g0466(.A1(new_n663), .A2(new_n664), .A3(new_n666), .ZN(G399));
  INV_X1    g0467(.A(new_n209), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(G41), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n502), .A2(G116), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G1), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n230), .B2(new_n670), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT28), .ZN(new_n674));
  INV_X1    g0474(.A(new_n524), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n620), .B1(new_n611), .B2(new_n612), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n675), .B1(new_n676), .B2(KEYINPUT26), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n563), .A2(new_n570), .A3(new_n603), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n484), .A2(new_n487), .A3(new_n489), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n653), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n612), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n524), .A2(new_n531), .A3(KEYINPUT87), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n678), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n620), .A2(new_n621), .A3(new_n533), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n677), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n660), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT29), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n609), .A2(new_n501), .A3(new_n533), .A4(new_n660), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT93), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n482), .A2(new_n369), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n690), .B1(new_n691), .B2(new_n521), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n525), .B1(new_n526), .B2(new_n298), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n693), .A2(KEYINPUT93), .A3(new_n369), .A4(new_n482), .ZN(new_n694));
  INV_X1    g0494(.A(new_n597), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n692), .A2(new_n547), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n541), .A2(new_n545), .A3(new_n546), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n595), .A2(new_n591), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n698), .A2(new_n521), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n697), .A2(KEYINPUT30), .A3(new_n488), .A4(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT30), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n488), .A2(new_n541), .A3(new_n545), .A4(new_n546), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n698), .A2(new_n521), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n696), .A2(new_n700), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n649), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT31), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n705), .A2(KEYINPUT31), .A3(new_n649), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n689), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G330), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT29), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n625), .A2(new_n712), .A3(new_n660), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n688), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  OR2_X1    g0514(.A1(new_n714), .A2(KEYINPUT94), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(KEYINPUT94), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n674), .B1(new_n717), .B2(G1), .ZN(G364));
  NAND2_X1  g0518(.A1(new_n640), .A2(G45), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n670), .A2(G1), .A3(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n721), .B1(new_n651), .B2(G330), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(G330), .B2(new_n651), .ZN(new_n723));
  NOR2_X1   g0523(.A1(G13), .A2(G33), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G20), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n226), .B1(G20), .B2(new_n367), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n250), .A2(G45), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n729), .A2(KEYINPUT95), .B1(new_n475), .B2(new_n231), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n668), .A2(new_n329), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n730), .B(new_n731), .C1(KEYINPUT95), .C2(new_n729), .ZN(new_n732));
  INV_X1    g0532(.A(G355), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n329), .A2(new_n209), .ZN(new_n734));
  OAI221_X1 g0534(.A(new_n732), .B1(G116), .B2(new_n209), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n369), .A2(G200), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n227), .A2(G190), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G311), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n319), .A2(G179), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(G283), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G179), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n737), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G329), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n742), .A2(new_n743), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n369), .A2(new_n319), .ZN(new_n748));
  NAND2_X1  g0548(.A1(G20), .A2(G190), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  XOR2_X1   g0552(.A(KEYINPUT98), .B(G326), .Z(new_n753));
  AOI211_X1 g0553(.A(new_n740), .B(new_n747), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n749), .A2(new_n369), .A3(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G322), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n227), .B1(new_n744), .B2(G190), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G294), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n741), .A2(new_n750), .ZN(new_n760));
  INV_X1    g0560(.A(G303), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n409), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n748), .A2(new_n737), .ZN(new_n763));
  XNOR2_X1  g0563(.A(KEYINPUT33), .B(G317), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n754), .A2(new_n756), .A3(new_n759), .A4(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n745), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G159), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT96), .ZN(new_n769));
  XOR2_X1   g0569(.A(new_n769), .B(KEYINPUT32), .Z(new_n770));
  AND2_X1   g0570(.A1(new_n757), .A2(KEYINPUT97), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n757), .A2(KEYINPUT97), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G97), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n763), .A2(G68), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n751), .A2(new_n202), .B1(new_n742), .B2(new_n244), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n760), .A2(new_n215), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n755), .ZN(new_n780));
  INV_X1    g0580(.A(G58), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n329), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n738), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n782), .B1(G77), .B2(new_n783), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n775), .A2(new_n776), .A3(new_n779), .A4(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n766), .B1(new_n770), .B2(new_n785), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n728), .A2(new_n735), .B1(new_n786), .B2(new_n727), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n726), .B(KEYINPUT99), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n721), .B(new_n787), .C1(new_n651), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n723), .A2(new_n789), .ZN(G396));
  NOR2_X1   g0590(.A1(new_n742), .A2(new_n220), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n760), .A2(new_n202), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n757), .A2(new_n781), .ZN(new_n793));
  OR4_X1    g0593(.A1(new_n409), .A2(new_n791), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n763), .A2(G150), .B1(G143), .B2(new_n755), .ZN(new_n795));
  INV_X1    g0595(.A(G137), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n795), .B1(new_n796), .B2(new_n751), .C1(new_n401), .C2(new_n738), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT34), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n794), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G132), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n799), .B1(new_n798), .B2(new_n797), .C1(new_n800), .C2(new_n745), .ZN(new_n801));
  INV_X1    g0601(.A(G294), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n780), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n742), .A2(new_n215), .ZN(new_n804));
  INV_X1    g0604(.A(new_n760), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n804), .B1(G107), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(new_n739), .B2(new_n745), .ZN(new_n807));
  XOR2_X1   g0607(.A(KEYINPUT100), .B(G283), .Z(new_n808));
  AOI21_X1  g0608(.A(new_n807), .B1(new_n763), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n409), .B1(new_n751), .B2(new_n761), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(G116), .B2(new_n783), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n809), .A2(new_n775), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n801), .B1(new_n803), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT101), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n720), .B1(new_n814), .B2(new_n727), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n727), .A2(new_n724), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n634), .A2(KEYINPUT102), .A3(new_n649), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n382), .A2(new_n649), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n394), .A2(new_n390), .A3(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT102), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n390), .B2(new_n660), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n818), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n815), .B1(G77), .B2(new_n817), .C1(new_n725), .C2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n649), .B1(new_n619), .B2(new_n624), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(new_n823), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(new_n711), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n824), .B1(new_n827), .B2(new_n721), .ZN(G384));
  OR2_X1    g0628(.A1(new_n282), .A2(KEYINPUT74), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n282), .A2(KEYINPUT74), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n829), .A2(new_n830), .A3(new_n649), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NOR3_X1   g0632(.A1(new_n317), .A2(new_n324), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n831), .B1(new_n314), .B2(new_n316), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n823), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT104), .ZN(new_n836));
  AND3_X1   g0636(.A1(new_n705), .A2(new_n836), .A3(new_n649), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n836), .B1(new_n705), .B2(new_n649), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n839), .A2(KEYINPUT105), .A3(new_n707), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n706), .A2(KEYINPUT104), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n705), .A2(new_n836), .A3(new_n649), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n841), .A2(new_n707), .A3(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT105), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n709), .A2(KEYINPUT106), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT106), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n705), .A2(new_n848), .A3(KEYINPUT31), .A4(new_n649), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n850), .A2(new_n689), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n835), .B1(new_n846), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT38), .ZN(new_n853));
  INV_X1    g0653(.A(new_n646), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n440), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT37), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n629), .A2(new_n855), .A3(new_n856), .A4(new_n436), .ZN(new_n857));
  INV_X1    g0657(.A(new_n436), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n423), .A2(new_n424), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n416), .A2(new_n859), .B1(new_n443), .B2(new_n646), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT37), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n646), .B1(new_n416), .B2(new_n859), .ZN(new_n862));
  AOI221_X4 g0662(.A(new_n853), .B1(new_n857), .B2(new_n861), .C1(new_n448), .C2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n855), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n445), .A2(new_n447), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n864), .B1(new_n865), .B2(new_n636), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n416), .A2(new_n427), .B1(new_n443), .B2(new_n646), .ZN(new_n867));
  OAI21_X1  g0667(.A(KEYINPUT37), .B1(new_n858), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n857), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT38), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT107), .B1(new_n863), .B2(new_n870), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n438), .A2(new_n439), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n855), .B1(new_n632), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n857), .A2(new_n868), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n853), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT107), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n448), .A2(new_n862), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n857), .A2(new_n861), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n877), .A2(KEYINPUT38), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n875), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n852), .A2(new_n871), .A3(KEYINPUT40), .A4(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT40), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT105), .B1(new_n839), .B2(new_n707), .ZN(new_n883));
  NOR4_X1   g0683(.A1(new_n837), .A2(new_n838), .A3(new_n844), .A4(KEYINPUT31), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n851), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n823), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n325), .A2(new_n831), .ZN(new_n887));
  INV_X1    g0687(.A(new_n834), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT38), .B1(new_n877), .B2(new_n878), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n863), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n882), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n881), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n449), .A2(new_n885), .ZN(new_n895));
  XOR2_X1   g0695(.A(new_n894), .B(new_n895), .Z(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(G330), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT39), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n863), .B2(new_n870), .ZN(new_n899));
  INV_X1    g0699(.A(new_n862), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n632), .B2(new_n872), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n857), .A2(new_n861), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n853), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(KEYINPUT39), .A3(new_n879), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n899), .A2(new_n317), .A3(new_n660), .A4(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n390), .A2(new_n649), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n825), .B2(new_n823), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n834), .B1(new_n325), .B2(new_n831), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n908), .B(new_n910), .C1(new_n891), .C2(new_n863), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n865), .A2(new_n646), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n905), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n688), .A2(new_n713), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n449), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n638), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n913), .B(new_n916), .Z(new_n917));
  XNOR2_X1  g0717(.A(new_n897), .B(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n275), .B2(new_n640), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n554), .A2(new_n555), .ZN(new_n920));
  OAI211_X1 g0720(.A(G116), .B(new_n228), .C1(new_n920), .C2(KEYINPUT35), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT103), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n920), .A2(KEYINPUT35), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT36), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n403), .A2(G77), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n230), .A2(new_n926), .B1(G50), .B2(new_n220), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n927), .A2(G1), .A3(new_n268), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n919), .A2(new_n925), .A3(new_n928), .ZN(G367));
  INV_X1    g0729(.A(new_n666), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n568), .A2(new_n649), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n563), .A2(new_n570), .A3(new_n931), .ZN(new_n932));
  OR3_X1    g0732(.A1(new_n930), .A2(KEYINPUT42), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n570), .B1(new_n932), .B2(new_n653), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n660), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT42), .B1(new_n930), .B2(new_n932), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n933), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n530), .A2(new_n509), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n649), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n683), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n524), .B2(new_n939), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n937), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n620), .A2(new_n649), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n932), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n663), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n943), .B(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n947), .A2(new_n948), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n669), .B(KEYINPUT41), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n945), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n666), .B2(new_n664), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(KEYINPUT108), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT108), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n956), .B(new_n953), .C1(new_n666), .C2(new_n664), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT44), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n955), .A2(KEYINPUT44), .A3(new_n957), .ZN(new_n961));
  NOR3_X1   g0761(.A1(new_n666), .A2(new_n664), .A3(new_n953), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT45), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n960), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n663), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n662), .A2(new_n665), .ZN(new_n966));
  AND3_X1   g0766(.A1(new_n966), .A2(new_n652), .A3(new_n930), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n652), .B1(new_n966), .B2(new_n930), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n715), .B2(new_n716), .ZN(new_n970));
  INV_X1    g0770(.A(new_n663), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n960), .A2(new_n963), .A3(new_n971), .A4(new_n961), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n965), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n952), .B1(new_n973), .B2(new_n717), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n719), .A2(G1), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n949), .B(new_n950), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n329), .B1(new_n742), .B2(new_n213), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n760), .A2(new_n781), .B1(new_n745), .B2(new_n796), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(G159), .B2(new_n763), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n202), .B2(new_n738), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n977), .B(new_n980), .C1(G143), .C2(new_n752), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(new_n220), .B2(new_n773), .C1(new_n350), .C2(new_n780), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n805), .A2(KEYINPUT46), .A3(G116), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT46), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n760), .B2(new_n246), .ZN(new_n985));
  INV_X1    g0785(.A(new_n763), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n983), .B(new_n985), .C1(new_n802), .C2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT110), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n468), .A2(new_n469), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n752), .A2(G311), .B1(new_n990), .B2(new_n755), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT109), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n987), .A2(new_n988), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n742), .A2(new_n457), .ZN(new_n994));
  INV_X1    g0794(.A(G317), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n409), .B1(new_n745), .B2(new_n995), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n994), .B(new_n996), .C1(G107), .C2(new_n758), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n989), .A2(new_n992), .A3(new_n993), .A4(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n808), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n999), .A2(new_n738), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n982), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT47), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n720), .B1(new_n1002), .B2(new_n727), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n731), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n728), .B1(new_n209), .B2(new_n379), .C1(new_n240), .C2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1003), .B(new_n1005), .C1(new_n788), .C2(new_n941), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n976), .A2(new_n1006), .ZN(G387));
  INV_X1    g0807(.A(new_n969), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n717), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n715), .A2(new_n716), .A3(new_n969), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n669), .B(KEYINPUT113), .Z(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1009), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n763), .A2(G311), .B1(G317), .B2(new_n755), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n783), .A2(new_n990), .ZN(new_n1015));
  INV_X1    g0815(.A(G322), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1014), .B(new_n1015), .C1(new_n1016), .C2(new_n751), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT48), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n802), .B2(new_n760), .C1(new_n757), .C2(new_n999), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT49), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n767), .A2(new_n753), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n742), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n329), .B1(new_n1024), .B2(G116), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n760), .A2(new_n213), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G159), .A2(new_n752), .B1(new_n763), .B2(new_n376), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n350), .B2(new_n745), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1027), .B(new_n1029), .C1(G50), .C2(new_n755), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n774), .A2(new_n378), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n409), .B(new_n994), .C1(G68), .C2(new_n783), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT112), .Z(new_n1034));
  NAND2_X1  g0834(.A1(new_n1026), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n720), .B1(new_n1035), .B2(new_n727), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n348), .A2(G50), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n475), .B1(new_n1038), .B2(KEYINPUT50), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G68), .B2(G77), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n671), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT111), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n1038), .A2(KEYINPUT50), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1040), .B(new_n1043), .C1(new_n1042), .C2(new_n1041), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1044), .B(new_n731), .C1(new_n236), .C2(new_n475), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(G107), .B2(new_n209), .C1(new_n671), .C2(new_n734), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n728), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n662), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1036), .B(new_n1047), .C1(new_n1048), .C2(new_n788), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n975), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1049), .B1(new_n969), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1013), .A2(new_n1052), .ZN(G393));
  NAND2_X1  g0853(.A1(new_n965), .A2(new_n972), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n1009), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1055), .A2(new_n973), .A3(new_n1012), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n965), .A2(new_n975), .A3(new_n972), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n752), .A2(G317), .B1(G311), .B2(new_n755), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT116), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT52), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G294), .A2(new_n783), .B1(new_n763), .B2(new_n990), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n1016), .B2(new_n745), .C1(new_n760), .C2(new_n999), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(G107), .B2(new_n1024), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n329), .B1(new_n758), .B2(G116), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1060), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT117), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n780), .A2(new_n401), .B1(new_n751), .B2(new_n350), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT51), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n774), .A2(G77), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n805), .A2(G68), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n409), .B(new_n804), .C1(G143), .C2(new_n767), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n376), .A2(new_n783), .B1(new_n763), .B2(G50), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT114), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT115), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1066), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n720), .B1(new_n1077), .B2(new_n727), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n728), .B1(new_n457), .B2(new_n209), .C1(new_n247), .C2(new_n1004), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n953), .A2(new_n726), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1057), .A2(KEYINPUT118), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(KEYINPUT118), .B1(new_n1057), .B2(new_n1081), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1056), .B1(new_n1083), .B2(new_n1084), .ZN(G390));
  AND3_X1   g0885(.A1(new_n903), .A2(KEYINPUT39), .A3(new_n879), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT39), .B1(new_n875), .B2(new_n879), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n724), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1069), .B1(new_n246), .B2(new_n780), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT120), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G283), .A2(new_n752), .B1(new_n763), .B2(G107), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n802), .B2(new_n745), .ZN(new_n1092));
  OR3_X1    g0892(.A1(new_n791), .A2(new_n778), .A3(new_n329), .ZN(new_n1093));
  NOR3_X1   g0893(.A1(new_n1090), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n783), .A2(G97), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n767), .A2(G125), .ZN(new_n1096));
  INV_X1    g0896(.A(G128), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n780), .A2(new_n800), .B1(new_n751), .B2(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT119), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n401), .B2(new_n773), .ZN(new_n1100));
  XOR2_X1   g0900(.A(KEYINPUT54), .B(G143), .Z(new_n1101));
  NAND2_X1  g0901(.A1(new_n783), .A2(new_n1101), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1102), .B1(new_n202), .B2(new_n742), .C1(new_n986), .C2(new_n796), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n760), .A2(new_n350), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT53), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n409), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n1105), .B2(new_n1104), .ZN(new_n1107));
  NOR3_X1   g0907(.A1(new_n1100), .A2(new_n1103), .A3(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1094), .A2(new_n1095), .B1(new_n1096), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1110), .A2(new_n727), .B1(new_n348), .B2(new_n816), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1088), .A2(new_n721), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n317), .A2(new_n660), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n907), .B2(new_n909), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n906), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n687), .B2(new_n886), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n910), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n871), .A2(new_n1118), .A3(new_n1113), .A4(new_n880), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n823), .A2(G330), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n910), .A2(new_n710), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n1115), .A2(new_n1119), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n823), .A2(G330), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1124), .B(new_n909), .C1(new_n846), .C2(new_n851), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1112), .B1(new_n1127), .B2(new_n1050), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n449), .A2(new_n885), .A3(G330), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1129), .A2(new_n915), .A3(new_n638), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n910), .B1(new_n710), .B2(new_n1120), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n908), .B1(new_n1125), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1117), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1124), .B1(new_n846), .B2(new_n851), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1121), .B(new_n1133), .C1(new_n1134), .C2(new_n910), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1130), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1136), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1011), .B1(new_n1127), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1128), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(G378));
  INV_X1    g0941(.A(new_n1130), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1137), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n881), .A2(new_n893), .A3(G330), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n353), .A2(new_n854), .ZN(new_n1145));
  XOR2_X1   g0945(.A(new_n1145), .B(KEYINPUT56), .Z(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n364), .A2(new_n371), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(KEYINPUT55), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1148), .A2(KEYINPUT55), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1147), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1151), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1153), .A2(new_n1149), .A3(new_n1146), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1144), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n881), .A2(new_n1155), .A3(new_n893), .A4(G330), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n913), .A2(KEYINPUT122), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1157), .A2(KEYINPUT122), .A3(new_n913), .A4(new_n1158), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1143), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT57), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1159), .A2(new_n913), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n913), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1168));
  OAI211_X1 g0968(.A(KEYINPUT57), .B(new_n1143), .C1(new_n1166), .C2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1165), .A2(new_n1012), .A3(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1161), .A2(new_n1162), .A3(new_n975), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G125), .A2(new_n752), .B1(new_n783), .B2(G137), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n800), .B2(new_n986), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n805), .A2(new_n1101), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT121), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1173), .B(new_n1175), .C1(G150), .C2(new_n774), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n1097), .B2(new_n780), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT59), .Z(new_n1178));
  AOI21_X1  g0978(.A(G41), .B1(new_n767), .B2(G124), .ZN(new_n1179));
  AOI21_X1  g0979(.A(G33), .B1(new_n1024), .B2(G159), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n202), .B1(new_n292), .B2(G41), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n742), .A2(new_n781), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n378), .B2(new_n783), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(new_n244), .B2(new_n780), .C1(new_n743), .C2(new_n745), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n986), .A2(new_n457), .B1(new_n246), .B2(new_n751), .ZN(new_n1186));
  NOR4_X1   g0986(.A1(new_n1185), .A2(G41), .A3(new_n1027), .A4(new_n1186), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1187), .B(new_n409), .C1(new_n220), .C2(new_n773), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT58), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1181), .A2(new_n1182), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n720), .B1(new_n1190), .B2(new_n727), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1191), .B1(G50), .B2(new_n817), .C1(new_n1155), .C2(new_n725), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1171), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1170), .A2(new_n1193), .ZN(G375));
  OAI221_X1 g0994(.A(new_n409), .B1(new_n213), .B2(new_n742), .C1(new_n986), .C2(new_n246), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n752), .A2(G294), .B1(new_n767), .B2(G303), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n244), .B2(new_n738), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1195), .B(new_n1197), .C1(G283), .C2(new_n755), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1198), .B(new_n1031), .C1(new_n457), .C2(new_n760), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT123), .Z(new_n1200));
  NOR2_X1   g1000(.A1(new_n738), .A2(new_n350), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n751), .A2(new_n800), .B1(new_n745), .B2(new_n1097), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(G159), .C2(new_n805), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n409), .B(new_n1183), .C1(new_n763), .C2(new_n1101), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(new_n202), .C2(new_n773), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G137), .B2(new_n755), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n727), .B1(new_n1200), .B2(new_n1206), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n721), .B(new_n1207), .C1(new_n910), .C2(new_n725), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n220), .B2(new_n816), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1209), .B1(new_n1210), .B2(new_n975), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1132), .A2(new_n1130), .A3(new_n1135), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n951), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1211), .B1(new_n1213), .B2(new_n1136), .ZN(G381));
  NOR2_X1   g1014(.A1(G375), .A2(G378), .ZN(new_n1215));
  INV_X1    g1015(.A(G396), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1013), .A2(new_n1216), .A3(new_n1052), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(G387), .A2(G390), .A3(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(G381), .A2(G384), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1215), .A2(new_n1218), .A3(new_n1219), .ZN(G407));
  NAND2_X1  g1020(.A1(new_n1215), .A2(new_n648), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(G407), .A2(G213), .A3(new_n1221), .ZN(G409));
  NAND3_X1  g1022(.A1(new_n648), .A2(G213), .A3(G2897), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1140), .B1(new_n1170), .B2(new_n1193), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1143), .A2(new_n1161), .A3(new_n951), .A4(new_n1162), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n975), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1140), .A2(new_n1192), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n648), .A2(G213), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1223), .B1(new_n1224), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT60), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1136), .B1(new_n1231), .B2(new_n1212), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1232), .B(new_n1012), .C1(new_n1231), .C2(new_n1212), .ZN(new_n1233));
  AND3_X1   g1033(.A1(new_n1233), .A2(G384), .A3(new_n1211), .ZN(new_n1234));
  AOI21_X1  g1034(.A(G384), .B1(new_n1233), .B2(new_n1211), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1230), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT62), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1236), .B(new_n1223), .C1(new_n1224), .C2(new_n1229), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(G375), .A2(G378), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1229), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1242), .A2(new_n1236), .A3(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(KEYINPUT61), .B1(new_n1244), .B2(KEYINPUT62), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1241), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT124), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1013), .A2(new_n1216), .A3(new_n1052), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1216), .B1(new_n1013), .B2(new_n1052), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1247), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(G393), .A2(G396), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1251), .A2(KEYINPUT124), .A3(new_n1217), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1250), .A2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(G390), .A2(new_n976), .A3(new_n1006), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(G390), .B1(new_n1006), .B2(new_n976), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1253), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1084), .ZN(new_n1258));
  AND2_X1   g1058(.A1(new_n973), .A2(new_n1012), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n1258), .A2(new_n1082), .B1(new_n1259), .B2(new_n1055), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(G387), .A2(new_n1260), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1250), .A2(new_n1252), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT125), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .A4(new_n1254), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1256), .A2(KEYINPUT125), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1257), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1246), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1238), .A2(KEYINPUT63), .A3(new_n1240), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT61), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1257), .A2(new_n1264), .A3(new_n1269), .A4(new_n1265), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT63), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1270), .B1(new_n1271), .B2(new_n1244), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n1268), .A2(new_n1272), .A3(KEYINPUT126), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT126), .B1(new_n1268), .B2(new_n1272), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1267), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT127), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1267), .B(KEYINPUT127), .C1(new_n1273), .C2(new_n1274), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(G405));
  NOR2_X1   g1079(.A1(new_n1215), .A2(new_n1224), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1280), .B(new_n1236), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(new_n1266), .ZN(G402));
endmodule


