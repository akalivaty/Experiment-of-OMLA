

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767;

  INV_X1 U381 ( .A(n564), .ZN(n580) );
  XNOR2_X1 U382 ( .A(n493), .B(n494), .ZN(n752) );
  XNOR2_X1 U383 ( .A(n534), .B(G469), .ZN(n611) );
  NOR2_X1 U384 ( .A1(n670), .A2(n580), .ZN(n579) );
  INV_X2 U385 ( .A(G953), .ZN(n756) );
  NOR2_X1 U386 ( .A1(n618), .A2(n617), .ZN(n708) );
  NOR2_X2 U387 ( .A1(n630), .A2(n629), .ZN(n706) );
  XNOR2_X2 U388 ( .A(G143), .B(G128), .ZN(n535) );
  NOR2_X1 U389 ( .A1(n643), .A2(n608), .ZN(n407) );
  NAND2_X1 U390 ( .A1(n584), .A2(n583), .ZN(n608) );
  XNOR2_X1 U391 ( .A(n560), .B(KEYINPUT35), .ZN(n764) );
  NOR2_X1 U392 ( .A1(n763), .A2(n766), .ZN(n616) );
  XNOR2_X1 U393 ( .A(n407), .B(n366), .ZN(n763) );
  AND2_X1 U394 ( .A1(n396), .A2(n376), .ZN(n380) );
  XNOR2_X1 U395 ( .A(n471), .B(n470), .ZN(n766) );
  NAND2_X1 U396 ( .A1(n473), .A2(n472), .ZN(n471) );
  INV_X1 U397 ( .A(n618), .ZN(n472) );
  INV_X1 U398 ( .A(n673), .ZN(n473) );
  AND2_X1 U399 ( .A1(n606), .A2(n605), .ZN(n626) );
  AND2_X1 U400 ( .A1(n408), .A2(n604), .ZN(n605) );
  NOR2_X1 U401 ( .A1(n611), .A2(n660), .ZN(n601) );
  BUF_X1 U402 ( .A(n567), .Z(n426) );
  XNOR2_X1 U403 ( .A(n558), .B(n557), .ZN(n584) );
  XNOR2_X1 U404 ( .A(n439), .B(G122), .ZN(n539) );
  XNOR2_X1 U405 ( .A(n485), .B(G110), .ZN(n739) );
  XNOR2_X1 U406 ( .A(n427), .B(G146), .ZN(n510) );
  XNOR2_X1 U407 ( .A(KEYINPUT42), .B(KEYINPUT107), .ZN(n470) );
  XNOR2_X1 U408 ( .A(G104), .B(KEYINPUT86), .ZN(n485) );
  XNOR2_X1 U409 ( .A(G107), .B(G116), .ZN(n439) );
  NOR2_X1 U410 ( .A1(n455), .A2(n490), .ZN(n454) );
  XNOR2_X1 U411 ( .A(n510), .B(n509), .ZN(n552) );
  INV_X1 U412 ( .A(KEYINPUT10), .ZN(n509) );
  XNOR2_X1 U413 ( .A(n535), .B(n482), .ZN(n493) );
  INV_X1 U414 ( .A(KEYINPUT4), .ZN(n482) );
  NOR2_X1 U415 ( .A1(G902), .A2(n724), .ZN(n534) );
  NAND2_X1 U416 ( .A1(n447), .A2(n445), .ZN(n564) );
  AND2_X1 U417 ( .A1(n449), .A2(n448), .ZN(n447) );
  AND2_X1 U418 ( .A1(n453), .A2(n359), .ZN(n446) );
  XNOR2_X1 U419 ( .A(n383), .B(n382), .ZN(n381) );
  NOR2_X1 U420 ( .A1(n388), .A2(n767), .ZN(n387) );
  NAND2_X1 U421 ( .A1(n372), .A2(G472), .ZN(n462) );
  NAND2_X1 U422 ( .A1(n372), .A2(G217), .ZN(n476) );
  NOR2_X1 U423 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U424 ( .A1(n492), .A2(n592), .ZN(n475) );
  NOR2_X1 U425 ( .A1(n764), .A2(KEYINPUT44), .ZN(n571) );
  XOR2_X1 U426 ( .A(G101), .B(KEYINPUT66), .Z(n495) );
  XNOR2_X1 U427 ( .A(G131), .B(G134), .ZN(n494) );
  XNOR2_X1 U428 ( .A(n514), .B(n513), .ZN(n515) );
  INV_X1 U429 ( .A(KEYINPUT24), .ZN(n513) );
  XOR2_X1 U430 ( .A(G110), .B(G128), .Z(n516) );
  NAND2_X1 U431 ( .A1(n390), .A2(n389), .ZN(n388) );
  XNOR2_X1 U432 ( .A(n561), .B(KEYINPUT84), .ZN(n389) );
  AND2_X1 U433 ( .A1(n570), .A2(n362), .ZN(n390) );
  NAND2_X1 U434 ( .A1(n429), .A2(n465), .ZN(n645) );
  NOR2_X1 U435 ( .A1(n720), .A2(n466), .ZN(n465) );
  INV_X1 U436 ( .A(n718), .ZN(n466) );
  XOR2_X1 U437 ( .A(G137), .B(G140), .Z(n529) );
  XNOR2_X1 U438 ( .A(n752), .B(G146), .ZN(n528) );
  INV_X1 U439 ( .A(G107), .ZN(n525) );
  INV_X1 U440 ( .A(G125), .ZN(n427) );
  XNOR2_X1 U441 ( .A(n486), .B(n495), .ZN(n531) );
  XNOR2_X1 U442 ( .A(n739), .B(KEYINPUT72), .ZN(n486) );
  XNOR2_X1 U443 ( .A(n479), .B(n478), .ZN(n477) );
  XNOR2_X1 U444 ( .A(n480), .B(KEYINPUT17), .ZN(n479) );
  NAND2_X1 U445 ( .A1(n756), .A2(G224), .ZN(n478) );
  INV_X1 U446 ( .A(n490), .ZN(n458) );
  XNOR2_X1 U447 ( .A(n544), .B(G478), .ZN(n583) );
  XNOR2_X1 U448 ( .A(n522), .B(n521), .ZN(n664) );
  XNOR2_X1 U449 ( .A(n520), .B(KEYINPUT25), .ZN(n521) );
  XNOR2_X1 U450 ( .A(n436), .B(n435), .ZN(n499) );
  XNOR2_X1 U451 ( .A(KEYINPUT3), .B(KEYINPUT71), .ZN(n435) );
  XNOR2_X1 U452 ( .A(n437), .B(G119), .ZN(n436) );
  INV_X1 U453 ( .A(G113), .ZN(n437) );
  NOR2_X1 U454 ( .A1(n687), .A2(n361), .ZN(n394) );
  XNOR2_X1 U455 ( .A(n489), .B(KEYINPUT88), .ZN(n650) );
  AND2_X1 U456 ( .A1(n377), .A2(n627), .ZN(n376) );
  NAND2_X1 U457 ( .A1(n564), .A2(n395), .ZN(n379) );
  BUF_X1 U458 ( .A(n661), .Z(n433) );
  XNOR2_X1 U459 ( .A(n374), .B(n373), .ZN(n568) );
  INV_X1 U460 ( .A(KEYINPUT22), .ZN(n373) );
  NAND2_X1 U461 ( .A1(n564), .A2(n375), .ZN(n374) );
  AND2_X1 U462 ( .A1(n652), .A2(n663), .ZN(n375) );
  INV_X1 U463 ( .A(n457), .ZN(n452) );
  NOR2_X1 U464 ( .A1(n650), .A2(n458), .ZN(n456) );
  XNOR2_X1 U465 ( .A(n403), .B(n613), .ZN(n614) );
  NAND2_X1 U466 ( .A1(n398), .A2(n405), .ZN(n397) );
  NAND2_X1 U467 ( .A1(n399), .A2(n747), .ZN(n398) );
  INV_X1 U468 ( .A(KEYINPUT69), .ZN(n412) );
  INV_X1 U469 ( .A(KEYINPUT18), .ZN(n480) );
  XNOR2_X1 U470 ( .A(n463), .B(KEYINPUT105), .ZN(n655) );
  NAND2_X1 U471 ( .A1(n649), .A2(n650), .ZN(n463) );
  AND2_X1 U472 ( .A1(n441), .A2(n459), .ZN(n440) );
  OR2_X1 U473 ( .A1(n442), .A2(n454), .ZN(n441) );
  XNOR2_X1 U474 ( .A(n497), .B(n496), .ZN(n498) );
  INV_X1 U475 ( .A(KEYINPUT5), .ZN(n496) );
  XNOR2_X1 U476 ( .A(n501), .B(n500), .ZN(n504) );
  NOR2_X1 U477 ( .A1(G953), .A2(G237), .ZN(n502) );
  XNOR2_X1 U478 ( .A(G113), .B(G122), .ZN(n548) );
  XOR2_X1 U479 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n549) );
  XNOR2_X1 U480 ( .A(G104), .B(G143), .ZN(n546) );
  XOR2_X1 U481 ( .A(G131), .B(G140), .Z(n547) );
  XNOR2_X1 U482 ( .A(n552), .B(n432), .ZN(n553) );
  XNOR2_X1 U483 ( .A(KEYINPUT90), .B(KEYINPUT91), .ZN(n432) );
  INV_X1 U484 ( .A(KEYINPUT73), .ZN(n382) );
  NAND2_X1 U485 ( .A1(G234), .A2(G237), .ZN(n481) );
  XNOR2_X1 U486 ( .A(n628), .B(n464), .ZN(n649) );
  INV_X1 U487 ( .A(KEYINPUT38), .ZN(n464) );
  OR2_X1 U488 ( .A1(G902), .A2(G237), .ZN(n488) );
  NOR2_X1 U489 ( .A1(n584), .A2(n582), .ZN(n652) );
  NOR2_X1 U490 ( .A1(n661), .A2(n660), .ZN(n578) );
  XNOR2_X1 U491 ( .A(n602), .B(n409), .ZN(n408) );
  INV_X1 U492 ( .A(KEYINPUT30), .ZN(n409) );
  INV_X1 U493 ( .A(n583), .ZN(n582) );
  XNOR2_X1 U494 ( .A(n645), .B(KEYINPUT82), .ZN(n755) );
  XNOR2_X1 U495 ( .A(n517), .B(n428), .ZN(n646) );
  XNOR2_X1 U496 ( .A(n518), .B(n516), .ZN(n428) );
  XNOR2_X1 U497 ( .A(G902), .B(KEYINPUT15), .ZN(n644) );
  NOR2_X1 U498 ( .A1(n645), .A2(n405), .ZN(n404) );
  XNOR2_X1 U499 ( .A(n533), .B(n532), .ZN(n724) );
  XNOR2_X1 U500 ( .A(n528), .B(n527), .ZN(n533) );
  XNOR2_X1 U501 ( .A(n371), .B(n487), .ZN(n722) );
  XNOR2_X1 U502 ( .A(n740), .B(n531), .ZN(n371) );
  AND2_X1 U503 ( .A1(n707), .A2(n430), .ZN(n631) );
  INV_X1 U504 ( .A(n612), .ZN(n431) );
  XNOR2_X1 U505 ( .A(n631), .B(n411), .ZN(n632) );
  INV_X1 U506 ( .A(KEYINPUT108), .ZN(n411) );
  BUF_X1 U507 ( .A(n628), .Z(n410) );
  XNOR2_X1 U508 ( .A(n438), .B(n499), .ZN(n740) );
  XNOR2_X1 U509 ( .A(n539), .B(KEYINPUT16), .ZN(n438) );
  XNOR2_X1 U510 ( .A(n542), .B(n413), .ZN(n736) );
  XNOR2_X1 U511 ( .A(n541), .B(n543), .ZN(n413) );
  INV_X1 U512 ( .A(KEYINPUT120), .ZN(n391) );
  NAND2_X1 U513 ( .A1(n393), .A2(n360), .ZN(n392) );
  NAND2_X1 U514 ( .A1(n380), .A2(n378), .ZN(n560) );
  NAND2_X1 U515 ( .A1(n565), .A2(n568), .ZN(n566) );
  NAND2_X1 U516 ( .A1(n452), .A2(n363), .ZN(n617) );
  XNOR2_X1 U517 ( .A(KEYINPUT99), .B(n608), .ZN(n707) );
  XNOR2_X1 U518 ( .A(n577), .B(KEYINPUT96), .ZN(n767) );
  NOR2_X1 U519 ( .A1(n576), .A2(n575), .ZN(n577) );
  OR2_X1 U520 ( .A1(n574), .A2(n573), .ZN(n576) );
  NAND2_X1 U521 ( .A1(n406), .A2(n461), .ZN(n460) );
  XNOR2_X1 U522 ( .A(n462), .B(n691), .ZN(n406) );
  XNOR2_X1 U523 ( .A(n690), .B(KEYINPUT62), .ZN(n691) );
  INV_X1 U524 ( .A(KEYINPUT124), .ZN(n416) );
  XNOR2_X1 U525 ( .A(n476), .B(n367), .ZN(n421) );
  INV_X1 U526 ( .A(KEYINPUT60), .ZN(n424) );
  INV_X1 U527 ( .A(KEYINPUT56), .ZN(n418) );
  AND2_X1 U528 ( .A1(n451), .A2(KEYINPUT0), .ZN(n359) );
  XOR2_X1 U529 ( .A(n683), .B(KEYINPUT119), .Z(n360) );
  AND2_X1 U530 ( .A1(n755), .A2(n685), .ZN(n361) );
  XNOR2_X1 U531 ( .A(n609), .B(n610), .ZN(n673) );
  XOR2_X1 U532 ( .A(n586), .B(KEYINPUT95), .Z(n362) );
  AND2_X1 U533 ( .A1(n453), .A2(n450), .ZN(n363) );
  AND2_X1 U534 ( .A1(n488), .A2(G210), .ZN(n364) );
  XNOR2_X1 U535 ( .A(KEYINPUT97), .B(KEYINPUT33), .ZN(n365) );
  XOR2_X1 U536 ( .A(n600), .B(KEYINPUT104), .Z(n366) );
  INV_X1 U537 ( .A(KEYINPUT0), .ZN(n459) );
  XOR2_X1 U538 ( .A(n647), .B(KEYINPUT123), .Z(n367) );
  XOR2_X1 U539 ( .A(n723), .B(n721), .Z(n368) );
  NOR2_X1 U540 ( .A1(G952), .A2(n756), .ZN(n738) );
  INV_X1 U541 ( .A(n738), .ZN(n461) );
  XOR2_X1 U542 ( .A(n688), .B(KEYINPUT121), .Z(n369) );
  INV_X1 U543 ( .A(KEYINPUT2), .ZN(n405) );
  INV_X1 U544 ( .A(n685), .ZN(n422) );
  XNOR2_X2 U545 ( .A(n370), .B(n364), .ZN(n628) );
  NAND2_X1 U546 ( .A1(n722), .A2(n644), .ZN(n370) );
  NAND2_X1 U547 ( .A1(n372), .A2(G475), .ZN(n733) );
  NAND2_X1 U548 ( .A1(n372), .A2(G210), .ZN(n474) );
  NAND2_X1 U549 ( .A1(n372), .A2(G469), .ZN(n727) );
  NAND2_X1 U550 ( .A1(n372), .A2(G478), .ZN(n735) );
  AND2_X2 U551 ( .A1(n400), .A2(n397), .ZN(n372) );
  NAND2_X1 U552 ( .A1(n580), .A2(KEYINPUT34), .ZN(n377) );
  OR2_X1 U553 ( .A1(n648), .A2(n379), .ZN(n378) );
  XNOR2_X2 U554 ( .A(n414), .B(n365), .ZN(n648) );
  NAND2_X1 U555 ( .A1(n387), .A2(n381), .ZN(n587) );
  NAND2_X1 U556 ( .A1(n385), .A2(n384), .ZN(n383) );
  INV_X1 U557 ( .A(n572), .ZN(n384) );
  XNOR2_X1 U558 ( .A(n571), .B(n386), .ZN(n385) );
  INV_X1 U559 ( .A(KEYINPUT67), .ZN(n386) );
  XNOR2_X1 U560 ( .A(n392), .B(n391), .ZN(n423) );
  NAND2_X1 U561 ( .A1(n686), .A2(n394), .ZN(n393) );
  INV_X1 U562 ( .A(KEYINPUT34), .ZN(n395) );
  NAND2_X1 U563 ( .A1(n648), .A2(KEYINPUT34), .ZN(n396) );
  INV_X1 U564 ( .A(n755), .ZN(n399) );
  NOR2_X1 U565 ( .A1(n687), .A2(n644), .ZN(n400) );
  AND2_X2 U566 ( .A1(n747), .A2(n404), .ZN(n687) );
  XNOR2_X2 U567 ( .A(n587), .B(KEYINPUT45), .ZN(n747) );
  NAND2_X1 U568 ( .A1(n626), .A2(n649), .ZN(n402) );
  XNOR2_X1 U569 ( .A(n402), .B(n607), .ZN(n643) );
  XNOR2_X1 U570 ( .A(n401), .B(n369), .ZN(G75) );
  NAND2_X1 U571 ( .A1(n423), .A2(n756), .ZN(n401) );
  XNOR2_X1 U572 ( .A(n616), .B(KEYINPUT46), .ZN(n469) );
  NAND2_X1 U573 ( .A1(n578), .A2(n575), .ZN(n414) );
  XNOR2_X1 U574 ( .A(n640), .B(n412), .ZN(n468) );
  NAND2_X1 U575 ( .A1(n426), .A2(n612), .ZN(n403) );
  NAND2_X1 U576 ( .A1(n421), .A2(n461), .ZN(n417) );
  XNOR2_X1 U577 ( .A(n733), .B(n734), .ZN(n434) );
  NAND2_X1 U578 ( .A1(n446), .A2(n452), .ZN(n445) );
  XNOR2_X1 U579 ( .A(n467), .B(n641), .ZN(n429) );
  XNOR2_X1 U580 ( .A(n567), .B(KEYINPUT6), .ZN(n596) );
  XNOR2_X1 U581 ( .A(n528), .B(n498), .ZN(n506) );
  BUF_X1 U582 ( .A(n755), .Z(n415) );
  XNOR2_X1 U583 ( .A(n417), .B(n416), .ZN(G66) );
  XNOR2_X1 U584 ( .A(n611), .B(KEYINPUT1), .ZN(n661) );
  XNOR2_X1 U585 ( .A(n419), .B(n418), .ZN(G51) );
  NAND2_X1 U586 ( .A1(n420), .A2(n461), .ZN(n419) );
  XNOR2_X1 U587 ( .A(n474), .B(n368), .ZN(n420) );
  NAND2_X1 U588 ( .A1(n469), .A2(n468), .ZN(n467) );
  NOR2_X1 U589 ( .A1(n747), .A2(n422), .ZN(n684) );
  XNOR2_X1 U590 ( .A(n425), .B(n424), .ZN(G60) );
  NAND2_X1 U591 ( .A1(n434), .A2(n461), .ZN(n425) );
  NOR2_X1 U592 ( .A1(n431), .A2(n596), .ZN(n430) );
  NAND2_X1 U593 ( .A1(n628), .A2(n454), .ZN(n453) );
  NAND2_X1 U594 ( .A1(n443), .A2(n440), .ZN(n448) );
  INV_X1 U595 ( .A(n451), .ZN(n442) );
  NAND2_X1 U596 ( .A1(n444), .A2(n451), .ZN(n443) );
  INV_X1 U597 ( .A(n628), .ZN(n444) );
  NAND2_X1 U598 ( .A1(n457), .A2(n459), .ZN(n449) );
  INV_X1 U599 ( .A(n456), .ZN(n450) );
  NOR2_X1 U600 ( .A1(n456), .A2(n475), .ZN(n451) );
  NAND2_X1 U601 ( .A1(n410), .A2(n650), .ZN(n633) );
  INV_X1 U602 ( .A(n650), .ZN(n455) );
  NOR2_X1 U603 ( .A1(n628), .A2(n458), .ZN(n457) );
  XNOR2_X1 U604 ( .A(n460), .B(KEYINPUT63), .ZN(G57) );
  NOR2_X1 U605 ( .A1(G902), .A2(n730), .ZN(n557) );
  XNOR2_X1 U606 ( .A(n493), .B(n477), .ZN(n484) );
  INV_X1 U607 ( .A(KEYINPUT74), .ZN(n500) );
  INV_X1 U608 ( .A(KEYINPUT48), .ZN(n641) );
  XNOR2_X1 U609 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U610 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U611 ( .A(n506), .B(n505), .ZN(n689) );
  XNOR2_X1 U612 ( .A(n531), .B(n530), .ZN(n532) );
  INV_X1 U613 ( .A(n603), .ZN(n604) );
  XNOR2_X1 U614 ( .A(n552), .B(n529), .ZN(n754) );
  XNOR2_X1 U615 ( .A(KEYINPUT83), .B(KEYINPUT39), .ZN(n607) );
  INV_X1 U616 ( .A(KEYINPUT53), .ZN(n688) );
  XOR2_X1 U617 ( .A(KEYINPUT14), .B(n481), .Z(n679) );
  XNOR2_X1 U618 ( .A(n510), .B(KEYINPUT87), .ZN(n483) );
  XNOR2_X1 U619 ( .A(n484), .B(n483), .ZN(n487) );
  NAND2_X1 U620 ( .A1(n488), .A2(G214), .ZN(n489) );
  XNOR2_X1 U621 ( .A(KEYINPUT19), .B(KEYINPUT65), .ZN(n490) );
  NAND2_X1 U622 ( .A1(G952), .A2(n756), .ZN(n590) );
  NOR2_X1 U623 ( .A1(G898), .A2(n756), .ZN(n742) );
  NAND2_X1 U624 ( .A1(G902), .A2(n742), .ZN(n491) );
  NAND2_X1 U625 ( .A1(n590), .A2(n491), .ZN(n492) );
  XNOR2_X1 U626 ( .A(n495), .B(G137), .ZN(n497) );
  XNOR2_X1 U627 ( .A(n499), .B(G116), .ZN(n501) );
  XOR2_X1 U628 ( .A(KEYINPUT75), .B(n502), .Z(n545) );
  NAND2_X1 U629 ( .A1(n545), .A2(G210), .ZN(n503) );
  NOR2_X1 U630 ( .A1(G902), .A2(n689), .ZN(n508) );
  XNOR2_X1 U631 ( .A(KEYINPUT89), .B(G472), .ZN(n507) );
  XNOR2_X1 U632 ( .A(n508), .B(n507), .ZN(n567) );
  INV_X1 U633 ( .A(n596), .ZN(n575) );
  XOR2_X1 U634 ( .A(KEYINPUT80), .B(KEYINPUT8), .Z(n512) );
  NAND2_X1 U635 ( .A1(G234), .A2(n756), .ZN(n511) );
  XNOR2_X1 U636 ( .A(n512), .B(n511), .ZN(n540) );
  NAND2_X1 U637 ( .A1(G221), .A2(n540), .ZN(n514) );
  XNOR2_X1 U638 ( .A(n754), .B(n515), .ZN(n517) );
  XOR2_X1 U639 ( .A(G119), .B(KEYINPUT23), .Z(n518) );
  NOR2_X1 U640 ( .A1(n646), .A2(G902), .ZN(n522) );
  NAND2_X1 U641 ( .A1(G234), .A2(n644), .ZN(n519) );
  XNOR2_X1 U642 ( .A(KEYINPUT20), .B(n519), .ZN(n523) );
  NAND2_X1 U643 ( .A1(n523), .A2(G217), .ZN(n520) );
  NAND2_X1 U644 ( .A1(n523), .A2(G221), .ZN(n524) );
  XNOR2_X1 U645 ( .A(n524), .B(KEYINPUT21), .ZN(n593) );
  INV_X1 U646 ( .A(n593), .ZN(n663) );
  NAND2_X1 U647 ( .A1(n664), .A2(n663), .ZN(n660) );
  NAND2_X1 U648 ( .A1(G227), .A2(n756), .ZN(n526) );
  INV_X1 U649 ( .A(n529), .ZN(n530) );
  XOR2_X1 U650 ( .A(n535), .B(KEYINPUT7), .Z(n543) );
  XOR2_X1 U651 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n537) );
  XNOR2_X1 U652 ( .A(G134), .B(KEYINPUT9), .ZN(n536) );
  XNOR2_X1 U653 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U654 ( .A(n539), .B(n538), .Z(n542) );
  NAND2_X1 U655 ( .A1(G217), .A2(n540), .ZN(n541) );
  NOR2_X1 U656 ( .A1(G902), .A2(n736), .ZN(n544) );
  XNOR2_X1 U657 ( .A(KEYINPUT13), .B(G475), .ZN(n558) );
  NAND2_X1 U658 ( .A1(n545), .A2(G214), .ZN(n556) );
  XNOR2_X1 U659 ( .A(n547), .B(n546), .ZN(n551) );
  XNOR2_X1 U660 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U661 ( .A(n551), .B(n550), .ZN(n554) );
  XNOR2_X1 U662 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U663 ( .A(n556), .B(n555), .ZN(n730) );
  NAND2_X1 U664 ( .A1(n582), .A2(n584), .ZN(n559) );
  XOR2_X1 U665 ( .A(KEYINPUT98), .B(n559), .Z(n627) );
  NAND2_X1 U666 ( .A1(n764), .A2(KEYINPUT44), .ZN(n561) );
  INV_X1 U667 ( .A(n664), .ZN(n573) );
  NAND2_X1 U668 ( .A1(n573), .A2(n596), .ZN(n562) );
  NOR2_X1 U669 ( .A1(n433), .A2(n562), .ZN(n563) );
  XNOR2_X1 U670 ( .A(n563), .B(KEYINPUT76), .ZN(n565) );
  XNOR2_X1 U671 ( .A(KEYINPUT32), .B(n566), .ZN(n765) );
  NAND2_X1 U672 ( .A1(n568), .A2(n433), .ZN(n574) );
  NOR2_X1 U673 ( .A1(n426), .A2(n574), .ZN(n569) );
  NAND2_X1 U674 ( .A1(n573), .A2(n569), .ZN(n699) );
  NAND2_X1 U675 ( .A1(n765), .A2(n699), .ZN(n572) );
  NAND2_X1 U676 ( .A1(n572), .A2(KEYINPUT44), .ZN(n570) );
  NAND2_X1 U677 ( .A1(n426), .A2(n578), .ZN(n670) );
  XNOR2_X1 U678 ( .A(n579), .B(KEYINPUT31), .ZN(n713) );
  NOR2_X1 U679 ( .A1(n426), .A2(n580), .ZN(n581) );
  NAND2_X1 U680 ( .A1(n601), .A2(n581), .ZN(n695) );
  NAND2_X1 U681 ( .A1(n713), .A2(n695), .ZN(n585) );
  NOR2_X1 U682 ( .A1(n584), .A2(n583), .ZN(n701) );
  XOR2_X1 U683 ( .A(KEYINPUT94), .B(n701), .Z(n642) );
  NAND2_X1 U684 ( .A1(n642), .A2(n608), .ZN(n654) );
  XNOR2_X1 U685 ( .A(KEYINPUT78), .B(n654), .ZN(n620) );
  NAND2_X1 U686 ( .A1(n585), .A2(n620), .ZN(n586) );
  INV_X1 U687 ( .A(n433), .ZN(n635) );
  INV_X1 U688 ( .A(n679), .ZN(n592) );
  NOR2_X1 U689 ( .A1(G900), .A2(n756), .ZN(n588) );
  NAND2_X1 U690 ( .A1(G902), .A2(n588), .ZN(n589) );
  NAND2_X1 U691 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U692 ( .A1(n592), .A2(n591), .ZN(n603) );
  NOR2_X1 U693 ( .A1(n593), .A2(n603), .ZN(n594) );
  XOR2_X1 U694 ( .A(KEYINPUT70), .B(n594), .Z(n595) );
  NOR2_X1 U695 ( .A1(n664), .A2(n595), .ZN(n612) );
  NAND2_X1 U696 ( .A1(n650), .A2(n631), .ZN(n597) );
  NOR2_X1 U697 ( .A1(n635), .A2(n597), .ZN(n598) );
  XNOR2_X1 U698 ( .A(n598), .B(KEYINPUT43), .ZN(n599) );
  NOR2_X1 U699 ( .A1(n410), .A2(n599), .ZN(n720) );
  XNOR2_X1 U700 ( .A(KEYINPUT103), .B(KEYINPUT40), .ZN(n600) );
  XNOR2_X1 U701 ( .A(n601), .B(KEYINPUT100), .ZN(n606) );
  NAND2_X1 U702 ( .A1(n567), .A2(n650), .ZN(n602) );
  XOR2_X1 U703 ( .A(KEYINPUT106), .B(KEYINPUT41), .Z(n610) );
  NAND2_X1 U704 ( .A1(n655), .A2(n652), .ZN(n609) );
  XNOR2_X1 U705 ( .A(KEYINPUT101), .B(n611), .ZN(n615) );
  XOR2_X1 U706 ( .A(KEYINPUT28), .B(KEYINPUT102), .Z(n613) );
  NAND2_X1 U707 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U708 ( .A1(n654), .A2(n708), .ZN(n619) );
  NAND2_X1 U709 ( .A1(n619), .A2(KEYINPUT47), .ZN(n625) );
  INV_X1 U710 ( .A(n620), .ZN(n622) );
  XNOR2_X1 U711 ( .A(KEYINPUT68), .B(KEYINPUT47), .ZN(n621) );
  NOR2_X1 U712 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U713 ( .A1(n623), .A2(n708), .ZN(n624) );
  NAND2_X1 U714 ( .A1(n625), .A2(n624), .ZN(n639) );
  INV_X1 U715 ( .A(n626), .ZN(n630) );
  NAND2_X1 U716 ( .A1(n410), .A2(n627), .ZN(n629) );
  XNOR2_X1 U717 ( .A(n706), .B(KEYINPUT79), .ZN(n637) );
  NOR2_X1 U718 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U719 ( .A(n634), .B(KEYINPUT36), .ZN(n636) );
  NAND2_X1 U720 ( .A1(n636), .A2(n635), .ZN(n717) );
  NAND2_X1 U721 ( .A1(n637), .A2(n717), .ZN(n638) );
  OR2_X1 U722 ( .A1(n643), .A2(n642), .ZN(n718) );
  INV_X1 U723 ( .A(n646), .ZN(n647) );
  NOR2_X1 U724 ( .A1(n673), .A2(n648), .ZN(n682) );
  INV_X1 U725 ( .A(n648), .ZN(n659) );
  OR2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U727 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U728 ( .A(n653), .B(KEYINPUT118), .ZN(n657) );
  NAND2_X1 U729 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U730 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U731 ( .A1(n659), .A2(n658), .ZN(n676) );
  NAND2_X1 U732 ( .A1(n433), .A2(n660), .ZN(n662) );
  XNOR2_X1 U733 ( .A(n662), .B(KEYINPUT50), .ZN(n669) );
  NOR2_X1 U734 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U735 ( .A(KEYINPUT49), .B(n665), .Z(n666) );
  NOR2_X1 U736 ( .A1(n426), .A2(n666), .ZN(n667) );
  XOR2_X1 U737 ( .A(KEYINPUT117), .B(n667), .Z(n668) );
  NAND2_X1 U738 ( .A1(n669), .A2(n668), .ZN(n671) );
  NAND2_X1 U739 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U740 ( .A(KEYINPUT51), .B(n672), .Z(n674) );
  NAND2_X1 U741 ( .A1(n674), .A2(n473), .ZN(n675) );
  NAND2_X1 U742 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U743 ( .A(KEYINPUT52), .B(n677), .ZN(n678) );
  NAND2_X1 U744 ( .A1(n678), .A2(G952), .ZN(n680) );
  NOR2_X1 U745 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U746 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U747 ( .A(KEYINPUT2), .B(KEYINPUT77), .ZN(n685) );
  XNOR2_X1 U748 ( .A(n684), .B(KEYINPUT81), .ZN(n686) );
  XNOR2_X1 U749 ( .A(n689), .B(KEYINPUT109), .ZN(n690) );
  INV_X1 U750 ( .A(n707), .ZN(n710) );
  NOR2_X1 U751 ( .A1(n710), .A2(n695), .ZN(n693) );
  XNOR2_X1 U752 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n692) );
  XNOR2_X1 U753 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U754 ( .A(G104), .B(n694), .ZN(G6) );
  INV_X1 U755 ( .A(n701), .ZN(n714) );
  NOR2_X1 U756 ( .A1(n714), .A2(n695), .ZN(n697) );
  XNOR2_X1 U757 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n696) );
  XNOR2_X1 U758 ( .A(n697), .B(n696), .ZN(n698) );
  XNOR2_X1 U759 ( .A(G107), .B(n698), .ZN(G9) );
  XNOR2_X1 U760 ( .A(G110), .B(KEYINPUT112), .ZN(n700) );
  XNOR2_X1 U761 ( .A(n700), .B(n699), .ZN(G12) );
  XOR2_X1 U762 ( .A(KEYINPUT29), .B(KEYINPUT114), .Z(n703) );
  NAND2_X1 U763 ( .A1(n708), .A2(n701), .ZN(n702) );
  XNOR2_X1 U764 ( .A(n703), .B(n702), .ZN(n705) );
  XOR2_X1 U765 ( .A(G128), .B(KEYINPUT113), .Z(n704) );
  XNOR2_X1 U766 ( .A(n705), .B(n704), .ZN(G30) );
  XOR2_X1 U767 ( .A(G143), .B(n706), .Z(G45) );
  NAND2_X1 U768 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U769 ( .A(n709), .B(G146), .ZN(G48) );
  NOR2_X1 U770 ( .A1(n710), .A2(n713), .ZN(n712) );
  XNOR2_X1 U771 ( .A(G113), .B(KEYINPUT115), .ZN(n711) );
  XNOR2_X1 U772 ( .A(n712), .B(n711), .ZN(G15) );
  NOR2_X1 U773 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U774 ( .A(G116), .B(n715), .Z(G18) );
  XOR2_X1 U775 ( .A(G125), .B(KEYINPUT37), .Z(n716) );
  XNOR2_X1 U776 ( .A(n717), .B(n716), .ZN(G27) );
  XNOR2_X1 U777 ( .A(G134), .B(KEYINPUT116), .ZN(n719) );
  XNOR2_X1 U778 ( .A(n719), .B(n718), .ZN(G36) );
  XOR2_X1 U779 ( .A(G140), .B(n720), .Z(G42) );
  XOR2_X1 U780 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n721) );
  INV_X1 U781 ( .A(n722), .ZN(n723) );
  XNOR2_X1 U782 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n726) );
  XNOR2_X1 U783 ( .A(n724), .B(KEYINPUT57), .ZN(n725) );
  XNOR2_X1 U784 ( .A(n726), .B(n725), .ZN(n728) );
  XOR2_X1 U785 ( .A(n728), .B(n727), .Z(n729) );
  NOR2_X1 U786 ( .A1(n738), .A2(n729), .ZN(G54) );
  XOR2_X1 U787 ( .A(KEYINPUT59), .B(KEYINPUT64), .Z(n732) );
  XNOR2_X1 U788 ( .A(n730), .B(KEYINPUT85), .ZN(n731) );
  XNOR2_X1 U789 ( .A(n732), .B(n731), .ZN(n734) );
  XNOR2_X1 U790 ( .A(n736), .B(n735), .ZN(n737) );
  NOR2_X1 U791 ( .A1(n738), .A2(n737), .ZN(G63) );
  XNOR2_X1 U792 ( .A(n739), .B(G101), .ZN(n741) );
  XNOR2_X1 U793 ( .A(n741), .B(n740), .ZN(n743) );
  NOR2_X1 U794 ( .A1(n743), .A2(n742), .ZN(n751) );
  XOR2_X1 U795 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n745) );
  NAND2_X1 U796 ( .A1(G224), .A2(G953), .ZN(n744) );
  XNOR2_X1 U797 ( .A(n745), .B(n744), .ZN(n746) );
  NAND2_X1 U798 ( .A1(n746), .A2(G898), .ZN(n749) );
  NAND2_X1 U799 ( .A1(n747), .A2(n756), .ZN(n748) );
  NAND2_X1 U800 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U801 ( .A(n751), .B(n750), .ZN(G69) );
  XOR2_X1 U802 ( .A(KEYINPUT126), .B(n752), .Z(n753) );
  XNOR2_X1 U803 ( .A(n754), .B(n753), .ZN(n758) );
  XNOR2_X1 U804 ( .A(n758), .B(n415), .ZN(n757) );
  NAND2_X1 U805 ( .A1(n757), .A2(n756), .ZN(n762) );
  XNOR2_X1 U806 ( .A(G227), .B(n758), .ZN(n759) );
  NAND2_X1 U807 ( .A1(n759), .A2(G900), .ZN(n760) );
  NAND2_X1 U808 ( .A1(G953), .A2(n760), .ZN(n761) );
  NAND2_X1 U809 ( .A1(n762), .A2(n761), .ZN(G72) );
  XOR2_X1 U810 ( .A(n763), .B(G131), .Z(G33) );
  XOR2_X1 U811 ( .A(n764), .B(G122), .Z(G24) );
  XNOR2_X1 U812 ( .A(G119), .B(n765), .ZN(G21) );
  XOR2_X1 U813 ( .A(n766), .B(G137), .Z(G39) );
  XOR2_X1 U814 ( .A(n767), .B(G101), .Z(G3) );
endmodule

