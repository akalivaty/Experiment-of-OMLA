//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 0 1 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985;
  XOR2_X1   g000(.A(G134gat), .B(G162gat), .Z(new_n202));
  AOI21_X1  g001(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT99), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G29gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n207), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n208));
  XOR2_X1   g007(.A(KEYINPUT14), .B(G29gat), .Z(new_n209));
  OAI21_X1  g008(.A(new_n208), .B1(new_n209), .B2(G36gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(G43gat), .B(G50gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT15), .ZN(new_n212));
  OR3_X1    g011(.A1(new_n210), .A2(KEYINPUT90), .A3(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT90), .B1(new_n210), .B2(new_n212), .ZN(new_n214));
  XOR2_X1   g013(.A(new_n211), .B(KEYINPUT15), .Z(new_n215));
  AOI22_X1  g014(.A1(new_n213), .A2(new_n214), .B1(new_n210), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT98), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(G85gat), .A3(G92gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT7), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G99gat), .A2(G106gat), .ZN(new_n222));
  INV_X1    g021(.A(G85gat), .ZN(new_n223));
  INV_X1    g022(.A(G92gat), .ZN(new_n224));
  AOI22_X1  g023(.A1(KEYINPUT8), .A2(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n218), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n221), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  XOR2_X1   g026(.A(G99gat), .B(G106gat), .Z(new_n228));
  XNOR2_X1  g027(.A(new_n227), .B(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n217), .B1(KEYINPUT17), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT17), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n232), .A3(new_n229), .ZN(new_n233));
  NAND3_X1  g032(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  XOR2_X1   g034(.A(G190gat), .B(G218gat), .Z(new_n236));
  OR2_X1    g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n236), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n206), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT99), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n204), .A2(new_n240), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n237), .A2(new_n238), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n239), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT9), .ZN(new_n245));
  INV_X1    g044(.A(G57gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G64gat), .ZN(new_n247));
  INV_X1    g046(.A(G64gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(G57gat), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n245), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  OR2_X1    g049(.A1(G71gat), .A2(G78gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(G71gat), .A2(G78gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OR3_X1    g052(.A1(new_n250), .A2(KEYINPUT93), .A3(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT93), .B1(new_n250), .B2(new_n253), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n252), .B1(new_n251), .B2(new_n245), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT94), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n247), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n246), .A2(KEYINPUT94), .A3(G64gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(new_n249), .A3(new_n259), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n254), .A2(new_n255), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n261), .A2(KEYINPUT21), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(KEYINPUT95), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(KEYINPUT96), .ZN(new_n264));
  XOR2_X1   g063(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  XOR2_X1   g065(.A(G183gat), .B(G211gat), .Z(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  OR2_X1    g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n266), .A2(new_n268), .ZN(new_n270));
  XNOR2_X1  g069(.A(G15gat), .B(G22gat), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT16), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n271), .B1(new_n272), .B2(G1gat), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n273), .B1(G1gat), .B2(new_n271), .ZN(new_n274));
  INV_X1    g073(.A(G8gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n261), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT21), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT97), .ZN(new_n280));
  XNOR2_X1  g079(.A(G127gat), .B(G155gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(G231gat), .A2(G233gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  XOR2_X1   g082(.A(new_n280), .B(new_n283), .Z(new_n284));
  AND3_X1   g083(.A1(new_n269), .A2(new_n270), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n284), .B1(new_n269), .B2(new_n270), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n244), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G230gat), .A2(G233gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT100), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n228), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n227), .B(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n261), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT101), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n229), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT10), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT101), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n261), .A2(new_n292), .A3(new_n297), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n294), .A2(new_n295), .A3(new_n296), .A4(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n230), .A2(KEYINPUT10), .A3(new_n261), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n289), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n294), .A2(new_n295), .A3(new_n298), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(new_n289), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G120gat), .B(G148gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(G176gat), .B(G204gat), .ZN(new_n307));
  XOR2_X1   g106(.A(new_n306), .B(new_n307), .Z(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n302), .A2(new_n304), .A3(new_n308), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT102), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n310), .A2(KEYINPUT102), .A3(new_n311), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n287), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G113gat), .B(G141gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G169gat), .B(G197gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n320), .B(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n322), .B(KEYINPUT12), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT18), .ZN(new_n324));
  OAI21_X1  g123(.A(KEYINPUT91), .B1(new_n216), .B2(KEYINPUT17), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT91), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n232), .B1(new_n276), .B2(new_n326), .ZN(new_n327));
  AOI22_X1  g126(.A1(new_n325), .A2(new_n276), .B1(new_n327), .B2(new_n216), .ZN(new_n328));
  NAND2_X1  g127(.A1(G229gat), .A2(G233gat), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n324), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT92), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n323), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NOR3_X1   g133(.A1(new_n328), .A2(new_n324), .A3(new_n330), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n216), .B(new_n276), .ZN(new_n337));
  XOR2_X1   g136(.A(new_n329), .B(KEYINPUT13), .Z(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n334), .A2(new_n331), .A3(new_n336), .A4(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n331), .A2(new_n339), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n333), .B1(new_n335), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n317), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT86), .ZN(new_n345));
  NOR2_X1   g144(.A1(G127gat), .A2(G134gat), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT70), .B(G134gat), .ZN(new_n348));
  INV_X1    g147(.A(G127gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(G120gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G113gat), .ZN(new_n352));
  INV_X1    g151(.A(G113gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(G120gat), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT1), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT71), .B1(new_n350), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n355), .ZN(new_n357));
  INV_X1    g156(.A(G134gat), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n358), .A2(KEYINPUT70), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(KEYINPUT70), .ZN(new_n360));
  OAI21_X1  g159(.A(G127gat), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT71), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n357), .A2(new_n361), .A3(new_n362), .A4(new_n347), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT1), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n349), .A2(new_n358), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT72), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n366), .B1(new_n351), .B2(G113gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(new_n352), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n354), .A2(new_n366), .ZN(new_n369));
  OAI221_X1 g168(.A(new_n364), .B1(new_n346), .B2(new_n365), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n356), .A2(new_n363), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT78), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT4), .ZN(new_n373));
  AND2_X1   g172(.A1(G155gat), .A2(G162gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(G155gat), .A2(G162gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G141gat), .B(G148gat), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT2), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n378), .B1(G155gat), .B2(G162gat), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n376), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(G141gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(G148gat), .ZN(new_n382));
  INV_X1    g181(.A(G148gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(G141gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G155gat), .B(G162gat), .ZN(new_n386));
  INV_X1    g185(.A(G155gat), .ZN(new_n387));
  INV_X1    g186(.A(G162gat), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT2), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n385), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n380), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n371), .A2(new_n372), .A3(new_n373), .A4(new_n391), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n391), .A2(new_n356), .A3(new_n363), .A4(new_n370), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT78), .B1(new_n393), .B2(KEYINPUT4), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(KEYINPUT4), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n392), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(G225gat), .A2(G233gat), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n380), .A2(new_n390), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT3), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n399), .B(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n356), .A2(new_n363), .A3(new_n370), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n398), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n396), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT5), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n402), .A2(new_n399), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n393), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n405), .B1(new_n407), .B2(new_n398), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G1gat), .B(G29gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(KEYINPUT0), .ZN(new_n411));
  XNOR2_X1  g210(.A(G57gat), .B(G85gat), .ZN(new_n412));
  XOR2_X1   g211(.A(new_n411), .B(new_n412), .Z(new_n413));
  NAND3_X1  g212(.A1(new_n371), .A2(new_n373), .A3(new_n391), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n395), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n401), .A2(new_n402), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n398), .A2(KEYINPUT5), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n409), .A2(new_n413), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT6), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n413), .B1(new_n409), .B2(new_n418), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n345), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(KEYINPUT6), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n418), .ZN(new_n425));
  INV_X1    g224(.A(new_n413), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n427), .A2(KEYINPUT86), .A3(new_n420), .A4(new_n419), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n423), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G78gat), .B(G106gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(KEYINPUT31), .B(G50gat), .ZN(new_n431));
  XOR2_X1   g230(.A(new_n430), .B(new_n431), .Z(new_n432));
  NAND2_X1  g231(.A1(G211gat), .A2(G218gat), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT22), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g234(.A1(G197gat), .A2(G204gat), .ZN(new_n436));
  AND2_X1   g235(.A1(G197gat), .A2(G204gat), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  XOR2_X1   g237(.A(G211gat), .B(G218gat), .Z(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G211gat), .B(G218gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(G197gat), .B(G204gat), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(new_n442), .A3(new_n435), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT29), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n400), .B1(new_n444), .B2(KEYINPUT80), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT80), .ZN(new_n446));
  AOI211_X1 g245(.A(new_n446), .B(KEYINPUT29), .C1(new_n440), .C2(new_n443), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n399), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n440), .A2(new_n443), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n380), .A2(new_n390), .A3(new_n400), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT29), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n448), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(G228gat), .ZN(new_n455));
  INV_X1    g254(.A(G233gat), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n400), .B1(new_n444), .B2(KEYINPUT81), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n449), .A2(KEYINPUT81), .A3(new_n451), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n399), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n452), .A2(new_n458), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n454), .A2(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(G22gat), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n461), .A2(new_n462), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n438), .A2(new_n439), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n441), .B1(new_n435), .B2(new_n442), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n451), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n446), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n444), .A2(KEYINPUT80), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n400), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n452), .B1(new_n472), .B2(new_n399), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n464), .B(new_n466), .C1(new_n473), .C2(new_n457), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n432), .B1(new_n465), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT83), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT82), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n466), .B1(new_n473), .B2(new_n457), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n478), .B1(new_n479), .B2(G22gat), .ZN(new_n480));
  INV_X1    g279(.A(new_n432), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n474), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n479), .A2(new_n478), .A3(G22gat), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n477), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT82), .B1(new_n463), .B2(new_n464), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n432), .B1(new_n463), .B2(new_n464), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n486), .A2(new_n487), .A3(new_n477), .A4(new_n484), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n476), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT35), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n429), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT77), .ZN(new_n493));
  NAND2_X1  g292(.A1(G226gat), .A2(G233gat), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT76), .ZN(new_n496));
  XNOR2_X1  g295(.A(KEYINPUT27), .B(G183gat), .ZN(new_n497));
  INV_X1    g296(.A(G190gat), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n497), .B(new_n498), .C1(KEYINPUT68), .C2(KEYINPUT28), .ZN(new_n499));
  NAND2_X1  g298(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(KEYINPUT69), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n499), .B(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(G169gat), .A2(G176gat), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n503), .A2(KEYINPUT26), .ZN(new_n504));
  NAND2_X1  g303(.A1(G169gat), .A2(G176gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n503), .A2(KEYINPUT26), .ZN(new_n507));
  NAND2_X1  g306(.A1(G183gat), .A2(G190gat), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n502), .A2(new_n506), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT25), .ZN(new_n510));
  NAND3_X1  g309(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n511), .B1(G183gat), .B2(G190gat), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT24), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n512), .B1(new_n513), .B2(new_n508), .ZN(new_n514));
  OR2_X1    g313(.A1(new_n503), .A2(KEYINPUT23), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n503), .A2(KEYINPUT23), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n505), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n510), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n515), .A2(KEYINPUT25), .A3(new_n505), .A4(new_n516), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n508), .A2(KEYINPUT64), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT64), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n521), .A2(G183gat), .A3(G190gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT65), .B(KEYINPUT24), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n512), .B1(new_n525), .B2(KEYINPUT66), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT66), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n523), .A2(new_n527), .A3(new_n524), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n519), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT67), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n518), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n523), .A2(new_n527), .A3(new_n524), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n527), .B1(new_n523), .B2(new_n524), .ZN(new_n533));
  NOR3_X1   g332(.A1(new_n532), .A2(new_n533), .A3(new_n512), .ZN(new_n534));
  NOR3_X1   g333(.A1(new_n534), .A2(KEYINPUT67), .A3(new_n519), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n496), .B(new_n509), .C1(new_n531), .C2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT67), .B1(new_n534), .B2(new_n519), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n526), .A2(new_n528), .ZN(new_n539));
  INV_X1    g338(.A(new_n519), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n539), .A2(new_n530), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n538), .A2(new_n541), .A3(new_n518), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n496), .B1(new_n542), .B2(new_n509), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n493), .B(new_n495), .C1(new_n537), .C2(new_n543), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n509), .B1(new_n531), .B2(new_n535), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT76), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n494), .B1(new_n546), .B2(new_n536), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n451), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT77), .B1(new_n548), .B2(new_n494), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n544), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n449), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n451), .B(new_n494), .C1(new_n537), .C2(new_n543), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n542), .A2(new_n495), .A3(new_n509), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n449), .ZN(new_n556));
  XNOR2_X1  g355(.A(G8gat), .B(G36gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(G64gat), .B(G92gat), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n557), .B(new_n558), .Z(new_n559));
  NAND4_X1  g358(.A1(new_n552), .A2(KEYINPUT30), .A3(new_n556), .A4(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n559), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n495), .B1(new_n537), .B2(new_n543), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT29), .B1(new_n542), .B2(new_n509), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n493), .B1(new_n563), .B2(new_n495), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n449), .B1(new_n565), .B2(new_n544), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n551), .B1(new_n553), .B2(new_n554), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n561), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n560), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n567), .B1(new_n550), .B2(new_n551), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT30), .B1(new_n570), .B2(new_n559), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n545), .A2(new_n371), .ZN(new_n573));
  INV_X1    g372(.A(G227gat), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n574), .A2(new_n456), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n402), .B(new_n509), .C1(new_n531), .C2(new_n535), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT32), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT33), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(KEYINPUT73), .B(G71gat), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(G99gat), .ZN(new_n582));
  XOR2_X1   g381(.A(G15gat), .B(G43gat), .Z(new_n583));
  XOR2_X1   g382(.A(new_n582), .B(new_n583), .Z(new_n584));
  NAND3_X1  g383(.A1(new_n578), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n584), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n577), .B(KEYINPUT32), .C1(new_n579), .C2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT75), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n575), .ZN(new_n591));
  INV_X1    g390(.A(new_n576), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n402), .B1(new_n542), .B2(new_n509), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT34), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT34), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n596), .B(new_n591), .C1(new_n592), .C2(new_n593), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n585), .A2(KEYINPUT75), .A3(new_n587), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n590), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n588), .A2(new_n589), .A3(new_n595), .A4(new_n597), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AND3_X1   g401(.A1(new_n492), .A2(new_n572), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT88), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n552), .A2(new_n556), .A3(new_n559), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT30), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT79), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n415), .A2(new_n416), .ZN(new_n610));
  AOI22_X1  g409(.A1(new_n610), .A2(new_n417), .B1(new_n404), .B2(new_n408), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n609), .B1(new_n611), .B2(new_n413), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT6), .B1(new_n611), .B2(new_n413), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n422), .A2(KEYINPUT79), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(new_n424), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n608), .A2(new_n616), .A3(new_n568), .A4(new_n560), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n598), .A2(KEYINPUT74), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n588), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n585), .A2(new_n598), .A3(KEYINPUT74), .A4(new_n587), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(new_n490), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n605), .B(KEYINPUT35), .C1(new_n617), .C2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n486), .A2(new_n487), .A3(new_n484), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT83), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(new_n488), .ZN(new_n627));
  AOI22_X1  g426(.A1(new_n619), .A2(new_n620), .B1(new_n627), .B2(new_n476), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n560), .A2(new_n568), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n628), .A2(new_n629), .A3(new_n616), .A4(new_n608), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n605), .B1(new_n630), .B2(KEYINPUT35), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n604), .B1(new_n624), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(KEYINPUT84), .B1(new_n610), .B2(new_n397), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n415), .A2(new_n416), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT84), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n634), .A2(new_n635), .A3(new_n398), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT39), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n426), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n406), .A2(new_n393), .A3(new_n397), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n633), .A2(KEYINPUT39), .A3(new_n636), .A4(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n639), .A2(KEYINPUT40), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT85), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n639), .A2(KEYINPUT85), .A3(KEYINPUT40), .A4(new_n641), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT40), .B1(new_n639), .B2(new_n641), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n647), .A2(new_n422), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n646), .B(new_n648), .C1(new_n571), .C2(new_n569), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n429), .B1(new_n570), .B2(new_n559), .ZN(new_n650));
  XOR2_X1   g449(.A(KEYINPUT87), .B(KEYINPUT37), .Z(new_n651));
  AOI21_X1  g450(.A(new_n559), .B1(new_n570), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT38), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n550), .A2(new_n449), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n555), .A2(new_n551), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n654), .A2(KEYINPUT37), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n652), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n650), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(KEYINPUT37), .B1(new_n566), .B2(new_n567), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n653), .B1(new_n652), .B2(new_n659), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n649), .B(new_n490), .C1(new_n658), .C2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT36), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n621), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n663), .B1(new_n662), .B2(new_n602), .ZN(new_n664));
  INV_X1    g463(.A(new_n490), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n617), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n661), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n344), .B1(new_n632), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n616), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(G1gat), .ZN(G1324gat));
  INV_X1    g470(.A(new_n572), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT103), .B(KEYINPUT16), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(G8gat), .ZN(new_n674));
  AND3_X1   g473(.A1(new_n668), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n275), .B1(new_n668), .B2(new_n672), .ZN(new_n676));
  OAI21_X1  g475(.A(KEYINPUT42), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n677), .B1(KEYINPUT42), .B2(new_n675), .ZN(G1325gat));
  INV_X1    g477(.A(G15gat), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n668), .A2(new_n679), .A3(new_n602), .ZN(new_n680));
  INV_X1    g479(.A(new_n664), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n668), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n680), .B1(new_n682), .B2(new_n679), .ZN(G1326gat));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n665), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT43), .B(G22gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  AOI21_X1  g485(.A(new_n244), .B1(new_n632), .B2(new_n667), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n285), .A2(new_n286), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n343), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n689), .A2(new_n690), .A3(new_n316), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n693), .A2(new_n207), .A3(new_n669), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT104), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  INV_X1    g497(.A(new_n667), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n632), .A2(KEYINPUT105), .ZN(new_n700));
  OAI21_X1  g499(.A(KEYINPUT35), .B1(new_n617), .B2(new_n622), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(KEYINPUT88), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n623), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(new_n704), .A3(new_n604), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n699), .B1(new_n700), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n244), .A2(KEYINPUT44), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709));
  OAI22_X1  g508(.A1(new_n706), .A2(new_n708), .B1(new_n709), .B2(new_n687), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n710), .A2(new_n691), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n711), .A2(new_n669), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n697), .B(new_n698), .C1(new_n207), .C2(new_n712), .ZN(G1328gat));
  NOR3_X1   g512(.A1(new_n692), .A2(G36gat), .A3(new_n572), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT46), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n711), .A2(new_n672), .ZN(new_n716));
  INV_X1    g515(.A(G36gat), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(G1329gat));
  AOI21_X1  g517(.A(G43gat), .B1(new_n693), .B2(new_n602), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n681), .A2(G43gat), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n719), .B1(new_n711), .B2(new_n720), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT47), .Z(G1330gat));
  NAND3_X1  g521(.A1(new_n710), .A2(new_n665), .A3(new_n691), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(G50gat), .ZN(new_n724));
  INV_X1    g523(.A(G50gat), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n665), .A2(new_n725), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n692), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT48), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT106), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n692), .B2(new_n726), .ZN(new_n731));
  OR3_X1    g530(.A1(new_n692), .A2(new_n730), .A3(new_n726), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n724), .A2(KEYINPUT48), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n729), .A2(KEYINPUT107), .A3(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n732), .A2(KEYINPUT48), .A3(new_n731), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n736), .B1(G50gat), .B2(new_n723), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n735), .B1(new_n728), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n734), .A2(new_n738), .ZN(G1331gat));
  AOI21_X1  g538(.A(new_n704), .B1(new_n703), .B2(new_n604), .ZN(new_n740));
  AOI211_X1 g539(.A(KEYINPUT105), .B(new_n603), .C1(new_n702), .C2(new_n623), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n667), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n316), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n287), .A2(new_n343), .A3(new_n743), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n669), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(G57gat), .ZN(G1332gat));
  AND2_X1   g546(.A1(new_n745), .A2(new_n672), .ZN(new_n748));
  NOR2_X1   g547(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n749));
  AND2_X1   g548(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(new_n748), .B2(new_n749), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT108), .ZN(G1333gat));
  NAND3_X1  g552(.A1(new_n745), .A2(G71gat), .A3(new_n681), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT109), .ZN(new_n755));
  INV_X1    g554(.A(G71gat), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n742), .A2(new_n744), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n602), .B(KEYINPUT110), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT50), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT50), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n755), .A2(new_n762), .A3(new_n759), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(G1334gat));
  NAND2_X1  g563(.A1(new_n745), .A2(new_n665), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g565(.A1(new_n689), .A2(new_n343), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n768), .A2(new_n743), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n710), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(G85gat), .B1(new_n770), .B2(new_n616), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n700), .A2(new_n705), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n244), .B1(new_n772), .B2(new_n667), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT51), .B1(new_n773), .B2(new_n767), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n768), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n742), .A2(new_n243), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT111), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n742), .A2(KEYINPUT111), .A3(new_n243), .A4(new_n776), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n774), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n669), .A2(new_n316), .A3(new_n223), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n771), .B1(new_n781), .B2(new_n782), .ZN(G1336gat));
  NAND3_X1  g582(.A1(new_n710), .A2(new_n672), .A3(new_n769), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G92gat), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT112), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n784), .A2(KEYINPUT112), .A3(G92gat), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n672), .A2(new_n224), .A3(new_n316), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT113), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n774), .A2(new_n791), .B1(new_n779), .B2(new_n780), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n742), .A2(new_n243), .A3(new_n767), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n775), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT113), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n790), .B1(new_n792), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT52), .B1(new_n789), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n785), .B(new_n798), .C1(new_n781), .C2(new_n790), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(G1337gat));
  OAI21_X1  g599(.A(G99gat), .B1(new_n770), .B2(new_n664), .ZN(new_n801));
  INV_X1    g600(.A(new_n602), .ZN(new_n802));
  OR3_X1    g601(.A1(new_n802), .A2(G99gat), .A3(new_n743), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n801), .B1(new_n781), .B2(new_n803), .ZN(G1338gat));
  NAND3_X1  g603(.A1(new_n710), .A2(new_n665), .A3(new_n769), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT53), .B1(new_n805), .B2(G106gat), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n743), .A2(G106gat), .A3(new_n490), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n806), .B(KEYINPUT114), .C1(new_n781), .C2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT111), .B1(new_n773), .B2(new_n776), .ZN(new_n811));
  INV_X1    g610(.A(new_n780), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n794), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n807), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT114), .B1(new_n814), .B2(new_n806), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n774), .A2(new_n791), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n779), .A2(new_n780), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n816), .A2(new_n817), .A3(new_n795), .ZN(new_n818));
  AOI22_X1  g617(.A1(new_n818), .A2(new_n807), .B1(G106gat), .B2(new_n805), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n820));
  OAI22_X1  g619(.A1(new_n810), .A2(new_n815), .B1(new_n819), .B2(new_n820), .ZN(G1339gat));
  NAND3_X1  g620(.A1(new_n299), .A2(new_n289), .A3(new_n300), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n299), .A2(KEYINPUT115), .A3(new_n289), .A4(new_n300), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n824), .A2(new_n302), .A3(KEYINPUT54), .A4(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n308), .B1(new_n301), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(KEYINPUT55), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n311), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(KEYINPUT116), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n829), .A2(new_n832), .A3(new_n311), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n826), .A2(new_n828), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n343), .A2(new_n831), .A3(new_n833), .A4(new_n836), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n336), .A2(new_n331), .A3(new_n323), .A4(new_n339), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n328), .A2(new_n330), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n839), .B1(new_n338), .B2(new_n337), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n322), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n316), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n837), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n244), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n831), .A2(new_n833), .A3(new_n836), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n842), .A2(KEYINPUT117), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n838), .A2(new_n841), .A3(KEYINPUT117), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n243), .A2(new_n848), .ZN(new_n849));
  OR3_X1    g648(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n845), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n243), .B1(new_n837), .B2(new_n843), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT118), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n852), .A2(new_n855), .A3(new_n688), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n317), .A2(new_n690), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n665), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AND4_X1   g657(.A1(new_n669), .A2(new_n858), .A3(new_n572), .A4(new_n602), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n353), .B1(new_n859), .B2(new_n343), .ZN(new_n860));
  XOR2_X1   g659(.A(new_n860), .B(KEYINPUT119), .Z(new_n861));
  AOI21_X1  g660(.A(new_n616), .B1(new_n856), .B2(new_n857), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n672), .A2(new_n622), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(new_n353), .A3(new_n343), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n861), .A2(new_n866), .ZN(G1340gat));
  AOI21_X1  g666(.A(G120gat), .B1(new_n865), .B2(new_n316), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n743), .A2(new_n351), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n868), .B1(new_n859), .B2(new_n869), .ZN(G1341gat));
  NOR3_X1   g669(.A1(new_n864), .A2(G127gat), .A3(new_n688), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n859), .A2(new_n689), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n871), .B1(G127gat), .B2(new_n872), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT120), .ZN(G1342gat));
  NAND3_X1  g673(.A1(new_n865), .A2(new_n348), .A3(new_n243), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n875), .A2(KEYINPUT56), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n358), .B1(new_n859), .B2(new_n243), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n878), .B1(KEYINPUT56), .B2(new_n875), .ZN(G1343gat));
  INV_X1    g678(.A(KEYINPUT58), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n681), .A2(new_n616), .A3(new_n672), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n856), .A2(new_n857), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT57), .B1(new_n882), .B2(new_n665), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n343), .A2(new_n836), .ZN(new_n884));
  INV_X1    g683(.A(new_n830), .ZN(new_n885));
  AOI22_X1  g684(.A1(new_n884), .A2(new_n885), .B1(new_n316), .B2(new_n842), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n850), .B1(new_n886), .B2(new_n243), .ZN(new_n887));
  AOI22_X1  g686(.A1(new_n887), .A2(new_n688), .B1(new_n317), .B2(new_n690), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n490), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n881), .B1(new_n883), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(G141gat), .B1(new_n893), .B2(new_n690), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT121), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n880), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n681), .A2(new_n490), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n898), .A2(new_n672), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n862), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(new_n381), .A3(new_n343), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n894), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n896), .B(new_n903), .ZN(G1344gat));
  NAND3_X1  g703(.A1(new_n901), .A2(new_n383), .A3(new_n316), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n889), .B1(new_n888), .B2(new_n490), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n891), .B1(new_n856), .B2(new_n857), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(KEYINPUT122), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n908), .A2(KEYINPUT122), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n316), .A3(new_n881), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n906), .B1(new_n912), .B2(G148gat), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n893), .A2(new_n743), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n914), .A2(KEYINPUT59), .A3(new_n383), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n905), .B1(new_n913), .B2(new_n915), .ZN(G1345gat));
  OAI21_X1  g715(.A(G155gat), .B1(new_n893), .B2(new_n688), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n901), .A2(new_n387), .A3(new_n689), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1346gat));
  NOR3_X1   g718(.A1(new_n893), .A2(new_n388), .A3(new_n244), .ZN(new_n920));
  AOI21_X1  g719(.A(G162gat), .B1(new_n901), .B2(new_n243), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n920), .A2(new_n921), .ZN(G1347gat));
  NAND2_X1  g721(.A1(new_n672), .A2(new_n616), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n758), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n858), .A2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(G169gat), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n925), .A2(new_n926), .A3(new_n690), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n669), .B1(new_n856), .B2(new_n857), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT123), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n672), .B1(new_n928), .B2(new_n929), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n628), .A3(new_n343), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n927), .B1(new_n934), .B2(new_n926), .ZN(G1348gat));
  INV_X1    g734(.A(G176gat), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n925), .A2(new_n936), .A3(new_n743), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n933), .A2(new_n628), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n936), .B1(new_n938), .B2(new_n743), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT124), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI211_X1 g740(.A(KEYINPUT124), .B(new_n936), .C1(new_n938), .C2(new_n743), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n937), .B1(new_n941), .B2(new_n942), .ZN(G1349gat));
  OAI21_X1  g742(.A(G183gat), .B1(new_n925), .B2(new_n688), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n689), .A2(new_n497), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n938), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g746(.A(G190gat), .B1(new_n925), .B2(new_n244), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT61), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n243), .A2(new_n498), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n938), .B2(new_n950), .ZN(G1351gat));
  XOR2_X1   g750(.A(KEYINPUT125), .B(G197gat), .Z(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n681), .A2(new_n923), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n911), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n953), .B1(new_n955), .B2(new_n690), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n882), .A2(new_n616), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n572), .B1(new_n957), .B2(KEYINPUT123), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n958), .A2(new_n897), .A3(new_n930), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n343), .A2(new_n952), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(G1352gat));
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n681), .A2(new_n743), .A3(new_n923), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n963), .B1(new_n909), .B2(new_n910), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI211_X1 g765(.A(KEYINPUT126), .B(new_n963), .C1(new_n909), .C2(new_n910), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n966), .A2(G204gat), .A3(new_n967), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n743), .A2(G204gat), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(KEYINPUT62), .B1(new_n959), .B2(new_n970), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT62), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n933), .A2(new_n972), .A3(new_n897), .A4(new_n969), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n962), .B1(new_n968), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n966), .A2(G204gat), .A3(new_n967), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n976), .A2(KEYINPUT127), .A3(new_n971), .A4(new_n973), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n975), .A2(new_n977), .ZN(G1353gat));
  OR3_X1    g777(.A1(new_n959), .A2(G211gat), .A3(new_n688), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n911), .A2(new_n689), .A3(new_n954), .ZN(new_n980));
  AND3_X1   g779(.A1(new_n980), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n981));
  AOI21_X1  g780(.A(KEYINPUT63), .B1(new_n980), .B2(G211gat), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(G1354gat));
  OAI21_X1  g782(.A(G218gat), .B1(new_n955), .B2(new_n244), .ZN(new_n984));
  OR2_X1    g783(.A1(new_n244), .A2(G218gat), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n984), .B1(new_n959), .B2(new_n985), .ZN(G1355gat));
endmodule


