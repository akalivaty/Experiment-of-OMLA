//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0 0 1 1 1 0 0 0 1 0 0 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007;
  INV_X1    g000(.A(KEYINPUT5), .ZN(new_n202));
  NAND2_X1  g001(.A1(G225gat), .A2(G233gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT80), .B(G148gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G141gat), .ZN(new_n205));
  INV_X1    g004(.A(G141gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G148gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT81), .B(G162gat), .ZN(new_n209));
  INV_X1    g008(.A(G155gat), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT2), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G155gat), .B(G162gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n208), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT2), .ZN(new_n215));
  INV_X1    g014(.A(G148gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G141gat), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n215), .A2(KEYINPUT79), .B1(new_n207), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n215), .A2(KEYINPUT79), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT78), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n221), .B1(G155gat), .B2(G162gat), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n222), .B1(new_n212), .B2(new_n221), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n213), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G127gat), .B(G134gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT67), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OR2_X1    g027(.A1(G127gat), .A2(G134gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(G127gat), .A2(G134gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n229), .A2(KEYINPUT67), .A3(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G113gat), .B(G120gat), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n228), .B(new_n231), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n226), .A2(KEYINPUT69), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT69), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n229), .A2(new_n235), .A3(new_n230), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n232), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G113gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n240), .A2(G120gat), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT1), .B1(new_n241), .B2(KEYINPUT68), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n233), .B1(new_n237), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n225), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n234), .A2(new_n236), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n246), .A2(new_n239), .A3(new_n242), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n213), .A2(new_n247), .A3(new_n224), .A4(new_n233), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n203), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n202), .B1(new_n249), .B2(KEYINPUT82), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n225), .A2(KEYINPUT3), .ZN(new_n251));
  INV_X1    g050(.A(new_n212), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n252), .B1(new_n205), .B2(new_n207), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n253), .A2(new_n211), .B1(new_n220), .B2(new_n223), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT3), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n251), .A2(new_n256), .A3(new_n244), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n248), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n244), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n260), .A2(KEYINPUT4), .A3(new_n254), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n257), .A2(new_n203), .A3(new_n259), .A4(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n203), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n225), .A2(new_n244), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n213), .A2(new_n224), .B1(new_n247), .B2(new_n233), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT82), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n262), .A3(new_n268), .ZN(new_n269));
  AND2_X1   g068(.A1(new_n261), .A2(new_n259), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n270), .A2(new_n202), .A3(new_n203), .A4(new_n257), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G1gat), .B(G29gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(KEYINPUT0), .ZN(new_n274));
  XNOR2_X1  g073(.A(G57gat), .B(G85gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n272), .A2(KEYINPUT6), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT83), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  XOR2_X1   g078(.A(new_n276), .B(KEYINPUT87), .Z(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n272), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n283));
  INV_X1    g082(.A(new_n276), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n269), .A2(new_n284), .A3(new_n271), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n282), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n284), .B1(new_n269), .B2(new_n271), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n287), .A2(KEYINPUT83), .A3(KEYINPUT6), .ZN(new_n288));
  AND3_X1   g087(.A1(new_n279), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n290));
  NOR2_X1   g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n291), .B1(KEYINPUT23), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT65), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G183gat), .A2(G190gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT24), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT24), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(G183gat), .A3(G190gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n293), .B1(new_n298), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n291), .A2(KEYINPUT23), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT66), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n291), .A2(KEYINPUT66), .A3(KEYINPUT23), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT25), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n294), .B1(new_n300), .B2(new_n302), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n305), .A2(KEYINPUT25), .ZN(new_n314));
  NOR3_X1   g113(.A1(new_n313), .A2(new_n314), .A3(new_n293), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(KEYINPUT27), .B(G183gat), .ZN(new_n317));
  INV_X1    g116(.A(G190gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT28), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n317), .A2(KEYINPUT28), .A3(new_n318), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n291), .A2(KEYINPUT26), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n299), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n291), .A2(KEYINPUT26), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n325), .B1(new_n292), .B2(new_n326), .ZN(new_n327));
  AOI22_X1  g126(.A1(new_n312), .A2(new_n316), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(G226gat), .A2(G233gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n329), .B(KEYINPUT71), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(KEYINPUT72), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n290), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n330), .B1(new_n328), .B2(KEYINPUT29), .ZN(new_n333));
  XNOR2_X1  g132(.A(G197gat), .B(G204gat), .ZN(new_n334));
  INV_X1    g133(.A(G211gat), .ZN(new_n335));
  INV_X1    g134(.A(G218gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n334), .B1(KEYINPUT22), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G211gat), .B(G218gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n323), .A2(new_n327), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT25), .B1(new_n304), .B2(new_n309), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n342), .B1(new_n343), .B2(new_n315), .ZN(new_n344));
  INV_X1    g143(.A(new_n331), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n344), .A2(KEYINPUT73), .A3(new_n345), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n332), .A2(new_n333), .A3(new_n341), .A4(new_n346), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n328), .A2(new_n330), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT29), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n345), .B1(new_n344), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n340), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n347), .A2(KEYINPUT74), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n312), .A2(new_n316), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n331), .B1(new_n353), .B2(new_n342), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n344), .A2(new_n349), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n354), .A2(KEYINPUT73), .B1(new_n355), .B2(new_n330), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT74), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n356), .A2(new_n357), .A3(new_n341), .A4(new_n332), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n352), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT37), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  XOR2_X1   g160(.A(G8gat), .B(G36gat), .Z(new_n362));
  XNOR2_X1  g161(.A(new_n362), .B(KEYINPUT75), .ZN(new_n363));
  XNOR2_X1  g162(.A(G64gat), .B(G92gat), .ZN(new_n364));
  XOR2_X1   g163(.A(new_n363), .B(new_n364), .Z(new_n365));
  NAND3_X1  g164(.A1(new_n352), .A2(KEYINPUT37), .A3(new_n358), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n361), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT38), .ZN(new_n368));
  INV_X1    g167(.A(new_n365), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT76), .B1(new_n359), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT76), .ZN(new_n371));
  AOI211_X1 g170(.A(new_n371), .B(new_n365), .C1(new_n352), .C2(new_n358), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  OR2_X1    g172(.A1(new_n348), .A2(new_n350), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n360), .B1(new_n374), .B2(new_n341), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n356), .A2(new_n340), .A3(new_n332), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT38), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n377), .A3(new_n365), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n289), .A2(new_n368), .A3(new_n373), .A4(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n225), .A2(KEYINPUT3), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n244), .B1(new_n254), .B2(new_n255), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n261), .B(new_n259), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n263), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT39), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n264), .A2(new_n265), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n384), .B1(new_n385), .B2(new_n203), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n387), .B(new_n280), .C1(KEYINPUT39), .C2(new_n383), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT40), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n282), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n388), .A2(new_n389), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT77), .B(KEYINPUT30), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NOR3_X1   g194(.A1(new_n370), .A2(new_n372), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n365), .B1(new_n352), .B2(new_n358), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT30), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n398), .B1(new_n369), .B2(new_n359), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n393), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n401));
  INV_X1    g200(.A(G22gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n255), .B1(new_n340), .B2(KEYINPUT29), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n225), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n256), .A2(KEYINPUT86), .A3(new_n349), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n340), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT86), .B1(new_n256), .B2(new_n349), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n406), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(G228gat), .ZN(new_n411));
  INV_X1    g210(.A(G233gat), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n340), .B1(new_n380), .B2(KEYINPUT29), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n415), .B(new_n406), .C1(new_n411), .C2(new_n412), .ZN(new_n416));
  XNOR2_X1  g215(.A(G78gat), .B(G106gat), .ZN(new_n417));
  INV_X1    g216(.A(G50gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT85), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n414), .A2(new_n416), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n421), .B1(new_n414), .B2(new_n416), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n404), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n424), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n426), .A2(new_n403), .A3(new_n422), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n379), .A2(new_n400), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n344), .A2(new_n260), .ZN(new_n431));
  NAND2_X1  g230(.A1(G227gat), .A2(G233gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(KEYINPUT64), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n244), .B(new_n342), .C1(new_n343), .C2(new_n315), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n431), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  XOR2_X1   g234(.A(KEYINPUT70), .B(KEYINPUT33), .Z(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  XOR2_X1   g236(.A(G15gat), .B(G43gat), .Z(new_n438));
  XNOR2_X1  g237(.A(G71gat), .B(G99gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n431), .A2(new_n434), .ZN(new_n442));
  INV_X1    g241(.A(new_n433), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT34), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT34), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n442), .A2(new_n446), .A3(new_n443), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n441), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n435), .A2(KEYINPUT32), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n440), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n451), .B1(new_n435), .B2(new_n436), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n446), .B1(new_n442), .B2(new_n443), .ZN(new_n453));
  AOI211_X1 g252(.A(KEYINPUT34), .B(new_n433), .C1(new_n431), .C2(new_n434), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n448), .A2(new_n450), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n450), .B1(new_n448), .B2(new_n455), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT36), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n455), .ZN(new_n460));
  NOR3_X1   g259(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n449), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n448), .A2(new_n450), .A3(new_n455), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT36), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n359), .A2(new_n369), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n371), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n397), .A2(KEYINPUT76), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(new_n468), .A3(new_n394), .ZN(new_n469));
  INV_X1    g268(.A(new_n287), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n470), .A2(new_n283), .A3(new_n285), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n471), .A2(new_n279), .A3(new_n288), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n359), .A2(new_n369), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n473), .B1(KEYINPUT30), .B2(new_n397), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n469), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n465), .B1(new_n475), .B2(new_n428), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n430), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n456), .A2(new_n457), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n478), .A2(new_n427), .A3(new_n425), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT35), .B1(new_n475), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n396), .A2(new_n399), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n478), .A2(new_n427), .A3(new_n425), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n287), .A2(KEYINPUT83), .A3(KEYINPUT6), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT83), .B1(new_n287), .B2(KEYINPUT6), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT35), .B1(new_n485), .B2(new_n286), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n481), .A2(new_n482), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n480), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n477), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT98), .ZN(new_n490));
  XOR2_X1   g289(.A(G183gat), .B(G211gat), .Z(new_n491));
  INV_X1    g290(.A(KEYINPUT91), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(G57gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(G64gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(G71gat), .A2(G78gat), .ZN(new_n495));
  OR2_X1    g294(.A1(G71gat), .A2(G78gat), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT9), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n496), .A2(new_n495), .ZN(new_n500));
  OR2_X1    g299(.A1(G57gat), .A2(G64gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(G57gat), .A2(G64gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(KEYINPUT9), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  XOR2_X1   g304(.A(KEYINPUT92), .B(KEYINPUT21), .Z(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(G231gat), .A2(G233gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(G127gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n509), .A2(new_n510), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n491), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n513), .ZN(new_n515));
  INV_X1    g314(.A(new_n491), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n511), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT89), .ZN(new_n519));
  XNOR2_X1  g318(.A(G15gat), .B(G22gat), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n519), .B1(new_n520), .B2(G1gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n402), .A2(G15gat), .ZN(new_n522));
  INV_X1    g321(.A(G15gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(G22gat), .ZN(new_n524));
  INV_X1    g323(.A(G1gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT16), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n522), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(G8gat), .B1(new_n521), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n522), .A2(new_n524), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT89), .B1(new_n529), .B2(new_n525), .ZN(new_n530));
  INV_X1    g329(.A(G8gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n520), .A2(new_n526), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT21), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n535), .B1(new_n536), .B2(new_n505), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT93), .ZN(new_n538));
  XNOR2_X1  g337(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(new_n210), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n538), .A2(new_n540), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n518), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n514), .A2(new_n541), .A3(new_n517), .A4(new_n542), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT17), .ZN(new_n548));
  INV_X1    g347(.A(G29gat), .ZN(new_n549));
  INV_X1    g348(.A(G36gat), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n549), .A2(new_n550), .A3(KEYINPUT14), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT14), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(G29gat), .B2(G36gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(G29gat), .A2(G36gat), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n551), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(G43gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(G50gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n418), .A2(G43gat), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n555), .A2(KEYINPUT15), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT88), .B1(new_n418), .B2(G43gat), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n418), .A2(G43gat), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n418), .A2(KEYINPUT88), .A3(G43gat), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT15), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n557), .A2(new_n558), .A3(KEYINPUT15), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n565), .A2(new_n553), .A3(new_n551), .A4(new_n554), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n548), .B(new_n559), .C1(new_n564), .C2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT88), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n569), .B1(new_n556), .B2(G50gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n570), .A2(new_n557), .A3(new_n563), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT15), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n555), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n573), .A2(new_n565), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n548), .B1(new_n575), .B2(new_n559), .ZN(new_n576));
  INV_X1    g375(.A(G92gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT95), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT95), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(G92gat), .ZN(new_n580));
  INV_X1    g379(.A(G85gat), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n578), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n583));
  NAND2_X1  g382(.A1(G85gat), .A2(G92gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(G99gat), .A2(G106gat), .ZN(new_n585));
  AOI22_X1  g384(.A1(new_n583), .A2(new_n584), .B1(new_n585), .B2(KEYINPUT8), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT94), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT7), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n590));
  AND2_X1   g389(.A1(G85gat), .A2(G92gat), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n582), .A2(new_n586), .A3(new_n592), .ZN(new_n593));
  AND2_X1   g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(G99gat), .A2(G106gat), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT96), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(G99gat), .ZN(new_n597));
  INV_X1    g396(.A(G106gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT96), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(new_n600), .A3(new_n585), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n593), .A2(new_n602), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n593), .A2(new_n602), .ZN(new_n604));
  OAI22_X1  g403(.A1(new_n568), .A2(new_n576), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n603), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n559), .B1(new_n564), .B2(new_n566), .ZN(new_n607));
  NAND2_X1  g406(.A1(G232gat), .A2(G233gat), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  AOI22_X1  g408(.A1(new_n606), .A2(new_n607), .B1(KEYINPUT41), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G190gat), .B(G218gat), .Z(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n609), .A2(KEYINPUT41), .ZN(new_n614));
  XNOR2_X1  g413(.A(G134gat), .B(G162gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n612), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n605), .A2(new_n610), .A3(new_n617), .ZN(new_n618));
  AND3_X1   g417(.A1(new_n613), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n616), .B1(new_n613), .B2(new_n618), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n505), .B1(new_n604), .B2(new_n603), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n582), .A2(new_n586), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n596), .A2(new_n601), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n624), .A2(new_n625), .A3(new_n592), .ZN(new_n626));
  AOI22_X1  g425(.A1(new_n494), .A2(new_n498), .B1(new_n503), .B2(new_n500), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n593), .A2(new_n602), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G230gat), .A2(G233gat), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G120gat), .B(G148gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(G176gat), .B(G204gat), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n634), .B(new_n635), .Z(new_n636));
  NAND2_X1  g435(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT10), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n623), .A2(new_n638), .A3(new_n629), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n606), .A2(KEYINPUT10), .A3(new_n627), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT97), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n632), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n639), .A2(KEYINPUT97), .A3(new_n640), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n637), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n641), .A2(new_n631), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n636), .B1(new_n646), .B2(new_n633), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n547), .A2(new_n622), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT90), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n534), .A2(new_n607), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n607), .A2(KEYINPUT17), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n567), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n652), .B1(new_n654), .B2(new_n535), .ZN(new_n655));
  NAND2_X1  g454(.A1(G229gat), .A2(G233gat), .ZN(new_n656));
  AOI21_X1  g455(.A(KEYINPUT18), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(G197gat), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n206), .A2(G113gat), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n240), .A2(G141gat), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n659), .A2(new_n660), .A3(new_n658), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT11), .B(G169gat), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n664), .ZN(new_n666));
  INV_X1    g465(.A(new_n663), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n666), .B1(new_n667), .B2(new_n661), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n665), .A2(new_n668), .A3(KEYINPUT12), .ZN(new_n669));
  AOI21_X1  g468(.A(KEYINPUT12), .B1(new_n665), .B2(new_n668), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n534), .A2(new_n607), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n528), .A2(new_n575), .A3(new_n533), .A4(new_n559), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n656), .B(KEYINPUT13), .Z(new_n675));
  AOI21_X1  g474(.A(new_n671), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n535), .B1(new_n568), .B2(new_n576), .ZN(new_n677));
  INV_X1    g476(.A(new_n656), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT18), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n677), .A2(new_n672), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n651), .B1(new_n657), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n677), .A2(new_n672), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n679), .B1(new_n684), .B2(new_n678), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n685), .A2(KEYINPUT90), .A3(new_n681), .A4(new_n676), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n674), .A2(new_n675), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n685), .A2(new_n681), .A3(new_n687), .ZN(new_n688));
  AOI22_X1  g487(.A1(new_n683), .A2(new_n686), .B1(new_n688), .B2(new_n671), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n650), .A2(new_n689), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n489), .A2(new_n490), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n490), .B1(new_n489), .B2(new_n690), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(new_n472), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(new_n525), .ZN(G1324gat));
  NOR2_X1   g494(.A1(new_n693), .A2(new_n481), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT16), .B(G8gat), .Z(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n698), .B1(new_n531), .B2(new_n696), .ZN(new_n699));
  MUX2_X1   g498(.A(new_n698), .B(new_n699), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g499(.A(new_n465), .ZN(new_n701));
  OAI21_X1  g500(.A(G15gat), .B1(new_n693), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n478), .A2(new_n523), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n702), .B1(new_n693), .B2(new_n703), .ZN(G1326gat));
  NOR2_X1   g503(.A1(new_n693), .A2(new_n429), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT43), .B(G22gat), .Z(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1327gat));
  NAND2_X1  g506(.A1(new_n489), .A2(new_n621), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n547), .A2(new_n689), .A3(new_n648), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n472), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n711), .A2(new_n549), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT45), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n430), .A2(new_n476), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n488), .A2(KEYINPUT99), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT99), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n480), .A2(new_n487), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n716), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n715), .B1(new_n720), .B2(new_n622), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n622), .B1(new_n477), .B2(new_n488), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(KEYINPUT44), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n724), .A2(new_n472), .A3(new_n710), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n714), .B1(new_n725), .B2(new_n549), .ZN(G1328gat));
  INV_X1    g525(.A(new_n481), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n550), .A3(new_n727), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n728), .B(KEYINPUT46), .Z(new_n729));
  NOR3_X1   g528(.A1(new_n724), .A2(new_n481), .A3(new_n710), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(new_n730), .B2(new_n550), .ZN(G1329gat));
  NAND4_X1  g530(.A1(new_n721), .A2(new_n465), .A3(new_n709), .A4(new_n723), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G43gat), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n456), .A2(new_n457), .A3(G43gat), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n722), .A2(new_n709), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT100), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT100), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n722), .A2(new_n737), .A3(new_n709), .A4(new_n734), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n733), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT47), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT101), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n739), .B1(new_n732), .B2(G43gat), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT101), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n744), .A2(new_n745), .A3(KEYINPUT47), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT102), .ZN(new_n747));
  AND4_X1   g546(.A1(new_n747), .A2(new_n733), .A3(KEYINPUT47), .A4(new_n740), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n747), .B1(new_n744), .B2(KEYINPUT47), .ZN(new_n749));
  OAI22_X1  g548(.A1(new_n743), .A2(new_n746), .B1(new_n748), .B2(new_n749), .ZN(G1330gat));
  NAND2_X1  g549(.A1(new_n428), .A2(new_n418), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT103), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n711), .A2(new_n752), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n724), .A2(new_n429), .A3(new_n710), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n753), .B1(new_n754), .B2(new_n418), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT48), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI211_X1 g556(.A(KEYINPUT48), .B(new_n753), .C1(new_n754), .C2(new_n418), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(G1331gat));
  AND3_X1   g558(.A1(new_n480), .A2(new_n487), .A3(new_n718), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n718), .B1(new_n480), .B2(new_n487), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n477), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n689), .ZN(new_n763));
  NOR4_X1   g562(.A1(new_n546), .A2(new_n763), .A3(new_n649), .A4(new_n621), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n712), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g567(.A1(new_n765), .A2(new_n481), .ZN(new_n769));
  NOR2_X1   g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  AND2_X1   g569(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n772), .B1(new_n769), .B2(new_n770), .ZN(G1333gat));
  AND3_X1   g572(.A1(new_n766), .A2(G71gat), .A3(new_n465), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n478), .B(KEYINPUT104), .ZN(new_n775));
  AOI21_X1  g574(.A(G71gat), .B1(new_n766), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  XOR2_X1   g576(.A(new_n777), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g577(.A1(new_n766), .A2(new_n428), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g579(.A(KEYINPUT44), .B1(new_n762), .B2(new_n621), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n708), .A2(new_n715), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n547), .A2(new_n763), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n648), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n781), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(G85gat), .B1(new_n786), .B2(new_n472), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n762), .A2(new_n621), .A3(new_n783), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n712), .A2(new_n581), .A3(new_n648), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n787), .B1(new_n791), .B2(new_n792), .ZN(G1336gat));
  AOI22_X1  g592(.A1(new_n785), .A2(new_n727), .B1(new_n578), .B2(new_n580), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(KEYINPUT52), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n481), .A2(G92gat), .A3(new_n649), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n790), .A2(KEYINPUT106), .A3(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT106), .B1(new_n790), .B2(new_n796), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n795), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  XOR2_X1   g598(.A(new_n796), .B(KEYINPUT105), .Z(new_n800));
  AND2_X1   g599(.A1(new_n790), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT52), .B1(new_n801), .B2(new_n794), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n799), .A2(new_n802), .ZN(G1337gat));
  OAI21_X1  g602(.A(G99gat), .B1(new_n786), .B2(new_n701), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n478), .A2(new_n597), .A3(new_n648), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n791), .B2(new_n805), .ZN(G1338gat));
  NAND2_X1  g605(.A1(new_n785), .A2(new_n428), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(G106gat), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n429), .A2(G106gat), .A3(new_n649), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n790), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT53), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n808), .A2(new_n813), .A3(new_n810), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(G1339gat));
  NAND2_X1  g614(.A1(new_n641), .A2(new_n642), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n816), .A2(new_n631), .A3(new_n644), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n639), .A2(new_n632), .A3(new_n640), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT54), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g620(.A(KEYINPUT107), .B(KEYINPUT54), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n641), .A2(new_n631), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n636), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n821), .A2(KEYINPUT55), .A3(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT108), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n825), .B1(new_n817), .B2(new_n820), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n830), .A2(KEYINPUT108), .A3(KEYINPUT55), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT55), .B1(new_n821), .B2(new_n826), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n645), .B1(new_n833), .B2(KEYINPUT109), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n819), .B1(new_n643), .B2(new_n644), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n836), .B2(new_n825), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT109), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n832), .A2(new_n834), .A3(new_n763), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n683), .A2(new_n686), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n655), .A2(new_n656), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n674), .A2(new_n675), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n665), .B(new_n668), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n648), .A2(new_n841), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n621), .B1(new_n840), .B2(new_n845), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n621), .A2(new_n841), .A3(new_n844), .ZN(new_n847));
  AND4_X1   g646(.A1(new_n832), .A2(new_n839), .A3(new_n834), .A4(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n546), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n650), .A2(new_n763), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n428), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n851), .A2(new_n712), .A3(new_n481), .A4(new_n478), .ZN(new_n852));
  OAI21_X1  g651(.A(G113gat), .B1(new_n852), .B2(new_n689), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n689), .A2(G113gat), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT110), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n853), .B1(new_n852), .B2(new_n855), .ZN(G1340gat));
  OAI21_X1  g655(.A(G120gat), .B1(new_n852), .B2(new_n649), .ZN(new_n857));
  XOR2_X1   g656(.A(new_n857), .B(KEYINPUT111), .Z(new_n858));
  NOR2_X1   g657(.A1(new_n649), .A2(G120gat), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT112), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n858), .B1(new_n852), .B2(new_n860), .ZN(G1341gat));
  NOR2_X1   g660(.A1(new_n852), .A2(new_n546), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(new_n510), .ZN(G1342gat));
  NOR2_X1   g662(.A1(new_n727), .A2(new_n622), .ZN(new_n864));
  INV_X1    g663(.A(new_n478), .ZN(new_n865));
  AOI211_X1 g664(.A(new_n472), .B(new_n865), .C1(KEYINPUT56), .C2(G134gat), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n851), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n868));
  XOR2_X1   g667(.A(new_n867), .B(new_n868), .Z(G1343gat));
  NAND2_X1  g668(.A1(new_n701), .A2(new_n428), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(KEYINPUT115), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n472), .B1(new_n849), .B2(new_n850), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n871), .B1(new_n872), .B2(KEYINPUT114), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n872), .A2(KEYINPUT114), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n689), .A2(G141gat), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n481), .A3(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT116), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n727), .A2(new_n472), .A3(new_n465), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n849), .A2(new_n850), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT57), .B1(new_n881), .B2(new_n428), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n650), .A2(new_n763), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n832), .A2(new_n834), .A3(new_n839), .A4(new_n847), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n648), .A2(new_n841), .A3(new_n844), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n689), .A2(new_n833), .A3(new_n645), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n885), .B1(new_n886), .B2(new_n832), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n884), .B1(new_n887), .B2(new_n621), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n883), .B1(new_n888), .B2(new_n546), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n428), .A2(KEYINPUT57), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n880), .B1(new_n882), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(G141gat), .B1(new_n892), .B2(new_n689), .ZN(new_n893));
  OAI22_X1  g692(.A1(new_n878), .A2(new_n879), .B1(KEYINPUT113), .B2(new_n893), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n893), .A2(KEYINPUT113), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT58), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(KEYINPUT116), .A2(KEYINPUT58), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n878), .B(new_n897), .C1(new_n893), .C2(KEYINPUT58), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(G1344gat));
  INV_X1    g698(.A(KEYINPUT119), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n892), .A2(new_n649), .ZN(new_n901));
  INV_X1    g700(.A(new_n204), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT117), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n688), .A2(new_n671), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n645), .B1(new_n841), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(KEYINPUT108), .B1(new_n830), .B2(KEYINPUT55), .ZN(new_n909));
  NOR4_X1   g708(.A1(new_n836), .A2(new_n825), .A3(new_n828), .A4(new_n835), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n908), .B(new_n837), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n621), .B1(new_n911), .B2(new_n845), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n546), .B1(new_n912), .B2(new_n848), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n429), .B1(new_n913), .B2(new_n850), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n906), .B1(new_n914), .B2(KEYINPUT57), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT57), .ZN(new_n916));
  OAI211_X1 g715(.A(KEYINPUT117), .B(new_n916), .C1(new_n889), .C2(new_n429), .ZN(new_n917));
  INV_X1    g716(.A(new_n890), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n881), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n915), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n880), .A2(new_n648), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT118), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n920), .A2(KEYINPUT118), .A3(new_n921), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n924), .A2(G148gat), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n905), .B1(new_n926), .B2(KEYINPUT59), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n875), .A2(new_n727), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n649), .A2(new_n902), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n900), .B1(new_n927), .B2(new_n931), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n925), .A2(G148gat), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n903), .B1(new_n933), .B2(new_n924), .ZN(new_n934));
  OAI211_X1 g733(.A(KEYINPUT119), .B(new_n930), .C1(new_n934), .C2(new_n905), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n932), .A2(new_n935), .ZN(G1345gat));
  NAND3_X1  g735(.A1(new_n928), .A2(new_n210), .A3(new_n547), .ZN(new_n937));
  OAI21_X1  g736(.A(G155gat), .B1(new_n892), .B2(new_n546), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1346gat));
  NAND3_X1  g738(.A1(new_n876), .A2(new_n209), .A3(new_n864), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n892), .A2(new_n622), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n209), .B2(new_n941), .ZN(G1347gat));
  NAND2_X1  g741(.A1(new_n881), .A2(new_n472), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n943), .A2(KEYINPUT120), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n943), .A2(KEYINPUT120), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n481), .A2(new_n479), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OR2_X1    g747(.A1(new_n689), .A2(G169gat), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n727), .A2(new_n472), .ZN(new_n950));
  INV_X1    g749(.A(new_n775), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n851), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(G169gat), .B1(new_n953), .B2(new_n689), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n954), .A2(KEYINPUT121), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n954), .A2(KEYINPUT121), .ZN(new_n956));
  OAI22_X1  g755(.A1(new_n948), .A2(new_n949), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT122), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n957), .B(new_n958), .ZN(G1348gat));
  OAI21_X1  g758(.A(G176gat), .B1(new_n953), .B2(new_n649), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n649), .A2(G176gat), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n960), .B1(new_n948), .B2(new_n961), .ZN(G1349gat));
  OAI21_X1  g761(.A(G183gat), .B1(new_n953), .B2(new_n546), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n547), .A2(new_n317), .ZN(new_n964));
  OAI211_X1 g763(.A(new_n947), .B(new_n964), .C1(new_n944), .C2(new_n945), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT123), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n965), .A2(new_n966), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n963), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(KEYINPUT60), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT60), .ZN(new_n971));
  OAI211_X1 g770(.A(new_n971), .B(new_n963), .C1(new_n967), .C2(new_n968), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(new_n972), .ZN(G1350gat));
  OAI21_X1  g772(.A(G190gat), .B1(new_n953), .B2(new_n622), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT61), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n622), .A2(G190gat), .ZN(new_n976));
  OAI211_X1 g775(.A(new_n947), .B(new_n976), .C1(new_n944), .C2(new_n945), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n977), .A2(KEYINPUT124), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n977), .A2(KEYINPUT124), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n975), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(KEYINPUT125), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT125), .ZN(new_n982));
  OAI211_X1 g781(.A(new_n982), .B(new_n975), .C1(new_n978), .C2(new_n979), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n981), .A2(new_n983), .ZN(G1351gat));
  NOR2_X1   g783(.A1(new_n870), .A2(new_n481), .ZN(new_n985));
  AND2_X1   g784(.A1(new_n946), .A2(new_n985), .ZN(new_n986));
  XOR2_X1   g785(.A(KEYINPUT126), .B(G197gat), .Z(new_n987));
  NAND3_X1  g786(.A1(new_n986), .A2(new_n763), .A3(new_n987), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n920), .A2(new_n472), .A3(new_n727), .A4(new_n701), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n989), .A2(new_n689), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n988), .B1(new_n990), .B2(new_n987), .ZN(G1352gat));
  NOR2_X1   g790(.A1(new_n649), .A2(G204gat), .ZN(new_n992));
  OAI211_X1 g791(.A(new_n985), .B(new_n992), .C1(new_n944), .C2(new_n945), .ZN(new_n993));
  OR2_X1    g792(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n994));
  OAI21_X1  g793(.A(G204gat), .B1(new_n989), .B2(new_n649), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT127), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g798(.A1(new_n994), .A2(KEYINPUT127), .A3(new_n995), .A4(new_n996), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(G1353gat));
  OAI21_X1  g800(.A(G211gat), .B1(new_n989), .B2(new_n546), .ZN(new_n1002));
  XOR2_X1   g801(.A(new_n1002), .B(KEYINPUT63), .Z(new_n1003));
  NAND3_X1  g802(.A1(new_n986), .A2(new_n335), .A3(new_n547), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(new_n1004), .ZN(G1354gat));
  NAND3_X1  g804(.A1(new_n986), .A2(new_n336), .A3(new_n621), .ZN(new_n1006));
  OAI21_X1  g805(.A(G218gat), .B1(new_n989), .B2(new_n622), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1006), .A2(new_n1007), .ZN(G1355gat));
endmodule


