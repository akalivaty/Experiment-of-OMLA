//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n787, new_n788, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005;
  INV_X1    g000(.A(KEYINPUT15), .ZN(new_n202));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203));
  XOR2_X1   g002(.A(KEYINPUT87), .B(G36gat), .Z(new_n204));
  AOI22_X1  g003(.A1(new_n202), .A2(new_n203), .B1(new_n204), .B2(G29gat), .ZN(new_n205));
  OR3_X1    g004(.A1(KEYINPUT86), .A2(G29gat), .A3(G36gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT86), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(KEYINPUT14), .A3(new_n207), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n205), .B(new_n208), .C1(KEYINPUT14), .C2(new_n207), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n203), .A2(new_n202), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n210), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT17), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G15gat), .B(G22gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n216), .B(KEYINPUT88), .ZN(new_n217));
  INV_X1    g016(.A(G1gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n218), .A2(KEYINPUT16), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n219), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G8gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n221), .B(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n211), .A2(KEYINPUT17), .A3(new_n212), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n215), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G229gat), .A2(G233gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n221), .B(G8gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(new_n213), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n225), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT18), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n225), .A2(KEYINPUT18), .A3(new_n226), .A4(new_n228), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n227), .B(new_n213), .ZN(new_n233));
  XOR2_X1   g032(.A(new_n226), .B(KEYINPUT13), .Z(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n231), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G113gat), .B(G141gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n237), .B(G197gat), .ZN(new_n238));
  XOR2_X1   g037(.A(KEYINPUT11), .B(G169gat), .Z(new_n239));
  XNOR2_X1  g038(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n240), .B(KEYINPUT12), .Z(new_n241));
  NAND2_X1  g040(.A1(new_n236), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n241), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n231), .A2(new_n243), .A3(new_n232), .A4(new_n235), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT85), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT82), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT22), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n248), .A2(KEYINPUT76), .B1(G211gat), .B2(G218gat), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n249), .B1(KEYINPUT76), .B2(new_n248), .ZN(new_n250));
  INV_X1    g049(.A(G204gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G197gat), .ZN(new_n252));
  INV_X1    g051(.A(G197gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(G204gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT75), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n252), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n255), .B1(new_n252), .B2(new_n254), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n250), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G211gat), .B(G218gat), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n259), .B(new_n250), .C1(new_n256), .C2(new_n257), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G226gat), .A2(G233gat), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT28), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT27), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(G183gat), .ZN(new_n269));
  INV_X1    g068(.A(G183gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT27), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT67), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT67), .B1(new_n270), .B2(KEYINPUT27), .ZN(new_n273));
  INV_X1    g072(.A(G190gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n267), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n269), .A2(new_n271), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n277), .A2(KEYINPUT28), .A3(new_n274), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(G169gat), .ZN(new_n280));
  INV_X1    g079(.A(G176gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT26), .ZN(new_n283));
  NAND2_X1  g082(.A1(G169gat), .A2(G176gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT26), .ZN(new_n286));
  NAND2_X1  g085(.A1(G183gat), .A2(G190gat), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n279), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT66), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n287), .B1(new_n294), .B2(KEYINPUT24), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n294), .A2(KEYINPUT24), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n292), .B(new_n293), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT23), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT23), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n299), .B1(G169gat), .B2(G176gat), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n298), .A2(new_n300), .A3(new_n284), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n297), .A2(new_n301), .A3(KEYINPUT25), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n304), .A2(new_n292), .A3(new_n293), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT25), .B1(new_n301), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n302), .B1(new_n306), .B2(KEYINPUT65), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT25), .ZN(new_n308));
  AND3_X1   g107(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n309));
  NOR3_X1   g108(.A1(new_n309), .A2(new_n303), .A3(new_n291), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n298), .A2(new_n300), .A3(new_n284), .ZN(new_n311));
  OAI211_X1 g110(.A(KEYINPUT65), .B(new_n308), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n290), .B1(new_n307), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n266), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n308), .B1(new_n310), .B2(new_n311), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT65), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n311), .A2(new_n308), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n317), .A2(new_n318), .B1(new_n319), .B2(new_n297), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(new_n312), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n265), .B1(new_n321), .B2(new_n290), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n264), .B1(new_n316), .B2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G8gat), .B(G36gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(G64gat), .B(G92gat), .ZN(new_n325));
  XOR2_X1   g124(.A(new_n324), .B(new_n325), .Z(new_n326));
  AOI21_X1  g125(.A(new_n288), .B1(new_n276), .B2(new_n278), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n327), .B1(new_n320), .B2(new_n312), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n265), .B1(new_n328), .B2(KEYINPUT29), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n266), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(new_n330), .A3(new_n263), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n323), .A2(new_n326), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT30), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT77), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n326), .ZN(new_n335));
  NOR3_X1   g134(.A1(new_n316), .A2(new_n264), .A3(new_n322), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n263), .B1(new_n329), .B2(new_n330), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n323), .A2(KEYINPUT30), .A3(new_n331), .A4(new_n326), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n334), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n332), .A2(KEYINPUT77), .A3(new_n333), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n247), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n332), .A2(new_n333), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT77), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n338), .A2(new_n339), .ZN(new_n347));
  AND4_X1   g146(.A1(new_n247), .A2(new_n346), .A3(new_n347), .A4(new_n342), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT31), .B(G50gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(G228gat), .A2(G233gat), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n352));
  NAND2_X1  g151(.A1(G155gat), .A2(G162gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT2), .ZN(new_n354));
  INV_X1    g153(.A(G155gat), .ZN(new_n355));
  INV_X1    g154(.A(G162gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI22_X1  g156(.A1(new_n352), .A2(new_n354), .B1(new_n357), .B2(new_n353), .ZN(new_n358));
  INV_X1    g157(.A(G148gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n359), .A2(G141gat), .ZN(new_n360));
  INV_X1    g159(.A(G141gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n361), .A2(G148gat), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n354), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n361), .A2(G148gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n359), .A2(G141gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n353), .ZN(new_n368));
  NOR2_X1   g167(.A1(G155gat), .A2(G162gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n354), .B(new_n367), .C1(new_n370), .C2(new_n352), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n364), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT3), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT29), .B1(new_n261), .B2(new_n262), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT81), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AOI211_X1 g175(.A(KEYINPUT81), .B(KEYINPUT29), .C1(new_n261), .C2(new_n262), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n372), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n364), .A2(new_n371), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT29), .B1(new_n379), .B2(new_n373), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(new_n263), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n351), .B1(new_n378), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n372), .B1(new_n374), .B2(KEYINPUT3), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n382), .A2(new_n351), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n350), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G78gat), .B(G106gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n388), .B(G22gat), .ZN(new_n389));
  INV_X1    g188(.A(new_n350), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n252), .A2(new_n254), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT75), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n252), .A2(new_n254), .A3(new_n255), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n259), .B1(new_n394), .B2(new_n250), .ZN(new_n395));
  INV_X1    g194(.A(new_n262), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n315), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT81), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n374), .A2(new_n375), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n373), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n381), .B1(new_n400), .B2(new_n372), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n385), .B(new_n390), .C1(new_n401), .C2(new_n351), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n387), .A2(new_n389), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n389), .B1(new_n387), .B2(new_n402), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n406));
  INV_X1    g205(.A(G134gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(G127gat), .ZN(new_n408));
  INV_X1    g207(.A(G127gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(G134gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT72), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT1), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT70), .ZN(new_n414));
  INV_X1    g213(.A(G113gat), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n414), .B1(new_n415), .B2(G120gat), .ZN(new_n416));
  INV_X1    g215(.A(G120gat), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n417), .A2(KEYINPUT70), .A3(G113gat), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n415), .A2(KEYINPUT71), .A3(G120gat), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT71), .B1(new_n415), .B2(G120gat), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n416), .B(new_n418), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(G127gat), .B(G134gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT72), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n413), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT68), .B(KEYINPUT69), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT68), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n426), .A2(G134gat), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n425), .B1(new_n422), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT69), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT68), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n426), .A2(KEYINPUT69), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n427), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n411), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT1), .ZN(new_n435));
  XOR2_X1   g234(.A(G113gat), .B(G120gat), .Z(new_n436));
  AOI22_X1  g235(.A1(new_n428), .A2(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n424), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n314), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n428), .A2(new_n434), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n436), .A2(new_n435), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n413), .A2(new_n421), .A3(new_n423), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n321), .A2(new_n444), .A3(new_n290), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n439), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(G227gat), .A2(G233gat), .ZN(new_n447));
  XOR2_X1   g246(.A(new_n447), .B(KEYINPUT64), .Z(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n406), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n406), .ZN(new_n451));
  AOI211_X1 g250(.A(new_n448), .B(new_n451), .C1(new_n439), .C2(new_n445), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n439), .A2(new_n448), .A3(new_n445), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT32), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT33), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g256(.A(G15gat), .B(G43gat), .Z(new_n458));
  XNOR2_X1  g257(.A(G71gat), .B(G99gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n458), .B(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n455), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n460), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n454), .B(KEYINPUT32), .C1(new_n456), .C2(new_n462), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n453), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n452), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n446), .A2(new_n449), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n451), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n461), .A2(new_n463), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT74), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n453), .A2(new_n461), .A3(new_n463), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT74), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(G1gat), .B(G29gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(KEYINPUT0), .ZN(new_n474));
  XNOR2_X1  g273(.A(G57gat), .B(G85gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n379), .A2(new_n373), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n364), .A2(new_n371), .A3(KEYINPUT3), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n477), .B(new_n478), .C1(new_n437), .C2(new_n424), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT5), .ZN(new_n480));
  NAND2_X1  g279(.A1(G225gat), .A2(G233gat), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n442), .A2(new_n379), .A3(new_n443), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT80), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT4), .ZN(new_n485));
  XNOR2_X1  g284(.A(KEYINPUT79), .B(KEYINPUT4), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n438), .A2(new_n379), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n484), .B1(new_n483), .B2(KEYINPUT4), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n482), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n372), .B1(new_n424), .B2(new_n437), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n483), .ZN(new_n494));
  INV_X1    g293(.A(new_n481), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n480), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n483), .A2(new_n486), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n442), .A2(KEYINPUT4), .A3(new_n379), .A4(new_n443), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n497), .A2(new_n479), .A3(new_n481), .A4(new_n498), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n476), .B1(new_n492), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT6), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n496), .A2(new_n499), .ZN(new_n503));
  INV_X1    g302(.A(new_n476), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n488), .A2(new_n490), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n503), .B(new_n504), .C1(new_n505), .C2(new_n482), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n501), .A2(new_n502), .A3(new_n506), .ZN(new_n507));
  OAI211_X1 g306(.A(KEYINPUT6), .B(new_n476), .C1(new_n492), .C2(new_n500), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT35), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n405), .A2(new_n469), .A3(new_n472), .A4(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n246), .B1(new_n349), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n405), .A2(new_n509), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n346), .A2(new_n347), .A3(new_n342), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT82), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n341), .A2(new_n247), .A3(new_n342), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n461), .A2(new_n463), .ZN(new_n517));
  INV_X1    g316(.A(new_n453), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n453), .A2(new_n461), .A3(new_n463), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n471), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n472), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n512), .A2(new_n516), .A3(KEYINPUT85), .A4(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n464), .A2(new_n468), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n405), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n507), .A2(new_n508), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n527), .A2(new_n342), .A3(new_n341), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT35), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n511), .A2(new_n524), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT40), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n531), .A2(KEYINPUT83), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n479), .B1(new_n488), .B2(new_n490), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT39), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(new_n535), .A3(new_n495), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n476), .B1(KEYINPUT83), .B2(new_n531), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(KEYINPUT39), .B1(new_n494), .B2(new_n495), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n539), .B1(new_n534), .B2(new_n495), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n533), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n534), .A2(new_n495), .ZN(new_n542));
  INV_X1    g341(.A(new_n539), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n544), .A2(new_n536), .A3(new_n537), .A4(new_n532), .ZN(new_n545));
  AND3_X1   g344(.A1(new_n541), .A2(new_n501), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n514), .A2(new_n546), .A3(new_n515), .ZN(new_n547));
  INV_X1    g346(.A(new_n527), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n323), .A2(new_n331), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n335), .B1(new_n549), .B2(KEYINPUT37), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n550), .A2(KEYINPUT38), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT37), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n552), .B1(new_n323), .B2(new_n331), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT84), .ZN(new_n554));
  OR2_X1    g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n554), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n551), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT38), .B1(new_n550), .B2(new_n553), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n548), .A2(new_n557), .A3(new_n332), .A4(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n547), .A2(new_n405), .A3(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n404), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n387), .A2(new_n389), .A3(new_n402), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n528), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n525), .A2(KEYINPUT36), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n565), .B1(new_n523), .B2(KEYINPUT36), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n560), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n245), .B1(new_n530), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT97), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT90), .ZN(new_n570));
  XOR2_X1   g369(.A(G57gat), .B(G64gat), .Z(new_n571));
  NAND2_X1  g370(.A1(G71gat), .A2(G78gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT9), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n572), .A2(KEYINPUT89), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n572), .A2(KEYINPUT89), .ZN(new_n577));
  OR2_X1    g376(.A1(G71gat), .A2(G78gat), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n570), .B1(new_n575), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n579), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n571), .A2(new_n574), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(KEYINPUT90), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n578), .A2(new_n572), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n575), .A2(KEYINPUT91), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n571), .A2(new_n574), .A3(new_n584), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT91), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n580), .A2(new_n583), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n589), .A2(KEYINPUT21), .ZN(new_n590));
  NAND2_X1  g389(.A1(G231gat), .A2(G233gat), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n590), .B(new_n592), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n593), .A2(new_n409), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n409), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n227), .B1(KEYINPUT21), .B2(new_n589), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n597), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n594), .A2(new_n595), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(new_n355), .ZN(new_n602));
  XNOR2_X1  g401(.A(G183gat), .B(G211gat), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n602), .B(new_n603), .Z(new_n604));
  AND3_X1   g403(.A1(new_n598), .A2(new_n600), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n604), .B1(new_n598), .B2(new_n600), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(G85gat), .ZN(new_n608));
  INV_X1    g407(.A(G92gat), .ZN(new_n609));
  OAI21_X1  g408(.A(KEYINPUT92), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT92), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n611), .A2(G85gat), .A3(G92gat), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n610), .A2(new_n612), .A3(KEYINPUT7), .ZN(new_n613));
  OR2_X1    g412(.A1(G99gat), .A2(G106gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(G99gat), .A2(G106gat), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n614), .A2(KEYINPUT96), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT7), .ZN(new_n617));
  OAI211_X1 g416(.A(KEYINPUT92), .B(new_n617), .C1(new_n608), .C2(new_n609), .ZN(new_n618));
  AND3_X1   g417(.A1(new_n613), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT8), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n620), .B1(new_n615), .B2(KEYINPUT93), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n621), .B1(KEYINPUT93), .B2(new_n615), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT95), .ZN(new_n623));
  OR2_X1    g422(.A1(KEYINPUT94), .A2(G85gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(KEYINPUT94), .A2(G85gat), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n624), .A2(new_n609), .A3(new_n625), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n622), .A2(new_n623), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n623), .B1(new_n622), .B2(new_n626), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n619), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n615), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n631), .A2(KEYINPUT96), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n632), .ZN(new_n634));
  OAI211_X1 g433(.A(new_n619), .B(new_n634), .C1(new_n627), .C2(new_n628), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n215), .A2(new_n224), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n213), .A2(new_n636), .ZN(new_n639));
  AND2_X1   g438(.A1(G232gat), .A2(G233gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(KEYINPUT41), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n638), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(G190gat), .B(G218gat), .Z(new_n643));
  OR2_X1    g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n640), .A2(KEYINPUT41), .ZN(new_n646));
  XNOR2_X1  g445(.A(G134gat), .B(G162gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n644), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n648), .B1(new_n644), .B2(new_n645), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n569), .B1(new_n607), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n651), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n598), .A2(new_n600), .ZN(new_n654));
  INV_X1    g453(.A(new_n604), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n598), .A2(new_n600), .A3(new_n604), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n653), .A2(new_n658), .A3(KEYINPUT97), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n652), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n622), .A2(new_n626), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(KEYINPUT95), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n622), .A2(new_n623), .A3(new_n626), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n634), .B1(new_n664), .B2(new_n619), .ZN(new_n665));
  INV_X1    g464(.A(new_n635), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n589), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT10), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n580), .A2(new_n583), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n585), .A2(new_n588), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n671), .A2(new_n633), .A3(new_n635), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n667), .A2(new_n668), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n636), .A2(KEYINPUT10), .A3(new_n589), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(G230gat), .A2(G233gat), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n676), .B1(new_n667), .B2(new_n672), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g479(.A(G120gat), .B(G148gat), .Z(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT98), .ZN(new_n682));
  XNOR2_X1  g481(.A(G176gat), .B(G204gat), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n682), .B(new_n683), .Z(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(KEYINPUT99), .B1(new_n680), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n676), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n687), .B1(new_n673), .B2(new_n674), .ZN(new_n688));
  NOR4_X1   g487(.A1(new_n688), .A2(KEYINPUT99), .A3(new_n678), .A4(new_n685), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n680), .A2(new_n685), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n660), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n568), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(new_n527), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(new_n218), .ZN(G1324gat));
  NAND3_X1  g496(.A1(new_n568), .A2(new_n349), .A3(new_n694), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  XOR2_X1   g498(.A(KEYINPUT16), .B(G8gat), .Z(new_n700));
  NAND3_X1  g499(.A1(new_n699), .A2(KEYINPUT42), .A3(new_n700), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n699), .A2(new_n700), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT42), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n703), .B1(new_n698), .B2(G8gat), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n701), .B(KEYINPUT100), .C1(new_n702), .C2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT101), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n701), .A2(KEYINPUT100), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n706), .B1(new_n705), .B2(new_n707), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(G1325gat));
  OR2_X1    g509(.A1(new_n566), .A2(KEYINPUT102), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n566), .A2(KEYINPUT102), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(G15gat), .B1(new_n695), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n523), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n716), .A2(G15gat), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n715), .B1(new_n695), .B2(new_n717), .ZN(G1326gat));
  AND2_X1   g517(.A1(new_n568), .A2(new_n563), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n694), .ZN(new_n720));
  XNOR2_X1  g519(.A(KEYINPUT43), .B(G22gat), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1327gat));
  AND2_X1   g521(.A1(new_n691), .A2(new_n692), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n607), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(new_n653), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n568), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(G29gat), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n726), .A2(new_n727), .A3(new_n548), .ZN(new_n728));
  XOR2_X1   g527(.A(KEYINPUT103), .B(KEYINPUT45), .Z(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n564), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n528), .A2(KEYINPUT104), .A3(new_n563), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n560), .A2(new_n566), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n653), .B1(new_n530), .B2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n530), .A2(new_n567), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n653), .A2(new_n738), .ZN(new_n740));
  AOI22_X1  g539(.A1(new_n737), .A2(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n724), .A2(new_n245), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n731), .B1(new_n743), .B2(new_n527), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(G29gat), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n743), .A2(new_n731), .A3(new_n527), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n730), .B1(new_n745), .B2(new_n746), .ZN(G1328gat));
  NOR2_X1   g546(.A1(new_n516), .A2(new_n204), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n726), .A2(new_n748), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(KEYINPUT46), .Z(new_n750));
  OAI21_X1  g549(.A(new_n204), .B1(new_n743), .B2(new_n516), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(G1329gat));
  OAI21_X1  g551(.A(G43gat), .B1(new_n743), .B2(new_n566), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n568), .A2(new_n725), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n754), .A2(G43gat), .A3(new_n716), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT47), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n741), .A2(new_n713), .A3(new_n742), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n755), .B1(new_n759), .B2(G43gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(KEYINPUT47), .B2(new_n760), .ZN(G1330gat));
  OAI21_X1  g560(.A(G50gat), .B1(new_n743), .B2(new_n405), .ZN(new_n762));
  INV_X1    g561(.A(G50gat), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n719), .A2(new_n763), .A3(new_n725), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(KEYINPUT106), .B(KEYINPUT48), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n765), .B(new_n767), .ZN(G1331gat));
  NAND2_X1  g567(.A1(new_n242), .A2(new_n244), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n660), .A2(new_n769), .A3(new_n723), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n530), .A2(new_n735), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n527), .B(KEYINPUT107), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g573(.A1(new_n770), .A2(new_n771), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n775), .A2(new_n516), .ZN(new_n776));
  NOR2_X1   g575(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n777));
  AND2_X1   g576(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(new_n776), .B2(new_n777), .ZN(G1333gat));
  OAI21_X1  g579(.A(G71gat), .B1(new_n775), .B2(new_n714), .ZN(new_n781));
  INV_X1    g580(.A(G71gat), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n523), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n775), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n785));
  XOR2_X1   g584(.A(new_n784), .B(new_n785), .Z(G1334gat));
  NOR2_X1   g585(.A1(new_n775), .A2(new_n405), .ZN(new_n787));
  XOR2_X1   g586(.A(KEYINPUT109), .B(G78gat), .Z(new_n788));
  XNOR2_X1  g587(.A(new_n787), .B(new_n788), .ZN(G1335gat));
  NAND2_X1  g588(.A1(new_n624), .A2(new_n625), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n739), .A2(new_n740), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n658), .A2(new_n723), .A3(new_n769), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n791), .B(new_n792), .C1(KEYINPUT44), .C2(new_n736), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n790), .B1(new_n793), .B2(new_n527), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n658), .A2(new_n769), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n771), .A2(new_n651), .A3(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n736), .A2(KEYINPUT51), .A3(new_n795), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n723), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n527), .A2(new_n790), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n794), .B1(new_n801), .B2(new_n802), .ZN(G1336gat));
  OAI21_X1  g602(.A(G92gat), .B1(new_n793), .B2(new_n516), .ZN(new_n804));
  XNOR2_X1  g603(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT111), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n516), .A2(G92gat), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n800), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n806), .B1(new_n800), .B2(new_n807), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n804), .B(new_n805), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT110), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n798), .A2(new_n811), .A3(new_n799), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT51), .B1(new_n736), .B2(new_n795), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT110), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n812), .A2(new_n693), .A3(new_n814), .A4(new_n807), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n804), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(KEYINPUT52), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n810), .A2(new_n817), .ZN(G1337gat));
  OAI21_X1  g617(.A(G99gat), .B1(new_n793), .B2(new_n714), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n716), .A2(G99gat), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n819), .B1(new_n801), .B2(new_n820), .ZN(G1338gat));
  NOR2_X1   g620(.A1(new_n405), .A2(G106gat), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n822), .A2(new_n693), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n812), .A2(new_n814), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(G106gat), .B1(new_n793), .B2(new_n405), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT53), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n736), .A2(KEYINPUT51), .A3(new_n795), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n693), .B(new_n822), .C1(new_n829), .C2(new_n813), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n825), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n827), .A2(new_n828), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n831), .B1(new_n824), .B2(new_n825), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n825), .A2(new_n830), .A3(new_n831), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT113), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n833), .A2(new_n836), .ZN(G1339gat));
  NAND3_X1  g636(.A1(new_n673), .A2(new_n674), .A3(new_n687), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n677), .A2(KEYINPUT54), .A3(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n684), .B1(new_n688), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n839), .A2(KEYINPUT55), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT99), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n688), .A2(new_n678), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n843), .B1(new_n844), .B2(new_n684), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n842), .B1(new_n845), .B2(new_n689), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT55), .B1(new_n839), .B2(new_n841), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT114), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n847), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT114), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n691), .A2(new_n849), .A3(new_n850), .A4(new_n842), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n848), .A2(new_n851), .A3(new_n769), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n225), .A2(new_n228), .ZN(new_n853));
  OAI22_X1  g652(.A1(new_n853), .A2(new_n226), .B1(new_n233), .B2(new_n234), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n240), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n693), .A2(new_n244), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n651), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n244), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n858), .A2(new_n649), .A3(new_n650), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n848), .A3(new_n851), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n607), .B1(new_n857), .B2(new_n861), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n652), .A2(new_n659), .A3(new_n245), .A4(new_n723), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n526), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n772), .A2(new_n516), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n867), .A2(G113gat), .A3(new_n245), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n563), .B1(new_n862), .B2(new_n863), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n516), .A2(new_n548), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n870), .A2(new_n716), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n769), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n868), .B1(new_n873), .B2(G113gat), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT115), .ZN(G1340gat));
  OR2_X1    g674(.A1(new_n867), .A2(new_n723), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n723), .A2(new_n417), .ZN(new_n877));
  AOI22_X1  g676(.A1(new_n876), .A2(new_n417), .B1(new_n872), .B2(new_n877), .ZN(G1341gat));
  NOR2_X1   g677(.A1(new_n867), .A2(new_n607), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n879), .A2(KEYINPUT116), .ZN(new_n880));
  AOI21_X1  g679(.A(G127gat), .B1(new_n879), .B2(KEYINPUT116), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n607), .A2(new_n409), .ZN(new_n882));
  AOI22_X1  g681(.A1(new_n880), .A2(new_n881), .B1(new_n872), .B2(new_n882), .ZN(G1342gat));
  NOR2_X1   g682(.A1(new_n653), .A2(G134gat), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n864), .A2(new_n865), .A3(new_n866), .A4(new_n884), .ZN(new_n885));
  XOR2_X1   g684(.A(new_n885), .B(KEYINPUT56), .Z(new_n886));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT117), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n869), .A2(new_n651), .A3(new_n871), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(G134gat), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n889), .A2(new_n888), .A3(G134gat), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n886), .B(new_n887), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n891), .A2(new_n890), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n885), .B(KEYINPUT56), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT118), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n892), .A2(new_n895), .ZN(G1343gat));
  INV_X1    g695(.A(new_n863), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n723), .A2(new_n858), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n691), .A2(new_n849), .A3(new_n842), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n245), .B1(KEYINPUT119), .B2(new_n899), .ZN(new_n900));
  OR3_X1    g699(.A1(new_n846), .A2(KEYINPUT119), .A3(new_n847), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n860), .B1(new_n902), .B2(new_n651), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n897), .B1(new_n903), .B2(new_n607), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT57), .B1(new_n904), .B2(new_n405), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n405), .B1(new_n862), .B2(new_n863), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT57), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n566), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(new_n870), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n905), .A2(new_n769), .A3(new_n908), .A4(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(G141gat), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n713), .A2(new_n405), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n864), .A2(new_n866), .A3(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(new_n361), .A3(new_n769), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(KEYINPUT58), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT58), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n912), .A2(new_n919), .A3(new_n916), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1344gat));
  NAND3_X1  g720(.A1(new_n915), .A2(new_n359), .A3(new_n693), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n359), .A2(KEYINPUT59), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n905), .A2(new_n908), .A3(new_n910), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n923), .B1(new_n925), .B2(new_n693), .ZN(new_n926));
  XOR2_X1   g725(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n927));
  NAND2_X1  g726(.A1(new_n899), .A2(KEYINPUT119), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n901), .A2(new_n928), .A3(new_n769), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n651), .B1(new_n929), .B2(new_n856), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n653), .A2(new_n858), .A3(new_n899), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n607), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n863), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n907), .A3(new_n563), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n909), .A2(new_n723), .A3(new_n870), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n934), .B(new_n935), .C1(new_n906), .C2(new_n907), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n927), .B1(new_n936), .B2(G148gat), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n922), .B1(new_n926), .B2(new_n937), .ZN(G1345gat));
  AOI21_X1  g737(.A(G155gat), .B1(new_n915), .B2(new_n658), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n658), .A2(G155gat), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT121), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n939), .B1(new_n925), .B2(new_n941), .ZN(G1346gat));
  OAI21_X1  g741(.A(new_n356), .B1(new_n914), .B2(new_n653), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n651), .A2(G162gat), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n924), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT122), .ZN(G1347gat));
  AOI21_X1  g745(.A(new_n548), .B1(new_n862), .B2(new_n863), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n349), .A2(new_n865), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT123), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(G169gat), .B1(new_n950), .B2(new_n769), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n716), .A2(new_n772), .A3(new_n516), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n869), .A2(new_n952), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n953), .A2(new_n280), .A3(new_n245), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n951), .A2(new_n954), .ZN(G1348gat));
  NAND3_X1  g754(.A1(new_n950), .A2(new_n281), .A3(new_n693), .ZN(new_n956));
  OAI21_X1  g755(.A(G176gat), .B1(new_n953), .B2(new_n723), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(G1349gat));
  INV_X1    g757(.A(KEYINPUT125), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n959), .A2(KEYINPUT60), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n959), .A2(KEYINPUT60), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n864), .A2(new_n405), .A3(new_n658), .A4(new_n952), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(KEYINPUT124), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT124), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n869), .A2(new_n964), .A3(new_n658), .A4(new_n952), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n963), .A2(G183gat), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n950), .A2(new_n277), .A3(new_n658), .ZN(new_n967));
  AOI211_X1 g766(.A(new_n960), .B(new_n961), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  AND4_X1   g767(.A1(new_n959), .A2(new_n966), .A3(KEYINPUT60), .A4(new_n967), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n968), .A2(new_n969), .ZN(G1350gat));
  NAND3_X1  g769(.A1(new_n950), .A2(new_n274), .A3(new_n651), .ZN(new_n971));
  OAI21_X1  g770(.A(G190gat), .B1(new_n953), .B2(new_n653), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n972), .A2(KEYINPUT61), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n972), .A2(KEYINPUT61), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n971), .B1(new_n973), .B2(new_n974), .ZN(G1351gat));
  OAI211_X1 g774(.A(new_n934), .B(KEYINPUT126), .C1(new_n906), .C2(new_n907), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n977));
  AOI211_X1 g776(.A(KEYINPUT57), .B(new_n405), .C1(new_n932), .C2(new_n863), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n906), .A2(new_n907), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NOR3_X1   g779(.A1(new_n713), .A2(new_n516), .A3(new_n772), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n245), .A2(new_n253), .ZN(new_n982));
  NAND4_X1  g781(.A1(new_n976), .A2(new_n980), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  NOR3_X1   g782(.A1(new_n713), .A2(new_n405), .A3(new_n516), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n947), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n253), .B1(new_n985), .B2(new_n245), .ZN(new_n986));
  AND2_X1   g785(.A1(new_n983), .A2(new_n986), .ZN(G1352gat));
  NOR3_X1   g786(.A1(new_n985), .A2(G204gat), .A3(new_n723), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n988), .B(KEYINPUT62), .ZN(new_n989));
  AND4_X1   g788(.A1(new_n693), .A2(new_n976), .A3(new_n980), .A4(new_n981), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n989), .B1(new_n990), .B2(new_n251), .ZN(G1353gat));
  INV_X1    g790(.A(G211gat), .ZN(new_n992));
  NAND4_X1  g791(.A1(new_n947), .A2(new_n992), .A3(new_n658), .A4(new_n984), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT127), .ZN(new_n994));
  AND2_X1   g793(.A1(new_n981), .A2(new_n658), .ZN(new_n995));
  OAI211_X1 g794(.A(new_n934), .B(new_n995), .C1(new_n906), .C2(new_n907), .ZN(new_n996));
  AND4_X1   g795(.A1(new_n994), .A2(new_n996), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT63), .ZN(new_n998));
  AOI21_X1  g797(.A(new_n992), .B1(KEYINPUT127), .B2(new_n998), .ZN(new_n999));
  AOI22_X1  g798(.A1(new_n996), .A2(new_n999), .B1(new_n994), .B2(KEYINPUT63), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n993), .B1(new_n997), .B2(new_n1000), .ZN(G1354gat));
  INV_X1    g800(.A(G218gat), .ZN(new_n1002));
  NOR2_X1   g801(.A1(new_n653), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g802(.A1(new_n976), .A2(new_n980), .A3(new_n981), .A4(new_n1003), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n1002), .B1(new_n985), .B2(new_n653), .ZN(new_n1005));
  AND2_X1   g804(.A1(new_n1004), .A2(new_n1005), .ZN(G1355gat));
endmodule


