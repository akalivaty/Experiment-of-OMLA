

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U550 ( .A(KEYINPUT75), .B(n580), .Z(n954) );
  AND2_X1 U551 ( .A1(n954), .A2(n701), .ZN(n685) );
  INV_X1 U552 ( .A(n951), .ZN(n756) );
  NOR2_X1 U553 ( .A1(n757), .A2(n756), .ZN(n514) );
  NAND2_X1 U554 ( .A1(n753), .A2(n752), .ZN(n515) );
  NOR2_X1 U555 ( .A1(n694), .A2(n693), .ZN(n705) );
  NOR2_X1 U556 ( .A1(n708), .A2(n707), .ZN(n709) );
  INV_X1 U557 ( .A(KEYINPUT29), .ZN(n711) );
  XNOR2_X1 U558 ( .A(n712), .B(n711), .ZN(n718) );
  INV_X1 U559 ( .A(KEYINPUT103), .ZN(n737) );
  XNOR2_X1 U560 ( .A(n738), .B(n737), .ZN(n739) );
  XOR2_X1 U561 ( .A(n680), .B(KEYINPUT64), .Z(n713) );
  INV_X1 U562 ( .A(n713), .ZN(n720) );
  NOR2_X1 U563 ( .A1(G164), .A2(G1384), .ZN(n789) );
  NOR2_X1 U564 ( .A1(G651), .A2(n620), .ZN(n630) );
  XOR2_X1 U565 ( .A(KEYINPUT1), .B(n527), .Z(n635) );
  AND2_X1 U566 ( .A1(n823), .A2(n822), .ZN(n824) );
  NOR2_X1 U567 ( .A1(n526), .A2(n525), .ZN(G164) );
  NAND2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n516) );
  XOR2_X2 U569 ( .A(KEYINPUT66), .B(n516), .Z(n891) );
  NAND2_X1 U570 ( .A1(G114), .A2(n891), .ZN(n518) );
  INV_X1 U571 ( .A(G2105), .ZN(n522) );
  NOR2_X2 U572 ( .A1(G2104), .A2(n522), .ZN(n890) );
  NAND2_X1 U573 ( .A1(G126), .A2(n890), .ZN(n517) );
  NAND2_X1 U574 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U575 ( .A(n519), .B(KEYINPUT92), .ZN(n526) );
  XNOR2_X1 U576 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n521) );
  NOR2_X1 U577 ( .A1(G2104), .A2(G2105), .ZN(n520) );
  XNOR2_X1 U578 ( .A(n521), .B(n520), .ZN(n886) );
  NAND2_X1 U579 ( .A1(G138), .A2(n886), .ZN(n524) );
  AND2_X1 U580 ( .A1(n522), .A2(G2104), .ZN(n887) );
  NAND2_X1 U581 ( .A1(G102), .A2(n887), .ZN(n523) );
  NAND2_X1 U582 ( .A1(n524), .A2(n523), .ZN(n525) );
  INV_X1 U583 ( .A(G651), .ZN(n533) );
  NOR2_X1 U584 ( .A1(G543), .A2(n533), .ZN(n527) );
  NAND2_X1 U585 ( .A1(n635), .A2(G63), .ZN(n528) );
  XNOR2_X1 U586 ( .A(n528), .B(KEYINPUT78), .ZN(n530) );
  XOR2_X1 U587 ( .A(G543), .B(KEYINPUT0), .Z(n620) );
  NAND2_X1 U588 ( .A1(G51), .A2(n630), .ZN(n529) );
  NAND2_X1 U589 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U590 ( .A(KEYINPUT6), .B(n531), .ZN(n540) );
  NOR2_X1 U591 ( .A1(G651), .A2(G543), .ZN(n631) );
  NAND2_X1 U592 ( .A1(n631), .A2(G89), .ZN(n532) );
  XOR2_X1 U593 ( .A(KEYINPUT4), .B(n532), .Z(n536) );
  NOR2_X1 U594 ( .A1(n620), .A2(n533), .ZN(n632) );
  NAND2_X1 U595 ( .A1(n632), .A2(G76), .ZN(n534) );
  XOR2_X1 U596 ( .A(n534), .B(KEYINPUT76), .Z(n535) );
  NOR2_X1 U597 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U598 ( .A(KEYINPUT77), .B(n537), .Z(n538) );
  XNOR2_X1 U599 ( .A(n538), .B(KEYINPUT5), .ZN(n539) );
  NOR2_X1 U600 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U601 ( .A(n541), .B(KEYINPUT7), .ZN(n542) );
  XNOR2_X1 U602 ( .A(n542), .B(KEYINPUT79), .ZN(G168) );
  XOR2_X1 U603 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U604 ( .A1(G85), .A2(n631), .ZN(n544) );
  NAND2_X1 U605 ( .A1(G72), .A2(n632), .ZN(n543) );
  NAND2_X1 U606 ( .A1(n544), .A2(n543), .ZN(n548) );
  NAND2_X1 U607 ( .A1(G60), .A2(n635), .ZN(n546) );
  NAND2_X1 U608 ( .A1(G47), .A2(n630), .ZN(n545) );
  NAND2_X1 U609 ( .A1(n546), .A2(n545), .ZN(n547) );
  OR2_X1 U610 ( .A1(n548), .A2(n547), .ZN(G290) );
  INV_X1 U611 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U612 ( .A(KEYINPUT9), .B(KEYINPUT69), .ZN(n552) );
  NAND2_X1 U613 ( .A1(G90), .A2(n631), .ZN(n550) );
  NAND2_X1 U614 ( .A1(G77), .A2(n632), .ZN(n549) );
  NAND2_X1 U615 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n552), .B(n551), .ZN(n557) );
  NAND2_X1 U617 ( .A1(n635), .A2(G64), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n553), .B(KEYINPUT68), .ZN(n555) );
  NAND2_X1 U619 ( .A1(G52), .A2(n630), .ZN(n554) );
  NAND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U621 ( .A1(n557), .A2(n556), .ZN(G171) );
  NAND2_X1 U622 ( .A1(G94), .A2(G452), .ZN(n558) );
  XOR2_X1 U623 ( .A(KEYINPUT70), .B(n558), .Z(G173) );
  NAND2_X1 U624 ( .A1(G7), .A2(G661), .ZN(n559) );
  XOR2_X1 U625 ( .A(n559), .B(KEYINPUT10), .Z(n836) );
  NAND2_X1 U626 ( .A1(n836), .A2(G567), .ZN(n560) );
  XOR2_X1 U627 ( .A(KEYINPUT11), .B(n560), .Z(G234) );
  NAND2_X1 U628 ( .A1(G56), .A2(n635), .ZN(n561) );
  XOR2_X1 U629 ( .A(KEYINPUT14), .B(n561), .Z(n568) );
  NAND2_X1 U630 ( .A1(G81), .A2(n631), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n562), .B(KEYINPUT12), .ZN(n563) );
  XNOR2_X1 U632 ( .A(n563), .B(KEYINPUT72), .ZN(n565) );
  NAND2_X1 U633 ( .A1(G68), .A2(n632), .ZN(n564) );
  NAND2_X1 U634 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U635 ( .A(KEYINPUT13), .B(n566), .Z(n567) );
  NOR2_X1 U636 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U637 ( .A1(n630), .A2(G43), .ZN(n569) );
  NAND2_X1 U638 ( .A1(n570), .A2(n569), .ZN(n948) );
  INV_X1 U639 ( .A(G860), .ZN(n592) );
  OR2_X1 U640 ( .A1(n948), .A2(n592), .ZN(G153) );
  INV_X1 U641 ( .A(G868), .ZN(n653) );
  NOR2_X1 U642 ( .A1(n653), .A2(G171), .ZN(n571) );
  XNOR2_X1 U643 ( .A(n571), .B(KEYINPUT73), .ZN(n582) );
  NAND2_X1 U644 ( .A1(G54), .A2(n630), .ZN(n578) );
  NAND2_X1 U645 ( .A1(G92), .A2(n631), .ZN(n573) );
  NAND2_X1 U646 ( .A1(G79), .A2(n632), .ZN(n572) );
  NAND2_X1 U647 ( .A1(n573), .A2(n572), .ZN(n576) );
  NAND2_X1 U648 ( .A1(n635), .A2(G66), .ZN(n574) );
  XOR2_X1 U649 ( .A(KEYINPUT74), .B(n574), .Z(n575) );
  NOR2_X1 U650 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U651 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U652 ( .A(n579), .B(KEYINPUT15), .ZN(n580) );
  INV_X1 U653 ( .A(n954), .ZN(n699) );
  NAND2_X1 U654 ( .A1(n653), .A2(n699), .ZN(n581) );
  NAND2_X1 U655 ( .A1(n582), .A2(n581), .ZN(G284) );
  NAND2_X1 U656 ( .A1(G91), .A2(n631), .ZN(n584) );
  NAND2_X1 U657 ( .A1(G78), .A2(n632), .ZN(n583) );
  NAND2_X1 U658 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U659 ( .A(KEYINPUT71), .B(n585), .ZN(n589) );
  NAND2_X1 U660 ( .A1(G65), .A2(n635), .ZN(n587) );
  NAND2_X1 U661 ( .A1(G53), .A2(n630), .ZN(n586) );
  AND2_X1 U662 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U663 ( .A1(n589), .A2(n588), .ZN(G299) );
  NOR2_X1 U664 ( .A1(G286), .A2(n653), .ZN(n591) );
  NOR2_X1 U665 ( .A1(G868), .A2(G299), .ZN(n590) );
  NOR2_X1 U666 ( .A1(n591), .A2(n590), .ZN(G297) );
  NAND2_X1 U667 ( .A1(n592), .A2(G559), .ZN(n593) );
  NAND2_X1 U668 ( .A1(n593), .A2(n954), .ZN(n594) );
  XNOR2_X1 U669 ( .A(n594), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U670 ( .A1(G868), .A2(n948), .ZN(n597) );
  NAND2_X1 U671 ( .A1(G868), .A2(n954), .ZN(n595) );
  NOR2_X1 U672 ( .A1(G559), .A2(n595), .ZN(n596) );
  NOR2_X1 U673 ( .A1(n597), .A2(n596), .ZN(G282) );
  NAND2_X1 U674 ( .A1(G99), .A2(n887), .ZN(n598) );
  XNOR2_X1 U675 ( .A(n598), .B(KEYINPUT80), .ZN(n605) );
  NAND2_X1 U676 ( .A1(n886), .A2(G135), .ZN(n600) );
  NAND2_X1 U677 ( .A1(G111), .A2(n891), .ZN(n599) );
  NAND2_X1 U678 ( .A1(n600), .A2(n599), .ZN(n603) );
  NAND2_X1 U679 ( .A1(n890), .A2(G123), .ZN(n601) );
  XOR2_X1 U680 ( .A(KEYINPUT18), .B(n601), .Z(n602) );
  NOR2_X1 U681 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U682 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U683 ( .A(KEYINPUT81), .B(n606), .ZN(n926) );
  XNOR2_X1 U684 ( .A(n926), .B(G2096), .ZN(n607) );
  INV_X1 U685 ( .A(G2100), .ZN(n863) );
  NAND2_X1 U686 ( .A1(n607), .A2(n863), .ZN(G156) );
  NAND2_X1 U687 ( .A1(G67), .A2(n635), .ZN(n609) );
  NAND2_X1 U688 ( .A1(G93), .A2(n631), .ZN(n608) );
  NAND2_X1 U689 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U690 ( .A1(G80), .A2(n632), .ZN(n611) );
  NAND2_X1 U691 ( .A1(G55), .A2(n630), .ZN(n610) );
  NAND2_X1 U692 ( .A1(n611), .A2(n610), .ZN(n612) );
  OR2_X1 U693 ( .A1(n613), .A2(n612), .ZN(n652) );
  NAND2_X1 U694 ( .A1(G559), .A2(n954), .ZN(n614) );
  XOR2_X1 U695 ( .A(n948), .B(n614), .Z(n650) );
  XOR2_X1 U696 ( .A(n650), .B(KEYINPUT82), .Z(n615) );
  NOR2_X1 U697 ( .A1(G860), .A2(n615), .ZN(n616) );
  XOR2_X1 U698 ( .A(n652), .B(n616), .Z(G145) );
  NAND2_X1 U699 ( .A1(G49), .A2(n630), .ZN(n618) );
  NAND2_X1 U700 ( .A1(G74), .A2(G651), .ZN(n617) );
  NAND2_X1 U701 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U702 ( .A1(n635), .A2(n619), .ZN(n622) );
  NAND2_X1 U703 ( .A1(n620), .A2(G87), .ZN(n621) );
  NAND2_X1 U704 ( .A1(n622), .A2(n621), .ZN(G288) );
  NAND2_X1 U705 ( .A1(G61), .A2(n635), .ZN(n624) );
  NAND2_X1 U706 ( .A1(G86), .A2(n631), .ZN(n623) );
  NAND2_X1 U707 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U708 ( .A1(n632), .A2(G73), .ZN(n625) );
  XOR2_X1 U709 ( .A(KEYINPUT2), .B(n625), .Z(n626) );
  NOR2_X1 U710 ( .A1(n627), .A2(n626), .ZN(n629) );
  NAND2_X1 U711 ( .A1(n630), .A2(G48), .ZN(n628) );
  NAND2_X1 U712 ( .A1(n629), .A2(n628), .ZN(G305) );
  NAND2_X1 U713 ( .A1(n630), .A2(G50), .ZN(n640) );
  NAND2_X1 U714 ( .A1(G88), .A2(n631), .ZN(n634) );
  NAND2_X1 U715 ( .A1(G75), .A2(n632), .ZN(n633) );
  NAND2_X1 U716 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U717 ( .A1(G62), .A2(n635), .ZN(n636) );
  XNOR2_X1 U718 ( .A(KEYINPUT83), .B(n636), .ZN(n637) );
  NOR2_X1 U719 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U721 ( .A(KEYINPUT84), .B(n641), .ZN(G303) );
  XOR2_X1 U722 ( .A(KEYINPUT85), .B(KEYINPUT19), .Z(n642) );
  XNOR2_X1 U723 ( .A(G288), .B(n642), .ZN(n643) );
  XNOR2_X1 U724 ( .A(KEYINPUT87), .B(n643), .ZN(n645) );
  XNOR2_X1 U725 ( .A(G305), .B(KEYINPUT86), .ZN(n644) );
  XNOR2_X1 U726 ( .A(n645), .B(n644), .ZN(n646) );
  XOR2_X1 U727 ( .A(n652), .B(n646), .Z(n648) );
  XOR2_X1 U728 ( .A(G290), .B(G299), .Z(n647) );
  XNOR2_X1 U729 ( .A(n648), .B(n647), .ZN(n649) );
  XOR2_X1 U730 ( .A(n649), .B(G303), .Z(n909) );
  XNOR2_X1 U731 ( .A(n650), .B(n909), .ZN(n651) );
  NAND2_X1 U732 ( .A1(n651), .A2(G868), .ZN(n655) );
  NAND2_X1 U733 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U734 ( .A1(n655), .A2(n654), .ZN(G295) );
  NAND2_X1 U735 ( .A1(G2078), .A2(G2084), .ZN(n656) );
  XOR2_X1 U736 ( .A(KEYINPUT20), .B(n656), .Z(n657) );
  NAND2_X1 U737 ( .A1(G2090), .A2(n657), .ZN(n658) );
  XNOR2_X1 U738 ( .A(KEYINPUT21), .B(n658), .ZN(n659) );
  NAND2_X1 U739 ( .A1(n659), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U740 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U741 ( .A1(G69), .A2(G120), .ZN(n660) );
  XNOR2_X1 U742 ( .A(KEYINPUT90), .B(n660), .ZN(n661) );
  NOR2_X1 U743 ( .A1(G238), .A2(n661), .ZN(n662) );
  NAND2_X1 U744 ( .A1(G57), .A2(n662), .ZN(n841) );
  NAND2_X1 U745 ( .A1(n841), .A2(G567), .ZN(n669) );
  NAND2_X1 U746 ( .A1(G132), .A2(G82), .ZN(n663) );
  XNOR2_X1 U747 ( .A(n663), .B(KEYINPUT22), .ZN(n664) );
  XNOR2_X1 U748 ( .A(n664), .B(KEYINPUT88), .ZN(n665) );
  NOR2_X1 U749 ( .A1(G218), .A2(n665), .ZN(n666) );
  XOR2_X1 U750 ( .A(KEYINPUT89), .B(n666), .Z(n667) );
  NAND2_X1 U751 ( .A1(G96), .A2(n667), .ZN(n842) );
  NAND2_X1 U752 ( .A1(n842), .A2(G2106), .ZN(n668) );
  NAND2_X1 U753 ( .A1(n669), .A2(n668), .ZN(n843) );
  NAND2_X1 U754 ( .A1(G483), .A2(G661), .ZN(n670) );
  NOR2_X1 U755 ( .A1(n843), .A2(n670), .ZN(n671) );
  XOR2_X1 U756 ( .A(KEYINPUT91), .B(n671), .Z(n840) );
  NAND2_X1 U757 ( .A1(n840), .A2(G36), .ZN(G176) );
  NAND2_X1 U758 ( .A1(n886), .A2(G137), .ZN(n674) );
  NAND2_X1 U759 ( .A1(G101), .A2(n887), .ZN(n672) );
  XOR2_X1 U760 ( .A(KEYINPUT23), .B(n672), .Z(n673) );
  NAND2_X1 U761 ( .A1(n674), .A2(n673), .ZN(n678) );
  NAND2_X1 U762 ( .A1(G125), .A2(n890), .ZN(n676) );
  NAND2_X1 U763 ( .A1(G113), .A2(n891), .ZN(n675) );
  NAND2_X1 U764 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U765 ( .A1(n678), .A2(n677), .ZN(G160) );
  NAND2_X1 U766 ( .A1(G160), .A2(G40), .ZN(n788) );
  INV_X1 U767 ( .A(n788), .ZN(n679) );
  NAND2_X1 U768 ( .A1(n679), .A2(n789), .ZN(n680) );
  NAND2_X1 U769 ( .A1(n720), .A2(G1341), .ZN(n681) );
  XOR2_X1 U770 ( .A(KEYINPUT100), .B(n681), .Z(n682) );
  NOR2_X1 U771 ( .A1(n948), .A2(n682), .ZN(n700) );
  XOR2_X1 U772 ( .A(KEYINPUT65), .B(KEYINPUT26), .Z(n684) );
  NAND2_X1 U773 ( .A1(G1996), .A2(n713), .ZN(n683) );
  XNOR2_X1 U774 ( .A(n684), .B(n683), .ZN(n701) );
  NAND2_X1 U775 ( .A1(n700), .A2(n685), .ZN(n687) );
  INV_X1 U776 ( .A(KEYINPUT101), .ZN(n686) );
  XNOR2_X1 U777 ( .A(n687), .B(n686), .ZN(n697) );
  NOR2_X1 U778 ( .A1(G2067), .A2(n720), .ZN(n689) );
  NOR2_X1 U779 ( .A1(G1348), .A2(n713), .ZN(n688) );
  NOR2_X1 U780 ( .A1(n689), .A2(n688), .ZN(n695) );
  NAND2_X1 U781 ( .A1(n720), .A2(G1956), .ZN(n690) );
  XNOR2_X1 U782 ( .A(KEYINPUT99), .B(n690), .ZN(n694) );
  AND2_X1 U783 ( .A1(G2072), .A2(n713), .ZN(n692) );
  INV_X1 U784 ( .A(KEYINPUT27), .ZN(n691) );
  XNOR2_X1 U785 ( .A(n692), .B(n691), .ZN(n693) );
  INV_X1 U786 ( .A(G299), .ZN(n704) );
  NAND2_X1 U787 ( .A1(n705), .A2(n704), .ZN(n698) );
  AND2_X1 U788 ( .A1(n695), .A2(n698), .ZN(n696) );
  NAND2_X1 U789 ( .A1(n697), .A2(n696), .ZN(n710) );
  AND2_X1 U790 ( .A1(n699), .A2(n698), .ZN(n703) );
  NAND2_X1 U791 ( .A1(n701), .A2(n700), .ZN(n702) );
  AND2_X1 U792 ( .A1(n703), .A2(n702), .ZN(n708) );
  NOR2_X1 U793 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U794 ( .A(n706), .B(KEYINPUT28), .ZN(n707) );
  NAND2_X1 U795 ( .A1(n710), .A2(n709), .ZN(n712) );
  XNOR2_X1 U796 ( .A(G2078), .B(KEYINPUT25), .ZN(n995) );
  NAND2_X1 U797 ( .A1(n713), .A2(n995), .ZN(n715) );
  INV_X1 U798 ( .A(G1961), .ZN(n844) );
  NAND2_X1 U799 ( .A1(n720), .A2(n844), .ZN(n714) );
  NAND2_X1 U800 ( .A1(n715), .A2(n714), .ZN(n725) );
  AND2_X1 U801 ( .A1(n725), .A2(G171), .ZN(n716) );
  XOR2_X1 U802 ( .A(KEYINPUT98), .B(n716), .Z(n717) );
  NAND2_X1 U803 ( .A1(n718), .A2(n717), .ZN(n730) );
  INV_X1 U804 ( .A(G8), .ZN(n731) );
  OR2_X1 U805 ( .A1(G1966), .A2(n731), .ZN(n719) );
  NOR2_X1 U806 ( .A1(n713), .A2(n719), .ZN(n743) );
  NOR2_X1 U807 ( .A1(n720), .A2(G2084), .ZN(n744) );
  NOR2_X1 U808 ( .A1(n743), .A2(n744), .ZN(n721) );
  NAND2_X1 U809 ( .A1(G8), .A2(n721), .ZN(n722) );
  XNOR2_X1 U810 ( .A(KEYINPUT102), .B(n722), .ZN(n723) );
  XNOR2_X1 U811 ( .A(KEYINPUT30), .B(n723), .ZN(n724) );
  NOR2_X1 U812 ( .A1(n724), .A2(G168), .ZN(n727) );
  NOR2_X1 U813 ( .A1(G171), .A2(n725), .ZN(n726) );
  NOR2_X1 U814 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U815 ( .A(n728), .B(KEYINPUT31), .Z(n729) );
  NAND2_X1 U816 ( .A1(n730), .A2(n729), .ZN(n741) );
  NAND2_X1 U817 ( .A1(n741), .A2(G286), .ZN(n736) );
  NOR2_X1 U818 ( .A1(n720), .A2(G2090), .ZN(n733) );
  OR2_X1 U819 ( .A1(n713), .A2(n731), .ZN(n769) );
  NOR2_X1 U820 ( .A1(G1971), .A2(n769), .ZN(n732) );
  NOR2_X1 U821 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U822 ( .A1(G303), .A2(n734), .ZN(n735) );
  NAND2_X1 U823 ( .A1(n736), .A2(n735), .ZN(n738) );
  NAND2_X1 U824 ( .A1(G8), .A2(n739), .ZN(n740) );
  XNOR2_X1 U825 ( .A(n740), .B(KEYINPUT32), .ZN(n759) );
  INV_X1 U826 ( .A(n741), .ZN(n742) );
  NOR2_X1 U827 ( .A1(n743), .A2(n742), .ZN(n746) );
  NAND2_X1 U828 ( .A1(G8), .A2(n744), .ZN(n745) );
  NAND2_X1 U829 ( .A1(n746), .A2(n745), .ZN(n758) );
  NAND2_X1 U830 ( .A1(G1976), .A2(G288), .ZN(n961) );
  AND2_X1 U831 ( .A1(n758), .A2(n961), .ZN(n747) );
  NAND2_X1 U832 ( .A1(n759), .A2(n747), .ZN(n753) );
  INV_X1 U833 ( .A(n961), .ZN(n749) );
  NOR2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n754) );
  NOR2_X1 U835 ( .A1(G303), .A2(G1971), .ZN(n748) );
  NOR2_X1 U836 ( .A1(n754), .A2(n748), .ZN(n958) );
  OR2_X1 U837 ( .A1(n749), .A2(n958), .ZN(n750) );
  NOR2_X1 U838 ( .A1(n769), .A2(n750), .ZN(n751) );
  NOR2_X1 U839 ( .A1(n751), .A2(KEYINPUT33), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n754), .A2(KEYINPUT33), .ZN(n755) );
  NOR2_X1 U841 ( .A1(n755), .A2(n769), .ZN(n757) );
  XOR2_X1 U842 ( .A(G1981), .B(G305), .Z(n951) );
  NAND2_X1 U843 ( .A1(n515), .A2(n514), .ZN(n765) );
  NAND2_X1 U844 ( .A1(n759), .A2(n758), .ZN(n762) );
  NOR2_X1 U845 ( .A1(G2090), .A2(G303), .ZN(n760) );
  NAND2_X1 U846 ( .A1(G8), .A2(n760), .ZN(n761) );
  NAND2_X1 U847 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U848 ( .A1(n763), .A2(n769), .ZN(n764) );
  NAND2_X1 U849 ( .A1(n765), .A2(n764), .ZN(n813) );
  NOR2_X1 U850 ( .A1(G1981), .A2(G305), .ZN(n766) );
  XOR2_X1 U851 ( .A(n766), .B(KEYINPUT24), .Z(n767) );
  XNOR2_X1 U852 ( .A(KEYINPUT96), .B(n767), .ZN(n768) );
  NOR2_X1 U853 ( .A1(n769), .A2(n768), .ZN(n770) );
  XOR2_X1 U854 ( .A(KEYINPUT97), .B(n770), .Z(n811) );
  NAND2_X1 U855 ( .A1(G129), .A2(n890), .ZN(n772) );
  NAND2_X1 U856 ( .A1(G141), .A2(n886), .ZN(n771) );
  NAND2_X1 U857 ( .A1(n772), .A2(n771), .ZN(n775) );
  NAND2_X1 U858 ( .A1(n887), .A2(G105), .ZN(n773) );
  XOR2_X1 U859 ( .A(KEYINPUT38), .B(n773), .Z(n774) );
  NOR2_X1 U860 ( .A1(n775), .A2(n774), .ZN(n777) );
  NAND2_X1 U861 ( .A1(G117), .A2(n891), .ZN(n776) );
  NAND2_X1 U862 ( .A1(n777), .A2(n776), .ZN(n898) );
  NOR2_X1 U863 ( .A1(G1996), .A2(n898), .ZN(n939) );
  NAND2_X1 U864 ( .A1(G131), .A2(n886), .ZN(n778) );
  XNOR2_X1 U865 ( .A(n778), .B(KEYINPUT94), .ZN(n781) );
  NAND2_X1 U866 ( .A1(G95), .A2(n887), .ZN(n779) );
  XOR2_X1 U867 ( .A(KEYINPUT93), .B(n779), .Z(n780) );
  NAND2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n785) );
  NAND2_X1 U869 ( .A1(G119), .A2(n890), .ZN(n783) );
  NAND2_X1 U870 ( .A1(G107), .A2(n891), .ZN(n782) );
  NAND2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n897) );
  INV_X1 U873 ( .A(G1991), .ZN(n848) );
  NOR2_X1 U874 ( .A1(n897), .A2(n848), .ZN(n787) );
  AND2_X1 U875 ( .A1(G1996), .A2(n898), .ZN(n786) );
  NOR2_X1 U876 ( .A1(n787), .A2(n786), .ZN(n929) );
  NOR2_X1 U877 ( .A1(n789), .A2(n788), .ZN(n817) );
  XNOR2_X1 U878 ( .A(KEYINPUT95), .B(n817), .ZN(n790) );
  NOR2_X1 U879 ( .A1(n929), .A2(n790), .ZN(n814) );
  AND2_X1 U880 ( .A1(n848), .A2(n897), .ZN(n925) );
  NOR2_X1 U881 ( .A1(G1986), .A2(G290), .ZN(n791) );
  XNOR2_X1 U882 ( .A(KEYINPUT104), .B(n791), .ZN(n792) );
  NOR2_X1 U883 ( .A1(n925), .A2(n792), .ZN(n793) );
  NOR2_X1 U884 ( .A1(n814), .A2(n793), .ZN(n794) );
  XOR2_X1 U885 ( .A(KEYINPUT105), .B(n794), .Z(n795) );
  NOR2_X1 U886 ( .A1(n939), .A2(n795), .ZN(n796) );
  XNOR2_X1 U887 ( .A(n796), .B(KEYINPUT39), .ZN(n806) );
  NAND2_X1 U888 ( .A1(G140), .A2(n886), .ZN(n798) );
  NAND2_X1 U889 ( .A1(G104), .A2(n887), .ZN(n797) );
  NAND2_X1 U890 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U891 ( .A(KEYINPUT34), .B(n799), .ZN(n804) );
  NAND2_X1 U892 ( .A1(G128), .A2(n890), .ZN(n801) );
  NAND2_X1 U893 ( .A1(G116), .A2(n891), .ZN(n800) );
  NAND2_X1 U894 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U895 ( .A(KEYINPUT35), .B(n802), .Z(n803) );
  NOR2_X1 U896 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U897 ( .A(KEYINPUT36), .B(n805), .ZN(n903) );
  XNOR2_X1 U898 ( .A(KEYINPUT37), .B(G2067), .ZN(n807) );
  NOR2_X1 U899 ( .A1(n903), .A2(n807), .ZN(n923) );
  NAND2_X1 U900 ( .A1(n817), .A2(n923), .ZN(n816) );
  NAND2_X1 U901 ( .A1(n806), .A2(n816), .ZN(n808) );
  NAND2_X1 U902 ( .A1(n903), .A2(n807), .ZN(n922) );
  NAND2_X1 U903 ( .A1(n808), .A2(n922), .ZN(n809) );
  XNOR2_X1 U904 ( .A(KEYINPUT106), .B(n809), .ZN(n810) );
  AND2_X1 U905 ( .A1(n810), .A2(n817), .ZN(n821) );
  OR2_X1 U906 ( .A1(n811), .A2(n821), .ZN(n812) );
  OR2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n823) );
  INV_X1 U908 ( .A(n814), .ZN(n815) );
  NAND2_X1 U909 ( .A1(n816), .A2(n815), .ZN(n819) );
  XNOR2_X1 U910 ( .A(G1986), .B(G290), .ZN(n960) );
  AND2_X1 U911 ( .A1(n960), .A2(n817), .ZN(n818) );
  NOR2_X1 U912 ( .A1(n819), .A2(n818), .ZN(n820) );
  OR2_X1 U913 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U914 ( .A(n824), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U915 ( .A(G2427), .B(G2451), .ZN(n834) );
  XOR2_X1 U916 ( .A(G2430), .B(G2443), .Z(n826) );
  XNOR2_X1 U917 ( .A(KEYINPUT107), .B(G2438), .ZN(n825) );
  XNOR2_X1 U918 ( .A(n826), .B(n825), .ZN(n830) );
  XOR2_X1 U919 ( .A(G2435), .B(G2454), .Z(n828) );
  XNOR2_X1 U920 ( .A(G1341), .B(G1348), .ZN(n827) );
  XNOR2_X1 U921 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U922 ( .A(n830), .B(n829), .Z(n832) );
  XNOR2_X1 U923 ( .A(KEYINPUT108), .B(G2446), .ZN(n831) );
  XNOR2_X1 U924 ( .A(n832), .B(n831), .ZN(n833) );
  XNOR2_X1 U925 ( .A(n834), .B(n833), .ZN(n835) );
  NAND2_X1 U926 ( .A1(n835), .A2(G14), .ZN(n916) );
  XNOR2_X1 U927 ( .A(KEYINPUT109), .B(n916), .ZN(G401) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n836), .ZN(G217) );
  INV_X1 U929 ( .A(n836), .ZN(G223) );
  NAND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n837) );
  XOR2_X1 U931 ( .A(KEYINPUT110), .B(n837), .Z(n838) );
  NAND2_X1 U932 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U934 ( .A1(n840), .A2(n839), .ZN(G188) );
  XNOR2_X1 U935 ( .A(G120), .B(KEYINPUT111), .ZN(G236) );
  NOR2_X1 U936 ( .A1(n842), .A2(n841), .ZN(G325) );
  XOR2_X1 U937 ( .A(KEYINPUT112), .B(G325), .Z(G261) );
  INV_X1 U939 ( .A(G132), .ZN(G219) );
  INV_X1 U940 ( .A(G96), .ZN(G221) );
  INV_X1 U941 ( .A(G82), .ZN(G220) );
  INV_X1 U942 ( .A(G69), .ZN(G235) );
  INV_X1 U943 ( .A(n843), .ZN(G319) );
  XNOR2_X1 U944 ( .A(KEYINPUT116), .B(n844), .ZN(n846) );
  XNOR2_X1 U945 ( .A(G1986), .B(G1981), .ZN(n845) );
  XNOR2_X1 U946 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U947 ( .A(n847), .B(KEYINPUT41), .Z(n850) );
  XOR2_X1 U948 ( .A(G1996), .B(n848), .Z(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U950 ( .A(G1956), .B(G1966), .Z(n852) );
  XNOR2_X1 U951 ( .A(G1976), .B(G1971), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U953 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U954 ( .A(G2474), .B(KEYINPUT115), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(G229) );
  XOR2_X1 U956 ( .A(G2678), .B(KEYINPUT113), .Z(n858) );
  XNOR2_X1 U957 ( .A(KEYINPUT114), .B(KEYINPUT43), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U959 ( .A(KEYINPUT42), .B(G2090), .Z(n860) );
  XNOR2_X1 U960 ( .A(G2067), .B(G2072), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U962 ( .A(n862), .B(n861), .Z(n865) );
  XOR2_X1 U963 ( .A(G2096), .B(n863), .Z(n864) );
  XNOR2_X1 U964 ( .A(n865), .B(n864), .ZN(n867) );
  XOR2_X1 U965 ( .A(G2078), .B(G2084), .Z(n866) );
  XNOR2_X1 U966 ( .A(n867), .B(n866), .ZN(G227) );
  NAND2_X1 U967 ( .A1(n890), .A2(G124), .ZN(n868) );
  XNOR2_X1 U968 ( .A(n868), .B(KEYINPUT44), .ZN(n870) );
  NAND2_X1 U969 ( .A1(G112), .A2(n891), .ZN(n869) );
  NAND2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n874) );
  NAND2_X1 U971 ( .A1(G136), .A2(n886), .ZN(n872) );
  NAND2_X1 U972 ( .A1(G100), .A2(n887), .ZN(n871) );
  NAND2_X1 U973 ( .A1(n872), .A2(n871), .ZN(n873) );
  NOR2_X1 U974 ( .A1(n874), .A2(n873), .ZN(G162) );
  XOR2_X1 U975 ( .A(KEYINPUT118), .B(KEYINPUT46), .Z(n885) );
  NAND2_X1 U976 ( .A1(G130), .A2(n890), .ZN(n876) );
  NAND2_X1 U977 ( .A1(G118), .A2(n891), .ZN(n875) );
  NAND2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n882) );
  NAND2_X1 U979 ( .A1(G142), .A2(n886), .ZN(n878) );
  NAND2_X1 U980 ( .A1(G106), .A2(n887), .ZN(n877) );
  NAND2_X1 U981 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U982 ( .A(KEYINPUT45), .B(n879), .ZN(n880) );
  XNOR2_X1 U983 ( .A(KEYINPUT117), .B(n880), .ZN(n881) );
  NOR2_X1 U984 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U985 ( .A(G160), .B(n883), .ZN(n884) );
  XNOR2_X1 U986 ( .A(n885), .B(n884), .ZN(n902) );
  NAND2_X1 U987 ( .A1(G139), .A2(n886), .ZN(n889) );
  NAND2_X1 U988 ( .A1(G103), .A2(n887), .ZN(n888) );
  NAND2_X1 U989 ( .A1(n889), .A2(n888), .ZN(n896) );
  NAND2_X1 U990 ( .A1(G127), .A2(n890), .ZN(n893) );
  NAND2_X1 U991 ( .A1(G115), .A2(n891), .ZN(n892) );
  NAND2_X1 U992 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U993 ( .A(KEYINPUT47), .B(n894), .Z(n895) );
  NOR2_X1 U994 ( .A1(n896), .A2(n895), .ZN(n934) );
  XOR2_X1 U995 ( .A(G162), .B(n934), .Z(n900) );
  XOR2_X1 U996 ( .A(n898), .B(n897), .Z(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n905) );
  XNOR2_X1 U999 ( .A(n903), .B(KEYINPUT48), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(n905), .B(n904), .ZN(n907) );
  XNOR2_X1 U1001 ( .A(n926), .B(G164), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n908), .ZN(G395) );
  INV_X1 U1004 ( .A(G171), .ZN(G301) );
  XOR2_X1 U1005 ( .A(KEYINPUT119), .B(n909), .Z(n911) );
  XOR2_X1 U1006 ( .A(G301), .B(G286), .Z(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n912), .B(n954), .ZN(n913) );
  XNOR2_X1 U1009 ( .A(n948), .B(n913), .ZN(n914) );
  NOR2_X1 U1010 ( .A1(n914), .A2(G37), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(n915), .B(KEYINPUT120), .ZN(G397) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n916), .ZN(n919) );
  NOR2_X1 U1013 ( .A1(G229), .A2(G227), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1015 ( .A1(n919), .A2(n918), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(G395), .A2(G397), .ZN(n920) );
  NAND2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(G57), .ZN(G237) );
  INV_X1 U1020 ( .A(n922), .ZN(n924) );
  NOR2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n933) );
  NOR2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1023 ( .A(KEYINPUT121), .B(n927), .Z(n928) );
  NAND2_X1 U1024 ( .A1(n929), .A2(n928), .ZN(n931) );
  XOR2_X1 U1025 ( .A(G160), .B(G2084), .Z(n930) );
  NOR2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n944) );
  XOR2_X1 U1028 ( .A(G2072), .B(n934), .Z(n936) );
  XOR2_X1 U1029 ( .A(G164), .B(G2078), .Z(n935) );
  NOR2_X1 U1030 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1031 ( .A(KEYINPUT50), .B(n937), .ZN(n942) );
  XOR2_X1 U1032 ( .A(G2090), .B(G162), .Z(n938) );
  NOR2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1034 ( .A(KEYINPUT51), .B(n940), .Z(n941) );
  NAND2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1036 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1037 ( .A(KEYINPUT52), .B(n945), .ZN(n946) );
  INV_X1 U1038 ( .A(KEYINPUT55), .ZN(n1014) );
  NAND2_X1 U1039 ( .A1(n946), .A2(n1014), .ZN(n947) );
  NAND2_X1 U1040 ( .A1(n947), .A2(G29), .ZN(n1023) );
  XOR2_X1 U1041 ( .A(KEYINPUT56), .B(G16), .Z(n971) );
  XOR2_X1 U1042 ( .A(n948), .B(G1341), .Z(n950) );
  XOR2_X1 U1043 ( .A(G299), .B(G1956), .Z(n949) );
  NAND2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n968) );
  XNOR2_X1 U1045 ( .A(G1966), .B(G168), .ZN(n952) );
  NAND2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(n953), .B(KEYINPUT57), .ZN(n966) );
  XNOR2_X1 U1048 ( .A(n954), .B(G1348), .ZN(n956) );
  XOR2_X1 U1049 ( .A(G301), .B(G1961), .Z(n955) );
  NAND2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n964) );
  NAND2_X1 U1051 ( .A1(G303), .A2(G1971), .ZN(n957) );
  NAND2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n962) );
  NAND2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n963) );
  NOR2_X1 U1055 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1056 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1057 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1058 ( .A(KEYINPUT124), .B(n969), .ZN(n970) );
  NOR2_X1 U1059 ( .A1(n971), .A2(n970), .ZN(n1020) );
  XNOR2_X1 U1060 ( .A(G1986), .B(G24), .ZN(n973) );
  XNOR2_X1 U1061 ( .A(G22), .B(G1971), .ZN(n972) );
  NOR2_X1 U1062 ( .A1(n973), .A2(n972), .ZN(n976) );
  XNOR2_X1 U1063 ( .A(G1976), .B(KEYINPUT125), .ZN(n974) );
  XNOR2_X1 U1064 ( .A(n974), .B(G23), .ZN(n975) );
  NAND2_X1 U1065 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1066 ( .A(KEYINPUT58), .B(n977), .Z(n991) );
  XOR2_X1 U1067 ( .A(G1966), .B(G21), .Z(n979) );
  XOR2_X1 U1068 ( .A(G1961), .B(G5), .Z(n978) );
  NAND2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n989) );
  XOR2_X1 U1070 ( .A(G1348), .B(KEYINPUT59), .Z(n980) );
  XNOR2_X1 U1071 ( .A(G4), .B(n980), .ZN(n982) );
  XNOR2_X1 U1072 ( .A(G20), .B(G1956), .ZN(n981) );
  NOR2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n986) );
  XNOR2_X1 U1074 ( .A(G1981), .B(G6), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(G1341), .B(G19), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1078 ( .A(KEYINPUT60), .B(n987), .ZN(n988) );
  NOR2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(n992), .B(KEYINPUT61), .ZN(n993) );
  XNOR2_X1 U1082 ( .A(n993), .B(KEYINPUT126), .ZN(n994) );
  NOR2_X1 U1083 ( .A1(G16), .A2(n994), .ZN(n1017) );
  XNOR2_X1 U1084 ( .A(G27), .B(n995), .ZN(n1006) );
  XNOR2_X1 U1085 ( .A(KEYINPUT123), .B(G2067), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(n996), .B(G26), .ZN(n1001) );
  XOR2_X1 U1087 ( .A(G32), .B(G1996), .Z(n997) );
  NAND2_X1 U1088 ( .A1(n997), .A2(G28), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(G33), .B(G2072), .ZN(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(G25), .B(G1991), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(KEYINPUT122), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(n1007), .B(KEYINPUT53), .ZN(n1010) );
  XOR2_X1 U1097 ( .A(G2084), .B(G34), .Z(n1008) );
  XNOR2_X1 U1098 ( .A(KEYINPUT54), .B(n1008), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(G35), .B(G2090), .ZN(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(n1014), .B(n1013), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(G29), .A2(n1015), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(G11), .A2(n1018), .ZN(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1107 ( .A(KEYINPUT127), .B(n1021), .Z(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1024), .ZN(G150) );
  INV_X1 U1110 ( .A(G150), .ZN(G311) );
  INV_X1 U1111 ( .A(G303), .ZN(G166) );
endmodule

