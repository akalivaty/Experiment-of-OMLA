//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 1 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  AND2_X1   g002(.A1(KEYINPUT64), .A2(G143), .ZN(new_n189));
  NOR2_X1   g003(.A1(KEYINPUT64), .A2(G143), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT65), .A2(G146), .ZN(new_n192));
  NOR2_X1   g006(.A1(KEYINPUT65), .A2(G146), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n191), .B1(new_n194), .B2(G143), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT1), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n196), .B1(new_n194), .B2(G143), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n195), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT65), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(new_n188), .ZN(new_n201));
  NAND2_X1  g015(.A1(KEYINPUT65), .A2(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(G143), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n201), .A2(KEYINPUT66), .A3(G143), .A4(new_n202), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT64), .A2(G143), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(G146), .A3(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n205), .A2(new_n206), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n199), .A2(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(G125), .ZN(new_n215));
  INV_X1    g029(.A(G125), .ZN(new_n216));
  AND2_X1   g030(.A1(KEYINPUT0), .A2(G128), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n205), .A2(new_n206), .A3(new_n211), .A4(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(KEYINPUT0), .A2(G128), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n195), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n216), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n215), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G224), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(G953), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n223), .B(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(G110), .B(G122), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(KEYINPUT90), .ZN(new_n228));
  INV_X1    g042(.A(G104), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(KEYINPUT3), .ZN(new_n230));
  INV_X1    g044(.A(G107), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT80), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT80), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G107), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n230), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT81), .B(G101), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT3), .B1(new_n229), .B2(G107), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n229), .A2(G107), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n235), .A2(new_n236), .A3(new_n237), .A4(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT82), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G101), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT81), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT81), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G101), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n243), .A2(new_n245), .A3(new_n238), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n246), .A2(KEYINPUT82), .A3(new_n237), .A4(new_n235), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n241), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n249), .B1(new_n250), .B2(G101), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n250), .A2(new_n249), .A3(G101), .ZN(new_n253));
  XOR2_X1   g067(.A(KEYINPUT2), .B(G113), .Z(new_n254));
  XNOR2_X1  g068(.A(G116), .B(G119), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G119), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G116), .ZN(new_n258));
  INV_X1    g072(.A(G116), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G119), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT2), .B(G113), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n256), .A2(KEYINPUT68), .A3(new_n263), .ZN(new_n264));
  OR3_X1    g078(.A1(new_n254), .A2(KEYINPUT68), .A3(new_n255), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n253), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n252), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n232), .A2(new_n234), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n229), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n231), .A2(KEYINPUT83), .A3(G104), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT83), .B1(new_n231), .B2(G104), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n242), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n273), .B1(new_n241), .B2(new_n247), .ZN(new_n274));
  OR2_X1    g088(.A1(new_n258), .A2(KEYINPUT5), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n275), .A2(G113), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n255), .A2(KEYINPUT5), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n276), .A2(new_n277), .B1(new_n255), .B2(new_n254), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n267), .A2(KEYINPUT89), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT89), .B1(new_n267), .B2(new_n279), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n228), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n283));
  INV_X1    g097(.A(new_n279), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n253), .A2(new_n264), .A3(new_n265), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n285), .B1(new_n248), .B2(new_n251), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n282), .A2(new_n283), .B1(new_n287), .B2(new_n227), .ZN(new_n288));
  INV_X1    g102(.A(new_n228), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT89), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n290), .B1(new_n284), .B2(new_n286), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n267), .A2(KEYINPUT89), .A3(new_n279), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n289), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT6), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n226), .B1(new_n288), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(G210), .B1(G237), .B2(G902), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n273), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n248), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n278), .ZN(new_n300));
  XOR2_X1   g114(.A(KEYINPUT91), .B(KEYINPUT8), .Z(new_n301));
  XNOR2_X1  g115(.A(new_n301), .B(new_n227), .ZN(new_n302));
  OR2_X1    g116(.A1(new_n276), .A2(KEYINPUT92), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n276), .A2(KEYINPUT92), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n277), .A3(new_n304), .ZN(new_n305));
  AND2_X1   g119(.A1(new_n305), .A2(new_n256), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n300), .B(new_n302), .C1(new_n306), .C2(new_n299), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n287), .A2(new_n227), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT7), .B1(new_n224), .B2(G953), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n309), .B1(new_n215), .B2(new_n222), .ZN(new_n310));
  OR3_X1    g124(.A1(new_n215), .A2(new_n222), .A3(new_n309), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n307), .A2(new_n308), .A3(new_n310), .A4(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G902), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR3_X1   g128(.A1(new_n295), .A2(new_n297), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n226), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n308), .B1(new_n293), .B2(KEYINPUT6), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n282), .A2(new_n283), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n314), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n296), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n187), .B1(new_n315), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT97), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT20), .ZN(new_n324));
  XNOR2_X1  g138(.A(G113), .B(G122), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n325), .B(new_n229), .ZN(new_n326));
  NOR3_X1   g140(.A1(new_n216), .A2(KEYINPUT16), .A3(G140), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n327), .A2(KEYINPUT74), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(G125), .B(G140), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n327), .B1(new_n330), .B2(KEYINPUT16), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT74), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n329), .B(G146), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G237), .ZN(new_n334));
  INV_X1    g148(.A(G953), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n334), .A2(new_n335), .A3(G143), .A4(G214), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n209), .A2(new_n210), .ZN(new_n337));
  INV_X1    g151(.A(G214), .ZN(new_n338));
  NOR3_X1   g152(.A1(new_n338), .A2(G237), .A3(G953), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n336), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G131), .ZN(new_n341));
  INV_X1    g155(.A(G131), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n342), .B(new_n336), .C1(new_n337), .C2(new_n339), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n330), .B(KEYINPUT77), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT19), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT94), .ZN(new_n348));
  INV_X1    g162(.A(new_n330), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT19), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT94), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n345), .A2(new_n351), .A3(new_n346), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n348), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n194), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n333), .B(new_n344), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(KEYINPUT18), .A2(G131), .ZN(new_n356));
  OR3_X1    g170(.A1(new_n340), .A2(KEYINPUT93), .A3(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n356), .B1(new_n340), .B2(KEYINPUT93), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n345), .A2(new_n194), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n349), .A2(G146), .ZN(new_n360));
  AOI22_X1  g174(.A1(new_n357), .A2(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n326), .B1(new_n355), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT17), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n341), .A2(new_n364), .A3(new_n343), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT95), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT95), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n341), .A2(new_n367), .A3(new_n364), .A4(new_n343), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G140), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G125), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n216), .A2(G140), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n372), .A3(KEYINPUT16), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT16), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(new_n370), .A3(G125), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n332), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n188), .B1(new_n376), .B2(new_n328), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT75), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n333), .A3(new_n378), .ZN(new_n379));
  OAI211_X1 g193(.A(KEYINPUT75), .B(new_n188), .C1(new_n376), .C2(new_n328), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n341), .A2(new_n364), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n369), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(new_n362), .A3(new_n326), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT96), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n382), .B1(new_n366), .B2(new_n368), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n361), .B1(new_n388), .B2(new_n381), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(KEYINPUT96), .A3(new_n326), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n363), .B1(new_n387), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(G475), .A2(G902), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n323), .B(new_n324), .C1(new_n391), .C2(new_n393), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n389), .A2(new_n326), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n395), .B1(new_n387), .B2(new_n390), .ZN(new_n396));
  OAI21_X1  g210(.A(G475), .B1(new_n396), .B2(G902), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n323), .B1(new_n391), .B2(new_n393), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n355), .A2(new_n362), .ZN(new_n400));
  INV_X1    g214(.A(new_n326), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AND4_X1   g216(.A1(KEYINPUT96), .A2(new_n384), .A3(new_n326), .A4(new_n362), .ZN(new_n403));
  AOI21_X1  g217(.A(KEYINPUT96), .B1(new_n389), .B2(new_n326), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(KEYINPUT97), .A3(new_n392), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n399), .A2(new_n406), .A3(KEYINPUT20), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n398), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n209), .A2(G128), .A3(new_n210), .ZN(new_n409));
  INV_X1    g223(.A(G134), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n198), .A2(G143), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n259), .A2(G122), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(KEYINPUT98), .ZN(new_n414));
  INV_X1    g228(.A(G122), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G116), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n268), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n414), .A2(new_n418), .A3(new_n416), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT13), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n411), .B1(new_n409), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n409), .ZN(new_n423));
  OR3_X1    g237(.A1(new_n423), .A2(KEYINPUT99), .A3(KEYINPUT13), .ZN(new_n424));
  OAI21_X1  g238(.A(KEYINPUT99), .B1(new_n423), .B2(KEYINPUT13), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n422), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI221_X1 g240(.A(new_n412), .B1(new_n419), .B2(new_n420), .C1(new_n426), .C2(new_n410), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n414), .A2(KEYINPUT14), .B1(G116), .B2(new_n415), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n428), .B1(KEYINPUT14), .B2(new_n414), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(G107), .ZN(new_n430));
  INV_X1    g244(.A(new_n420), .ZN(new_n431));
  INV_X1    g245(.A(new_n412), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n410), .B1(new_n409), .B2(new_n411), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n430), .B(new_n431), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n427), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT9), .B(G234), .ZN(new_n436));
  INV_X1    g250(.A(G217), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n436), .A2(new_n437), .A3(G953), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n427), .A2(new_n434), .A3(new_n438), .ZN(new_n441));
  AOI21_X1  g255(.A(G902), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G478), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(KEYINPUT15), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n442), .B(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n335), .A2(G952), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n448), .B1(G234), .B2(G237), .ZN(new_n449));
  AOI211_X1 g263(.A(new_n313), .B(new_n335), .C1(G234), .C2(G237), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(G898), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n447), .A2(new_n453), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n322), .A2(new_n408), .A3(new_n454), .ZN(new_n455));
  XOR2_X1   g269(.A(KEYINPUT26), .B(G101), .Z(new_n456));
  NAND3_X1  g270(.A1(new_n334), .A2(new_n335), .A3(G210), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n456), .B(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n458), .B(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT28), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n264), .A2(new_n265), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G137), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G134), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n410), .A2(G137), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n342), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n464), .A2(KEYINPUT11), .A3(G134), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n468), .A2(new_n466), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT67), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT11), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n471), .B1(new_n410), .B2(G137), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n469), .A2(new_n470), .A3(new_n342), .A4(new_n472), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n472), .A2(new_n468), .A3(new_n342), .A4(new_n466), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT67), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n467), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n214), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n472), .A2(new_n468), .A3(new_n466), .ZN(new_n478));
  AOI22_X1  g292(.A1(new_n473), .A2(new_n475), .B1(G131), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n218), .A2(new_n221), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n463), .B1(new_n477), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n478), .A2(G131), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n474), .A2(KEYINPUT67), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n474), .A2(KEYINPUT67), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n218), .A3(new_n221), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n214), .A2(new_n476), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n488), .A3(new_n462), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n461), .B1(new_n482), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n461), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n460), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT30), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n487), .A2(new_n494), .A3(new_n488), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n494), .B1(new_n487), .B2(new_n488), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n463), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n460), .ZN(new_n498));
  XOR2_X1   g312(.A(KEYINPUT71), .B(KEYINPUT31), .Z(new_n499));
  NAND4_X1  g313(.A1(new_n497), .A2(new_n489), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n493), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n497), .A2(new_n489), .A3(new_n498), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n502), .A2(KEYINPUT70), .A3(KEYINPUT31), .ZN(new_n503));
  AOI21_X1  g317(.A(KEYINPUT70), .B1(new_n502), .B2(KEYINPUT31), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(G472), .A2(G902), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(KEYINPUT32), .A3(new_n506), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n487), .A2(new_n488), .A3(new_n462), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n462), .B1(new_n487), .B2(new_n488), .ZN(new_n509));
  OAI21_X1  g323(.A(KEYINPUT28), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n510), .A2(KEYINPUT29), .A3(new_n491), .A4(new_n498), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n313), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT73), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT73), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n511), .A2(new_n514), .A3(new_n313), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n510), .A2(new_n491), .A3(new_n498), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT29), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT30), .B1(new_n477), .B2(new_n481), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n487), .A2(new_n488), .A3(new_n494), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n508), .B1(new_n520), .B2(new_n463), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n516), .B(new_n517), .C1(new_n521), .C2(new_n498), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n513), .A2(new_n515), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G472), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n507), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT32), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n493), .A2(new_n500), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n502), .A2(KEYINPUT31), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT70), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n502), .A2(KEYINPUT70), .A3(KEYINPUT31), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n527), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n506), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n526), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT72), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT32), .B1(new_n505), .B2(new_n506), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT72), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n525), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n437), .B1(G234), .B2(new_n313), .ZN(new_n540));
  XOR2_X1   g354(.A(KEYINPUT24), .B(G110), .Z(new_n541));
  XNOR2_X1  g355(.A(G119), .B(G128), .ZN(new_n542));
  OR3_X1    g356(.A1(new_n541), .A2(KEYINPUT76), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT76), .B1(new_n541), .B2(new_n542), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT23), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n257), .B2(G128), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n198), .A2(KEYINPUT23), .A3(G119), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n546), .B(new_n547), .C1(G119), .C2(new_n198), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n543), .B(new_n544), .C1(G110), .C2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n549), .A2(new_n333), .A3(new_n359), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT78), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT78), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n549), .A2(new_n552), .A3(new_n333), .A4(new_n359), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n541), .A2(new_n542), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n548), .A2(G110), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n379), .A2(new_n380), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT22), .B(G137), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n335), .A2(G221), .A3(G234), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n554), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n560), .B1(new_n554), .B2(new_n557), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n563), .A2(KEYINPUT25), .A3(new_n313), .ZN(new_n564));
  AOI21_X1  g378(.A(KEYINPUT25), .B1(new_n563), .B2(new_n313), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n540), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n540), .A2(G902), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(G221), .B1(new_n436), .B2(G902), .ZN(new_n571));
  XOR2_X1   g385(.A(new_n571), .B(KEYINPUT79), .Z(new_n572));
  NAND2_X1  g386(.A1(new_n206), .A2(new_n211), .ZN(new_n573));
  AOI21_X1  g387(.A(KEYINPUT66), .B1(new_n194), .B2(G143), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n196), .B1(new_n337), .B2(new_n188), .ZN(new_n575));
  OAI22_X1  g389(.A1(new_n573), .A2(new_n574), .B1(new_n575), .B2(new_n198), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n213), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n274), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT10), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n252), .A2(new_n218), .A3(new_n221), .A4(new_n253), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n579), .B1(new_n199), .B2(new_n213), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n274), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n580), .A2(new_n581), .A3(new_n479), .A4(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT12), .B1(new_n486), .B2(KEYINPUT84), .ZN(new_n585));
  INV_X1    g399(.A(new_n214), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n299), .A2(new_n586), .ZN(new_n587));
  AOI211_X1 g401(.A(new_n479), .B(new_n585), .C1(new_n587), .C2(new_n578), .ZN(new_n588));
  INV_X1    g402(.A(new_n585), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n578), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n589), .B1(new_n590), .B2(new_n486), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n584), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(G110), .B(G140), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n335), .A2(G227), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n595), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n584), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT85), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n599), .A2(new_n600), .A3(new_n486), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n600), .B1(new_n599), .B2(new_n486), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n598), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT86), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n596), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n604), .B1(new_n596), .B2(new_n603), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n313), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(G469), .ZN(new_n608));
  INV_X1    g422(.A(new_n584), .ZN(new_n609));
  AOI21_X1  g423(.A(KEYINPUT10), .B1(new_n577), .B2(new_n274), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n582), .A2(new_n274), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n253), .A2(new_n218), .A3(new_n221), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(new_n248), .B2(new_n251), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(KEYINPUT85), .B1(new_n614), .B2(new_n479), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n599), .A2(new_n600), .A3(new_n486), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n609), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(KEYINPUT88), .B1(new_n617), .B2(new_n597), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n584), .B1(new_n601), .B2(new_n602), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT88), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n619), .A2(new_n620), .A3(new_n595), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n598), .B1(new_n588), .B2(new_n591), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n618), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT87), .B(G469), .Z(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n313), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n572), .B1(new_n608), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n455), .A2(new_n539), .A3(new_n570), .A4(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(new_n627), .B(KEYINPUT100), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(new_n236), .ZN(G3));
  NOR2_X1   g443(.A1(new_n532), .A2(G902), .ZN(new_n630));
  INV_X1    g444(.A(G472), .ZN(new_n631));
  OAI22_X1  g445(.A1(new_n630), .A2(new_n631), .B1(new_n533), .B2(new_n532), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n569), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n453), .B(new_n187), .C1(new_n315), .C2(new_n321), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n440), .A2(new_n441), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(KEYINPUT33), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n440), .A2(new_n637), .A3(new_n441), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n636), .A2(G478), .A3(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n443), .A2(new_n313), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n640), .B1(new_n442), .B2(new_n443), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n399), .A2(new_n406), .A3(KEYINPUT20), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n394), .A2(new_n397), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n634), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n633), .A2(new_n626), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT34), .B(G104), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G6));
  NAND3_X1  g464(.A1(new_n398), .A2(new_n407), .A3(new_n446), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n634), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n633), .A2(new_n626), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT35), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  INV_X1    g469(.A(new_n632), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n554), .A2(new_n557), .ZN(new_n657));
  INV_X1    g471(.A(new_n560), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(KEYINPUT36), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n657), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n567), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n566), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n455), .A2(new_n626), .A3(new_n656), .A4(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT37), .B(G110), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G12));
  AND3_X1   g479(.A1(new_n539), .A2(new_n626), .A3(new_n662), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n449), .B(KEYINPUT102), .ZN(new_n667));
  INV_X1    g481(.A(G900), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(KEYINPUT101), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n668), .A2(KEYINPUT101), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n450), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n398), .A2(new_n407), .A3(new_n446), .A4(new_n672), .ZN(new_n673));
  OAI21_X1  g487(.A(KEYINPUT103), .B1(new_n673), .B2(new_n322), .ZN(new_n674));
  AND4_X1   g488(.A1(new_n407), .A2(new_n394), .A3(new_n446), .A4(new_n397), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n676));
  INV_X1    g490(.A(new_n187), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n297), .B1(new_n295), .B2(new_n314), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n319), .A2(new_n296), .A3(new_n320), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n675), .A2(new_n676), .A3(new_n680), .A4(new_n672), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n674), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n666), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G128), .ZN(G30));
  NAND2_X1  g498(.A1(new_n678), .A2(new_n679), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n662), .A2(new_n447), .A3(new_n677), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n687), .A2(new_n408), .A3(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n521), .A2(new_n460), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n482), .A2(new_n489), .A3(new_n460), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n313), .ZN(new_n692));
  OAI21_X1  g506(.A(G472), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n507), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n536), .A3(new_n538), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n672), .B(KEYINPUT39), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n626), .A2(new_n696), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n689), .B(new_n695), .C1(KEYINPUT40), .C2(new_n697), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n697), .A2(KEYINPUT40), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n337), .B(KEYINPUT105), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G45));
  OAI211_X1 g516(.A(new_n643), .B(new_n672), .C1(new_n644), .C2(new_n645), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n322), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n539), .A2(new_n704), .A3(new_n626), .A4(new_n662), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  AND3_X1   g520(.A1(new_n623), .A2(new_n313), .A3(new_n624), .ZN(new_n707));
  INV_X1    g521(.A(G469), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n623), .B2(new_n313), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n707), .A2(new_n709), .A3(new_n572), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n710), .A2(new_n539), .A3(new_n647), .A4(new_n570), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT41), .B(G113), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT106), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n711), .B(new_n713), .ZN(G15));
  NAND4_X1  g528(.A1(new_n710), .A2(new_n539), .A3(new_n570), .A4(new_n652), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G116), .ZN(G18));
  NOR2_X1   g530(.A1(new_n408), .A2(new_n454), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n539), .A2(new_n717), .A3(new_n662), .ZN(new_n718));
  INV_X1    g532(.A(new_n709), .ZN(new_n719));
  INV_X1    g533(.A(new_n572), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n719), .A2(new_n720), .A3(new_n625), .A4(new_n680), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(new_n257), .ZN(G21));
  NOR2_X1   g537(.A1(new_n644), .A2(new_n645), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n634), .A2(new_n724), .A3(new_n447), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT107), .B(G472), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n727), .B1(new_n505), .B2(new_n313), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n533), .B1(new_n501), .B2(new_n528), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n569), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n725), .A2(new_n710), .A3(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  NOR2_X1   g546(.A1(new_n728), .A2(new_n729), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n642), .B1(new_n398), .B2(new_n407), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n733), .A2(new_n734), .A3(new_n662), .A4(new_n672), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n721), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(new_n216), .ZN(G27));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n507), .B(new_n524), .C1(new_n537), .C2(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n534), .A2(KEYINPUT108), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n570), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n596), .A2(new_n603), .ZN(new_n742));
  OAI21_X1  g556(.A(G469), .B1(new_n742), .B2(G902), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n625), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n572), .A2(new_n677), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n678), .A2(new_n679), .A3(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n744), .A2(new_n734), .A3(new_n672), .A4(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT42), .B1(new_n741), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n703), .A2(KEYINPUT42), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n678), .A2(new_n679), .A3(new_n745), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n750), .B1(new_n625), .B2(new_n743), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n539), .A2(new_n749), .A3(new_n570), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n342), .ZN(G33));
  XNOR2_X1  g568(.A(new_n537), .B(new_n535), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n569), .B1(new_n755), .B2(new_n525), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT109), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n673), .B(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n756), .A2(new_n757), .A3(new_n751), .A4(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n539), .A2(new_n570), .A3(new_n751), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n673), .B(KEYINPUT109), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT110), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G134), .ZN(G36));
  NAND2_X1  g579(.A1(new_n632), .A2(new_n662), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT112), .ZN(new_n767));
  OR3_X1    g581(.A1(new_n644), .A2(KEYINPUT111), .A3(new_n645), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n408), .A2(KEYINPUT111), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n768), .A2(new_n769), .A3(KEYINPUT43), .A4(new_n643), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT43), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n408), .B2(new_n642), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n767), .A2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n767), .A2(KEYINPUT44), .A3(new_n773), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n678), .A2(new_n187), .A3(new_n679), .ZN(new_n778));
  XOR2_X1   g592(.A(new_n778), .B(KEYINPUT113), .Z(new_n779));
  NOR2_X1   g593(.A1(new_n708), .A2(new_n313), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT45), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n781), .B1(new_n605), .B2(new_n606), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n708), .B1(new_n742), .B2(KEYINPUT45), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n784), .A2(KEYINPUT46), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n625), .B1(new_n784), .B2(KEYINPUT46), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n720), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n696), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n776), .A2(new_n777), .A3(new_n779), .A4(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G137), .ZN(G39));
  NAND2_X1  g605(.A1(new_n787), .A2(KEYINPUT114), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n793), .B(new_n720), .C1(new_n785), .C2(new_n786), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n795), .A2(KEYINPUT47), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n792), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n795), .A3(KEYINPUT47), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n795), .A2(KEYINPUT47), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n792), .A2(new_n799), .A3(new_n794), .A4(new_n796), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  OR3_X1    g615(.A1(new_n703), .A2(new_n570), .A3(new_n778), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n539), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G140), .ZN(G42));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n736), .B1(new_n666), .B2(new_n682), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n566), .A2(new_n720), .A3(new_n661), .A4(new_n672), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n808), .B1(new_n625), .B2(new_n743), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n680), .A2(new_n408), .A3(new_n446), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n695), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n705), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT52), .B1(new_n807), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n539), .A2(new_n626), .A3(new_n662), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n674), .A2(new_n681), .ZN(new_n815));
  OAI22_X1  g629(.A1(new_n814), .A2(new_n815), .B1(new_n721), .B2(new_n735), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n705), .A2(new_n811), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n813), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n711), .A2(new_n715), .A3(new_n731), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n722), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n447), .A2(new_n672), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n408), .A2(new_n778), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n824), .A2(new_n539), .A3(new_n626), .A4(new_n662), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n733), .A2(new_n662), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n826), .A2(new_n734), .A3(new_n672), .A4(new_n751), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n748), .A2(new_n752), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n627), .A2(new_n663), .A3(new_n648), .A4(new_n653), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n822), .A2(new_n828), .A3(new_n764), .A4(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n806), .B1(new_n820), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n822), .A2(new_n764), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n807), .A2(new_n812), .A3(KEYINPUT52), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n818), .B1(new_n816), .B2(new_n817), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n827), .A2(new_n825), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n829), .A2(new_n753), .A3(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n834), .A2(new_n837), .A3(KEYINPUT53), .A4(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n832), .A2(new_n833), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n832), .A2(new_n840), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT54), .ZN(new_n843));
  INV_X1    g657(.A(new_n667), .ZN(new_n844));
  AOI21_X1  g658(.A(KEYINPUT116), .B1(new_n773), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n846));
  AOI211_X1 g660(.A(new_n846), .B(new_n667), .C1(new_n770), .C2(new_n772), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n741), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n719), .A2(new_n720), .A3(new_n625), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n850), .A2(new_n778), .ZN(new_n851));
  XOR2_X1   g665(.A(KEYINPUT121), .B(KEYINPUT48), .Z(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n848), .A2(new_n849), .A3(new_n851), .A4(new_n853), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n849), .B(new_n851), .C1(new_n845), .C2(new_n847), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n852), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n721), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n858), .B(new_n730), .C1(new_n845), .C2(new_n847), .ZN(new_n859));
  INV_X1    g673(.A(new_n695), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n570), .A2(new_n449), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n851), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n448), .B1(new_n862), .B2(new_n734), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT120), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n859), .A2(new_n866), .A3(new_n863), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n857), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n868), .A2(KEYINPUT122), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n868), .A2(KEYINPUT122), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n841), .B(new_n843), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT51), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n408), .A2(new_n643), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n862), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT119), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n862), .A2(new_n876), .A3(new_n873), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n848), .A2(new_n826), .A3(new_n851), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n687), .A2(new_n850), .A3(new_n187), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n730), .B(new_n881), .C1(new_n845), .C2(new_n847), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n884), .A2(KEYINPUT50), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(KEYINPUT50), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n880), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n848), .A2(new_n730), .A3(new_n779), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n719), .A2(new_n572), .A3(new_n625), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT117), .Z(new_n891));
  NAND3_X1  g705(.A1(new_n798), .A2(new_n891), .A3(new_n800), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n872), .B1(new_n887), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n798), .A2(new_n800), .A3(new_n890), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n872), .B1(new_n889), .B2(new_n895), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n896), .B(new_n880), .C1(new_n885), .C2(new_n886), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  OAI22_X1  g712(.A1(new_n871), .A2(new_n898), .B1(G952), .B2(G953), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n719), .A2(new_n625), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT49), .ZN(new_n901));
  INV_X1    g715(.A(new_n687), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n902), .A2(new_n570), .A3(new_n643), .A4(new_n745), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n768), .A2(new_n769), .ZN(new_n904));
  OR4_X1    g718(.A1(new_n695), .A2(new_n901), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n899), .A2(new_n905), .ZN(G75));
  NAND3_X1  g720(.A1(new_n842), .A2(G210), .A3(G902), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT56), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n317), .A2(new_n318), .A3(new_n316), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(new_n295), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT55), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n907), .A2(new_n908), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n911), .B1(new_n907), .B2(new_n908), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n335), .A2(G952), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(G51));
  INV_X1    g729(.A(KEYINPUT123), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n841), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n832), .A2(new_n840), .A3(KEYINPUT123), .A4(new_n833), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n917), .A2(new_n843), .A3(new_n918), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n780), .B(KEYINPUT57), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n623), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n832), .A2(new_n840), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n923), .A2(new_n313), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n924), .A2(new_n782), .A3(new_n783), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n914), .B1(new_n922), .B2(new_n925), .ZN(G54));
  NAND3_X1  g740(.A1(new_n924), .A2(KEYINPUT58), .A3(G475), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n391), .ZN(new_n928));
  INV_X1    g742(.A(new_n914), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n924), .A2(KEYINPUT58), .A3(G475), .A4(new_n405), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(G60));
  XOR2_X1   g745(.A(KEYINPUT124), .B(KEYINPUT59), .Z(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(new_n640), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n843), .B2(new_n841), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n636), .A2(new_n638), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n929), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n933), .B1(new_n636), .B2(new_n638), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n936), .B1(new_n919), .B2(new_n937), .ZN(G63));
  INV_X1    g752(.A(new_n562), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n554), .A2(new_n557), .A3(new_n560), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(G217), .A2(G902), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n942), .A2(KEYINPUT60), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(KEYINPUT60), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n941), .B1(new_n923), .B2(new_n945), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n842), .A2(new_n660), .A3(new_n943), .A4(new_n944), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n946), .A2(new_n929), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT61), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(G66));
  OAI21_X1  g764(.A(G953), .B1(new_n451), .B2(new_n224), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n822), .A2(new_n830), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n951), .B1(new_n953), .B2(G953), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n288), .B(new_n294), .C1(G898), .C2(new_n335), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(G69));
  XOR2_X1   g770(.A(new_n520), .B(new_n353), .Z(new_n957));
  NAND2_X1  g771(.A1(new_n807), .A2(new_n705), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n959), .B(KEYINPUT62), .C1(new_n699), .C2(new_n698), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT62), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(new_n700), .B2(new_n958), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n778), .B1(new_n646), .B2(new_n651), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n756), .A2(new_n626), .A3(new_n696), .A4(new_n964), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT125), .Z(new_n966));
  AND2_X1   g780(.A1(new_n966), .A2(new_n790), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n963), .A2(new_n967), .A3(new_n804), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n957), .B1(new_n968), .B2(new_n335), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  AOI211_X1 g784(.A(new_n539), .B(new_n802), .C1(new_n798), .C2(new_n800), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n849), .A2(new_n810), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n753), .B1(new_n789), .B2(new_n972), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n790), .A2(new_n764), .A3(new_n959), .A4(new_n973), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n335), .ZN(new_n976));
  INV_X1    g790(.A(new_n957), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(G900), .B2(G953), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n335), .B1(G227), .B2(G900), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n970), .A2(new_n979), .A3(KEYINPUT126), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(KEYINPUT126), .ZN(new_n982));
  OR2_X1    g796(.A1(new_n980), .A2(KEYINPUT126), .ZN(new_n983));
  INV_X1    g797(.A(new_n978), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n984), .B1(new_n975), .B2(new_n335), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n982), .B(new_n983), .C1(new_n985), .C2(new_n969), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n981), .A2(new_n986), .ZN(G72));
  NAND4_X1  g801(.A1(new_n963), .A2(new_n967), .A3(new_n804), .A4(new_n953), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT127), .ZN(new_n989));
  NAND2_X1  g803(.A1(G472), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT63), .Z(new_n991));
  NAND3_X1  g805(.A1(new_n988), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n690), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n989), .B1(new_n988), .B2(new_n991), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NOR3_X1   g809(.A1(new_n971), .A2(new_n974), .A3(new_n952), .ZN(new_n996));
  INV_X1    g810(.A(new_n991), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n460), .B(new_n521), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n521), .B(new_n498), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n842), .A2(new_n991), .A3(new_n999), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n998), .A2(new_n1000), .A3(new_n929), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n995), .A2(new_n1001), .ZN(G57));
endmodule


