//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 1 1 0 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G146), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT65), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT64), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT64), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n190), .B1(new_n195), .B2(G143), .ZN(new_n196));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G128), .Z(new_n197));
  NAND4_X1  g011(.A1(new_n192), .A2(new_n194), .A3(new_n189), .A4(new_n187), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n195), .A2(G143), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n191), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n200), .A2(KEYINPUT0), .A3(G128), .A4(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n199), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G125), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT68), .B(G128), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n187), .B1(new_n192), .B2(new_n194), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(new_n196), .A3(new_n198), .ZN(new_n210));
  INV_X1    g024(.A(G125), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n200), .A2(new_n208), .A3(G128), .A4(new_n202), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n205), .A2(new_n213), .ZN(new_n214));
  XOR2_X1   g028(.A(KEYINPUT90), .B(G224), .Z(new_n215));
  INV_X1    g029(.A(G953), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT91), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n217), .B(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n214), .B(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G107), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(KEYINPUT85), .A3(G104), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT3), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n221), .A2(G104), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n226), .A2(new_n221), .A3(KEYINPUT85), .A4(G104), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n223), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G101), .ZN(new_n229));
  INV_X1    g043(.A(G101), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n223), .A2(new_n225), .A3(new_n230), .A4(new_n227), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n229), .A2(KEYINPUT4), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G119), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G116), .ZN(new_n234));
  INV_X1    g048(.A(G116), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G119), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT2), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(G113), .ZN(new_n238));
  INV_X1    g052(.A(G113), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(KEYINPUT2), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n234), .B(new_n236), .C1(new_n238), .C2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n234), .A2(new_n236), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT2), .B(G113), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n241), .A2(new_n244), .A3(KEYINPUT69), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n241), .A2(new_n244), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n228), .A2(new_n249), .A3(G101), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n232), .A2(new_n245), .A3(new_n248), .A4(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n234), .A2(new_n236), .A3(KEYINPUT5), .ZN(new_n252));
  OR3_X1    g066(.A1(new_n235), .A2(KEYINPUT5), .A3(G119), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(G113), .ZN(new_n254));
  INV_X1    g068(.A(G104), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(G107), .ZN(new_n256));
  OAI21_X1  g070(.A(G101), .B1(new_n224), .B2(new_n256), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n231), .A2(new_n254), .A3(new_n241), .A4(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT88), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n231), .A2(new_n257), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n254), .A2(new_n241), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(new_n263), .A3(KEYINPUT88), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n251), .A2(new_n260), .A3(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(G110), .B(G122), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n258), .B(KEYINPUT88), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(new_n266), .A3(new_n251), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(KEYINPUT6), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT89), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n266), .B1(new_n269), .B2(new_n251), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AND4_X1   g089(.A1(new_n272), .A2(new_n265), .A3(new_n274), .A4(new_n267), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n220), .B(new_n271), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  XOR2_X1   g091(.A(KEYINPUT92), .B(KEYINPUT7), .Z(new_n278));
  OAI21_X1  g092(.A(new_n214), .B1(new_n219), .B2(new_n278), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n279), .A2(new_n270), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT7), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n217), .B(KEYINPUT91), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT93), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n219), .A2(KEYINPUT93), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n284), .A2(new_n205), .A3(new_n213), .A4(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n266), .B(KEYINPUT8), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n262), .A2(new_n263), .ZN(new_n288));
  INV_X1    g102(.A(new_n258), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(G902), .B1(new_n280), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n277), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(G210), .B1(G237), .B2(G902), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT94), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n277), .A2(new_n294), .A3(new_n292), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G214), .B1(G237), .B2(G902), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n293), .A2(KEYINPUT94), .A3(new_n295), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT95), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT95), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n299), .A2(new_n304), .A3(new_n300), .A4(new_n301), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G469), .ZN(new_n307));
  INV_X1    g121(.A(G902), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n232), .A2(new_n250), .ZN(new_n309));
  INV_X1    g123(.A(new_n204), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n261), .B1(new_n210), .B2(new_n212), .ZN(new_n311));
  AOI22_X1  g125(.A1(new_n309), .A2(new_n310), .B1(new_n311), .B2(KEYINPUT10), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT86), .ZN(new_n313));
  INV_X1    g127(.A(G134), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT11), .B1(new_n314), .B2(G137), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT11), .ZN(new_n316));
  INV_X1    g130(.A(G137), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n317), .A3(G134), .ZN(new_n318));
  AOI22_X1  g132(.A1(new_n315), .A2(new_n318), .B1(new_n314), .B2(G137), .ZN(new_n319));
  INV_X1    g133(.A(G131), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n319), .B(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(G128), .B1(new_n188), .B2(new_n208), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n323), .B1(new_n207), .B2(new_n201), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n212), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n262), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT10), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n312), .A2(new_n313), .A3(new_n322), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n311), .A2(KEYINPUT10), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n232), .A2(new_n199), .A3(new_n203), .A4(new_n250), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n330), .A2(new_n328), .A3(new_n322), .A4(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT86), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(G110), .B(G140), .ZN(new_n335));
  INV_X1    g149(.A(G227), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n336), .A2(G953), .ZN(new_n337));
  XOR2_X1   g151(.A(new_n335), .B(new_n337), .Z(new_n338));
  NAND2_X1  g152(.A1(new_n210), .A2(new_n212), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n326), .B1(new_n339), .B2(new_n262), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT12), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n322), .A2(KEYINPUT87), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n341), .B1(new_n340), .B2(new_n342), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n334), .A2(new_n338), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n312), .A2(new_n328), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n321), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n338), .B1(new_n334), .B2(new_n349), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n307), .B(new_n308), .C1(new_n347), .C2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(G469), .A2(G902), .ZN(new_n352));
  INV_X1    g166(.A(new_n338), .ZN(new_n353));
  INV_X1    g167(.A(new_n334), .ZN(new_n354));
  INV_X1    g168(.A(new_n345), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n353), .B1(new_n329), .B2(new_n333), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n349), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(G469), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n351), .A2(new_n352), .A3(new_n359), .ZN(new_n360));
  XOR2_X1   g174(.A(KEYINPUT9), .B(G234), .Z(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(G221), .B1(new_n362), .B2(G902), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G217), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n362), .A2(new_n365), .A3(G953), .ZN(new_n366));
  XNOR2_X1  g180(.A(G116), .B(G122), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n221), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n235), .A2(KEYINPUT14), .A3(G122), .ZN(new_n369));
  INV_X1    g183(.A(new_n367), .ZN(new_n370));
  OAI211_X1 g184(.A(G107), .B(new_n369), .C1(new_n370), .C2(KEYINPUT14), .ZN(new_n371));
  INV_X1    g185(.A(G128), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT68), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT68), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G128), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n187), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n372), .A2(G143), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT98), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT98), .ZN(new_n379));
  INV_X1    g193(.A(new_n377), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n379), .B(new_n380), .C1(new_n206), .C2(new_n187), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n378), .A2(new_n314), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n314), .B1(new_n378), .B2(new_n381), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n368), .B(new_n371), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n378), .A2(new_n314), .A3(new_n381), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n377), .A2(KEYINPUT13), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n386), .B1(new_n206), .B2(new_n187), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n377), .A2(KEYINPUT13), .ZN(new_n388));
  OAI21_X1  g202(.A(G134), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n367), .B(new_n221), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n385), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n366), .B1(new_n384), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n384), .A2(new_n391), .A3(new_n366), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n308), .ZN(new_n396));
  INV_X1    g210(.A(G478), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n397), .A2(KEYINPUT15), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n396), .B(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G475), .ZN(new_n400));
  INV_X1    g214(.A(G237), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n216), .A3(G214), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n187), .ZN(new_n403));
  NOR2_X1   g217(.A1(G237), .A2(G953), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(G143), .A3(G214), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  AND2_X1   g220(.A1(KEYINPUT18), .A2(G131), .ZN(new_n407));
  XOR2_X1   g221(.A(new_n406), .B(new_n407), .Z(new_n408));
  INV_X1    g222(.A(KEYINPUT79), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n409), .B(G140), .C1(new_n211), .C2(KEYINPUT78), .ZN(new_n410));
  INV_X1    g224(.A(G140), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT79), .B1(new_n411), .B2(G125), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(G125), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n410), .B(new_n412), .C1(KEYINPUT78), .C2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G146), .ZN(new_n415));
  XNOR2_X1  g229(.A(G125), .B(G140), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n195), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n415), .A2(KEYINPUT96), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT96), .B1(new_n415), .B2(new_n417), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n408), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(G113), .B(G122), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(new_n255), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT80), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n424), .B1(new_n413), .B2(KEYINPUT16), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT16), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n426), .A2(new_n411), .A3(KEYINPUT80), .A4(G125), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n425), .B(new_n427), .C1(new_n414), .C2(new_n426), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n191), .ZN(new_n429));
  OR2_X1    g243(.A1(new_n413), .A2(KEYINPUT78), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n430), .A2(KEYINPUT16), .A3(new_n412), .A4(new_n410), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n431), .A2(G146), .A3(new_n425), .A4(new_n427), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n406), .A2(KEYINPUT17), .A3(G131), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n406), .A2(G131), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT17), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n403), .A2(new_n320), .A3(new_n405), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n429), .A2(new_n432), .A3(new_n433), .A4(new_n437), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n421), .A2(new_n423), .A3(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n414), .A2(KEYINPUT19), .B1(new_n416), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n195), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n434), .A2(new_n436), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(new_n432), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n423), .B1(new_n421), .B2(new_n444), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n400), .B(new_n308), .C1(new_n439), .C2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n421), .A2(new_n423), .A3(new_n438), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n406), .B(new_n407), .ZN(new_n450));
  INV_X1    g264(.A(new_n420), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n450), .B1(new_n451), .B2(new_n418), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n442), .A2(new_n432), .A3(new_n443), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n449), .B1(new_n454), .B2(new_n423), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n455), .A2(KEYINPUT20), .A3(new_n400), .A4(new_n308), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n423), .B1(new_n421), .B2(new_n438), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n308), .B1(new_n439), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G475), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n448), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n399), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n216), .A2(G952), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n462), .B1(G234), .B2(G237), .ZN(new_n463));
  XOR2_X1   g277(.A(KEYINPUT21), .B(G898), .Z(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(G234), .A2(G237), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(G902), .A3(G953), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n463), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n461), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n364), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n306), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT99), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT24), .B(G110), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n475), .B(KEYINPUT77), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n233), .A2(G128), .ZN(new_n477));
  OAI211_X1 g291(.A(KEYINPUT75), .B(new_n477), .C1(new_n206), .C2(new_n233), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT76), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n233), .B1(new_n373), .B2(new_n375), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n478), .B(new_n479), .C1(new_n481), .C2(KEYINPUT75), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n477), .A2(KEYINPUT75), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n206), .A2(KEYINPUT75), .A3(new_n233), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT76), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n476), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n373), .A2(new_n375), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(KEYINPUT23), .A3(G119), .ZN(new_n489));
  INV_X1    g303(.A(G110), .ZN(new_n490));
  AOI21_X1  g304(.A(KEYINPUT23), .B1(new_n372), .B2(G119), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n489), .A2(new_n490), .A3(new_n477), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT81), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n491), .B1(new_n480), .B2(KEYINPUT23), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT81), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n495), .A2(new_n496), .A3(new_n490), .A4(new_n477), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n432), .B(new_n417), .C1(new_n487), .C2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT82), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n429), .A2(new_n432), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n482), .A2(new_n486), .A3(new_n476), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n495), .A2(new_n477), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(G110), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n501), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n499), .A2(new_n500), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n216), .A2(G221), .A3(G234), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(KEYINPUT22), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(G137), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n500), .B1(new_n499), .B2(new_n505), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI211_X1 g327(.A(new_n500), .B(new_n510), .C1(new_n499), .C2(new_n505), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n308), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT83), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT25), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n499), .A2(new_n505), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT82), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(new_n506), .A3(new_n510), .ZN(new_n522));
  INV_X1    g336(.A(new_n514), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n524), .A2(new_n516), .A3(new_n517), .A4(new_n308), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n365), .B1(G234), .B2(new_n308), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n519), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT84), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n526), .A2(G902), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n522), .A2(new_n523), .A3(KEYINPUT84), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT31), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n248), .A2(new_n245), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT30), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT66), .B1(new_n317), .B2(G134), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT66), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(new_n314), .A3(G137), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n317), .A2(G134), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n538), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G131), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT67), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n319), .A2(new_n320), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT67), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n542), .A2(new_n546), .A3(G131), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT70), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT70), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n544), .A2(new_n550), .A3(new_n545), .A4(new_n547), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n339), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n321), .A2(new_n199), .A3(new_n203), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n537), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n210), .A2(new_n212), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n553), .B(new_n537), .C1(new_n555), .C2(new_n548), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n536), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n552), .A2(new_n535), .A3(new_n553), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n559), .A2(KEYINPUT71), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT71), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n562), .B(new_n536), .C1(new_n554), .C2(new_n557), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(G101), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n404), .A2(G210), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n534), .B1(new_n564), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n568), .ZN(new_n570));
  AOI211_X1 g384(.A(KEYINPUT31), .B(new_n570), .C1(new_n561), .C2(new_n563), .ZN(new_n571));
  OR2_X1    g385(.A1(new_n559), .A2(KEYINPUT28), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n559), .A2(KEYINPUT28), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n553), .B1(new_n555), .B2(new_n548), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n572), .A2(new_n573), .B1(new_n536), .B2(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n568), .B(KEYINPUT72), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n569), .A2(new_n571), .A3(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(G472), .A2(G902), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT32), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n564), .A2(new_n568), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT31), .ZN(new_n583));
  INV_X1    g397(.A(new_n577), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n564), .A2(new_n534), .A3(new_n568), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT32), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(new_n587), .A3(new_n579), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n581), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(KEYINPUT73), .B1(new_n564), .B2(new_n568), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT73), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n561), .A2(new_n591), .A3(new_n570), .A4(new_n563), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT29), .B1(new_n575), .B2(new_n576), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n590), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n535), .B1(new_n552), .B2(new_n553), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n595), .B1(new_n572), .B2(new_n573), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n596), .A2(KEYINPUT29), .A3(new_n568), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT74), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n596), .A2(KEYINPUT74), .A3(KEYINPUT29), .A4(new_n568), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n594), .A2(new_n308), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(G472), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n533), .B1(new_n589), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT99), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n306), .A2(new_n472), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n474), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT100), .B(G101), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G3));
  INV_X1    g422(.A(G472), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n609), .B1(new_n586), .B2(new_n308), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n578), .A2(new_n580), .ZN(new_n611));
  NOR4_X1   g425(.A1(new_n610), .A2(new_n611), .A3(new_n364), .A4(new_n533), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n296), .A2(new_n298), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n300), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT101), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT101), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n613), .A2(new_n616), .A3(new_n300), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n615), .A2(new_n470), .A3(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n397), .A2(new_n308), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n384), .A2(new_n391), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT102), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(new_n394), .A3(new_n393), .ZN(new_n624));
  INV_X1    g438(.A(new_n394), .ZN(new_n625));
  AOI21_X1  g439(.A(KEYINPUT102), .B1(new_n384), .B2(new_n391), .ZN(new_n626));
  OAI22_X1  g440(.A1(new_n625), .A2(new_n392), .B1(new_n626), .B2(new_n620), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n619), .B1(new_n628), .B2(G478), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n395), .A2(new_n397), .A3(new_n308), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n460), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT103), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n618), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n612), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT34), .B(G104), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G6));
  INV_X1    g452(.A(new_n399), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n460), .ZN(new_n640));
  AND4_X1   g454(.A1(new_n470), .A2(new_n615), .A3(new_n617), .A4(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n612), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT35), .B(G107), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT104), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n642), .B(new_n644), .ZN(G9));
  NOR2_X1   g459(.A1(new_n610), .A2(new_n611), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n510), .A2(KEYINPUT36), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n520), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n530), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n527), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n474), .A2(new_n605), .A3(new_n646), .A4(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(new_n490), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT105), .B(KEYINPUT37), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G12));
  NOR3_X1   g468(.A1(new_n578), .A2(KEYINPUT32), .A3(new_n580), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n587), .B1(new_n586), .B2(new_n579), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n602), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n615), .A2(new_n617), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT106), .B(G900), .Z(new_n659));
  AOI21_X1  g473(.A(new_n463), .B1(new_n468), .B2(new_n659), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n639), .A2(new_n460), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n650), .A2(new_n363), .A3(new_n360), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n657), .A2(new_n658), .A3(new_n661), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G128), .ZN(G30));
  INV_X1    g479(.A(new_n364), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n660), .B(KEYINPUT39), .Z(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n668), .A2(KEYINPUT40), .ZN(new_n669));
  INV_X1    g483(.A(new_n582), .ZN(new_n670));
  INV_X1    g484(.A(new_n595), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n576), .B1(new_n671), .B2(new_n559), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n308), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(G472), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n674), .B1(new_n655), .B2(new_n656), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n299), .A2(new_n301), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT38), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n676), .A2(new_n678), .A3(new_n650), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n639), .A2(new_n632), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n300), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT107), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT107), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n679), .A2(new_n686), .A3(new_n683), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n669), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n668), .A2(KEYINPUT40), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G143), .ZN(G45));
  INV_X1    g505(.A(new_n660), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n629), .A2(new_n460), .A3(new_n630), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT108), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n657), .A2(new_n658), .A3(new_n663), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G146), .ZN(G48));
  NAND2_X1  g510(.A1(new_n334), .A2(new_n349), .ZN(new_n697));
  AOI22_X1  g511(.A1(new_n697), .A2(new_n353), .B1(new_n357), .B2(new_n345), .ZN(new_n698));
  OAI21_X1  g512(.A(G469), .B1(new_n698), .B2(G902), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n699), .A2(new_n363), .A3(new_n351), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(KEYINPUT109), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n699), .A2(new_n702), .A3(new_n363), .A4(new_n351), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n603), .A2(new_n635), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT110), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  INV_X1    g523(.A(new_n533), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n641), .A2(new_n657), .A3(new_n710), .A4(new_n705), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G116), .ZN(G18));
  AND4_X1   g526(.A1(new_n617), .A2(new_n701), .A3(new_n615), .A4(new_n703), .ZN(new_n713));
  INV_X1    g527(.A(new_n471), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n713), .A2(new_n657), .A3(new_n714), .A4(new_n650), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G119), .ZN(G21));
  NOR2_X1   g530(.A1(new_n704), .A2(new_n681), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n533), .B(KEYINPUT112), .ZN(new_n718));
  INV_X1    g532(.A(new_n618), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n586), .A2(new_n308), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n596), .A2(new_n576), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n583), .A2(new_n585), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n579), .B(KEYINPUT111), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n720), .A2(G472), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n717), .A2(new_n718), .A3(new_n719), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  OAI21_X1  g540(.A(G472), .B1(new_n578), .B2(G902), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n722), .A2(new_n723), .ZN(new_n728));
  AND4_X1   g542(.A1(new_n727), .A2(new_n694), .A3(new_n650), .A4(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n713), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G125), .ZN(G27));
  AND3_X1   g545(.A1(new_n657), .A2(new_n718), .A3(KEYINPUT42), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n633), .A2(KEYINPUT108), .A3(new_n692), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n693), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n733), .A2(new_n677), .A3(new_n300), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n352), .B(KEYINPUT113), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n351), .A2(new_n359), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT114), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT114), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n351), .A2(new_n359), .A3(new_n740), .A4(new_n737), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n739), .A2(new_n363), .A3(new_n741), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n736), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n657), .A3(new_n710), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT42), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n732), .A2(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n320), .ZN(G33));
  NAND2_X1  g561(.A1(new_n677), .A2(new_n300), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  AND4_X1   g563(.A1(new_n363), .A2(new_n739), .A3(new_n661), .A4(new_n741), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n603), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G134), .ZN(G36));
  NAND2_X1  g566(.A1(new_n356), .A2(new_n358), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n356), .A2(KEYINPUT45), .A3(new_n358), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(G469), .A3(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT46), .ZN(new_n759));
  INV_X1    g573(.A(new_n737), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(KEYINPUT46), .B1(new_n757), .B2(new_n737), .ZN(new_n762));
  INV_X1    g576(.A(new_n351), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n765), .A2(new_n363), .A3(new_n667), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT44), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n631), .A2(KEYINPUT43), .A3(new_n460), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n460), .B(KEYINPUT115), .ZN(new_n769));
  INV_X1    g583(.A(new_n631), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n768), .B1(new_n771), .B2(KEYINPUT43), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n772), .B(new_n650), .C1(new_n611), .C2(new_n610), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n766), .B1(new_n767), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n749), .B1(new_n773), .B2(new_n767), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT116), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n775), .A2(KEYINPUT116), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n774), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G137), .ZN(G39));
  INV_X1    g593(.A(new_n363), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n764), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT47), .ZN(new_n782));
  INV_X1    g596(.A(new_n736), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n657), .A2(new_n710), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G140), .ZN(G42));
  INV_X1    g600(.A(KEYINPUT120), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n718), .A2(new_n724), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n772), .A2(new_n463), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n705), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n678), .A2(new_n682), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(KEYINPUT50), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT50), .B1(new_n792), .B2(new_n794), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n787), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n797), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(new_n795), .A3(KEYINPUT120), .ZN(new_n800));
  INV_X1    g614(.A(new_n789), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n704), .A2(new_n748), .ZN(new_n802));
  AND4_X1   g616(.A1(new_n650), .A2(new_n801), .A3(new_n724), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n676), .A2(new_n463), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n710), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n804), .A2(new_n770), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n803), .B1(new_n806), .B2(new_n632), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n699), .A2(new_n351), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n363), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n749), .B(new_n790), .C1(new_n782), .C2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n798), .A2(new_n800), .A3(new_n807), .A4(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT51), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n810), .A2(new_n807), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n812), .B1(new_n799), .B2(new_n795), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n462), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n790), .A2(new_n713), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n657), .A2(new_n718), .ZN(new_n818));
  NOR4_X1   g632(.A1(new_n818), .A2(new_n704), .A3(new_n748), .A4(new_n789), .ZN(new_n819));
  XOR2_X1   g633(.A(new_n819), .B(KEYINPUT48), .Z(new_n820));
  NAND4_X1  g634(.A1(new_n813), .A2(new_n816), .A3(new_n817), .A4(new_n820), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n640), .A2(new_n633), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n612), .A2(new_n306), .A3(new_n470), .A4(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n651), .A2(new_n606), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n706), .A2(new_n715), .A3(new_n725), .A4(new_n711), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n824), .A2(new_n746), .A3(new_n825), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n399), .A2(new_n460), .A3(new_n660), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n657), .A2(new_n663), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n742), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n829), .A2(new_n724), .A3(new_n650), .A4(new_n694), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n748), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n603), .A2(new_n749), .A3(new_n750), .ZN(new_n832));
  OAI21_X1  g646(.A(KEYINPUT117), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n662), .B1(new_n589), .B2(new_n602), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n835), .A2(new_n827), .B1(new_n729), .B2(new_n829), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n834), .B(new_n751), .C1(new_n836), .C2(new_n748), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n615), .A2(new_n617), .A3(new_n680), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n527), .A2(new_n649), .A3(new_n692), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT118), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n527), .A2(new_n842), .A3(new_n649), .A4(new_n692), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n675), .A2(new_n829), .A3(new_n839), .A4(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n664), .A2(new_n695), .A3(new_n845), .A4(new_n730), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n835), .B(new_n658), .C1(new_n661), .C2(new_n694), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(KEYINPUT52), .A3(new_n730), .A4(new_n845), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  AND4_X1   g665(.A1(KEYINPUT53), .A2(new_n826), .A3(new_n838), .A4(new_n851), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n833), .A2(new_n837), .B1(new_n848), .B2(new_n850), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT53), .B1(new_n853), .B2(new_n826), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT54), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  OR3_X1    g669(.A1(new_n804), .A2(new_n634), .A3(new_n805), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n838), .A2(new_n851), .ZN(new_n858));
  INV_X1    g672(.A(new_n746), .ZN(new_n859));
  INV_X1    g673(.A(new_n825), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n606), .A2(new_n823), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n859), .A2(new_n860), .A3(new_n861), .A4(new_n651), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n857), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n853), .A2(KEYINPUT53), .A3(new_n826), .ZN(new_n864));
  XNOR2_X1  g678(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n855), .A2(new_n856), .A3(new_n867), .ZN(new_n868));
  OAI22_X1  g682(.A1(new_n821), .A2(new_n868), .B1(G952), .B2(G953), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n808), .A2(KEYINPUT49), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n678), .A2(new_n770), .A3(new_n769), .A4(new_n870), .ZN(new_n871));
  AOI211_X1 g685(.A(new_n675), .B(new_n871), .C1(KEYINPUT49), .C2(new_n808), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n872), .A2(new_n300), .A3(new_n363), .A4(new_n718), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n869), .A2(new_n873), .ZN(G75));
  AOI21_X1  g688(.A(new_n308), .B1(new_n863), .B2(new_n864), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(G210), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT56), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n271), .B1(new_n275), .B2(new_n276), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(new_n220), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT55), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n876), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n880), .B1(new_n876), .B2(new_n877), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n216), .A2(G952), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(G51));
  NOR2_X1   g698(.A1(new_n737), .A2(KEYINPUT57), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n865), .B1(new_n852), .B2(new_n854), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n885), .B1(new_n886), .B2(new_n867), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n737), .A2(KEYINPUT57), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n698), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n875), .A2(new_n758), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n883), .B1(new_n891), .B2(new_n892), .ZN(G54));
  NAND3_X1  g707(.A1(new_n875), .A2(KEYINPUT58), .A3(G475), .ZN(new_n894));
  INV_X1    g708(.A(new_n455), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n896), .A2(new_n897), .A3(new_n883), .ZN(G60));
  INV_X1    g712(.A(new_n883), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n619), .B(KEYINPUT59), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n855), .B2(new_n867), .ZN(new_n901));
  INV_X1    g715(.A(new_n628), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n900), .B1(new_n886), .B2(new_n867), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n903), .B1(new_n902), .B2(new_n904), .ZN(G63));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n906));
  NAND2_X1  g720(.A1(G217), .A2(G902), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT60), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(new_n852), .B2(new_n854), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n529), .A2(new_n531), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n883), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n908), .B1(new_n863), .B2(new_n864), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n648), .B(KEYINPUT121), .Z(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n906), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  OR2_X1    g730(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n917));
  INV_X1    g731(.A(new_n911), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n899), .B(new_n917), .C1(new_n913), .C2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n912), .B2(KEYINPUT123), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n915), .B(KEYINPUT122), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n916), .B1(new_n921), .B2(new_n922), .ZN(G66));
  NAND3_X1  g737(.A1(new_n860), .A2(new_n861), .A3(new_n651), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n216), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT124), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n216), .B1(new_n215), .B2(new_n464), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n878), .B1(G898), .B2(new_n216), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT125), .Z(new_n930));
  XNOR2_X1  g744(.A(new_n928), .B(new_n930), .ZN(G69));
  NAND3_X1  g745(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n554), .A2(new_n557), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT126), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(new_n441), .Z(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n785), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n849), .A2(new_n730), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n938), .B1(new_n688), .B2(new_n689), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n937), .B1(new_n940), .B2(KEYINPUT62), .ZN(new_n941));
  INV_X1    g755(.A(new_n778), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT62), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n942), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n668), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n603), .A2(new_n945), .A3(new_n749), .A4(new_n822), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n941), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n932), .B(new_n936), .C1(new_n947), .C2(G953), .ZN(new_n948));
  INV_X1    g762(.A(new_n839), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n766), .A2(new_n818), .A3(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n950), .A2(new_n938), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n746), .A2(new_n832), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n785), .A2(new_n778), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n216), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n336), .A2(G900), .A3(G953), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n954), .A2(new_n935), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n948), .A2(new_n956), .ZN(G72));
  INV_X1    g771(.A(new_n924), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n941), .A2(new_n944), .A3(new_n958), .A4(new_n946), .ZN(new_n959));
  XNOR2_X1  g773(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n960));
  NAND2_X1  g774(.A1(G472), .A2(G902), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(new_n962));
  AOI211_X1 g776(.A(new_n570), .B(new_n564), .C1(new_n959), .C2(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n962), .B1(new_n953), .B2(new_n924), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n964), .A2(new_n570), .A3(new_n564), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n590), .A2(new_n582), .A3(new_n592), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n962), .B(new_n966), .C1(new_n852), .C2(new_n854), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n965), .A2(new_n899), .A3(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n963), .A2(new_n968), .ZN(G57));
endmodule


