//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n621, new_n623, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191, new_n1192, new_n1193, new_n1194;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT65), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  OR2_X1    g029(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT66), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  AOI22_X1  g032(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT67), .Z(G319));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G137), .ZN(new_n464));
  OR3_X1    g039(.A1(new_n462), .A2(KEYINPUT68), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g040(.A(KEYINPUT68), .B1(new_n462), .B2(new_n464), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n462), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n463), .A2(G2104), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n470), .A2(G2105), .B1(G101), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  OAI21_X1  g049(.A(G2104), .B1(new_n463), .B2(G112), .ZN(new_n475));
  INV_X1    g050(.A(G100), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(new_n463), .ZN(new_n477));
  XNOR2_X1  g052(.A(KEYINPUT3), .B(G2104), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n478), .B(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(new_n463), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n477), .B1(new_n481), .B2(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n480), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  OAI21_X1  g061(.A(G2104), .B1(new_n463), .B2(G114), .ZN(new_n487));
  NOR2_X1   g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT70), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n490), .A2(new_n492), .A3(new_n493), .A4(G2104), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(G126), .A2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n460), .ZN(new_n497));
  INV_X1    g072(.A(new_n461), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n502), .B(new_n503), .C1(new_n461), .C2(new_n460), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n503), .B1(new_n478), .B2(new_n502), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n495), .B(new_n500), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n510), .A2(G543), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n520), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n516), .A2(new_n520), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n519), .A2(new_n525), .ZN(G166));
  INV_X1    g101(.A(new_n523), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G89), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n529));
  XOR2_X1   g104(.A(KEYINPUT74), .B(KEYINPUT7), .Z(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n530), .B(new_n531), .ZN(new_n532));
  XOR2_X1   g107(.A(KEYINPUT73), .B(G51), .Z(new_n533));
  NAND2_X1  g108(.A1(new_n521), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n528), .A2(new_n529), .A3(new_n532), .A4(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  NAND2_X1  g111(.A1(new_n521), .A2(G52), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n523), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT75), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(new_n518), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  NAND3_X1  g119(.A1(new_n516), .A2(G81), .A3(new_n520), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n521), .A2(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(KEYINPUT76), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT76), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n545), .A2(new_n549), .A3(new_n546), .ZN(new_n550));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n514), .A2(new_n515), .ZN(new_n552));
  INV_X1    g127(.A(G56), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n548), .A2(new_n550), .B1(G651), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND3_X1  g135(.A1(new_n521), .A2(KEYINPUT9), .A3(G53), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n520), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT77), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n552), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n527), .A2(G91), .B1(new_n570), .B2(G651), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n567), .A2(new_n571), .ZN(G299));
  OAI221_X1 g147(.A(new_n522), .B1(new_n523), .B2(new_n524), .C1(new_n517), .C2(new_n518), .ZN(G303));
  OAI21_X1  g148(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n516), .A2(G87), .A3(new_n520), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n521), .A2(G49), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  NAND3_X1  g152(.A1(new_n514), .A2(G61), .A3(new_n515), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G651), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n514), .A2(G86), .A3(new_n515), .A4(new_n520), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n520), .A2(G48), .A3(G543), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n581), .A2(new_n585), .ZN(G305));
  NAND2_X1  g161(.A1(G72), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G60), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n552), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G651), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(KEYINPUT78), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(KEYINPUT78), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n527), .A2(G85), .B1(G47), .B2(new_n521), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(KEYINPUT79), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(KEYINPUT79), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(G290));
  INV_X1    g172(.A(KEYINPUT80), .ZN(new_n598));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(G171), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(G301), .A2(KEYINPUT80), .A3(G868), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n516), .A2(G92), .A3(new_n520), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n602), .B(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(G79), .ZN(new_n605));
  OAI21_X1  g180(.A(KEYINPUT81), .B1(new_n605), .B2(new_n512), .ZN(new_n606));
  OR3_X1    g181(.A1(new_n605), .A2(new_n512), .A3(KEYINPUT81), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n606), .B(new_n607), .C1(new_n552), .C2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n609), .A2(G651), .B1(G54), .B2(new_n521), .ZN(new_n610));
  AND2_X1   g185(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  OAI211_X1 g186(.A(new_n600), .B(new_n601), .C1(G868), .C2(new_n611), .ZN(G284));
  OAI211_X1 g187(.A(new_n600), .B(new_n601), .C1(G868), .C2(new_n611), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT77), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n566), .B(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n571), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n614), .B1(new_n618), .B2(G868), .ZN(G297));
  OAI21_X1  g194(.A(new_n614), .B1(new_n618), .B2(G868), .ZN(G280));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n611), .B1(new_n621), .B2(G860), .ZN(G148));
  NOR2_X1   g197(.A1(new_n555), .A2(G868), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n611), .A2(new_n621), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(G868), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT82), .Z(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n478), .A2(new_n471), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT12), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(G2100), .Z(new_n631));
  NAND2_X1  g206(.A1(new_n483), .A2(G135), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n481), .A2(G123), .ZN(new_n633));
  NOR2_X1   g208(.A1(G99), .A2(G2105), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(new_n463), .B2(G111), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(G2096), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n631), .A2(new_n638), .ZN(G156));
  XOR2_X1   g214(.A(KEYINPUT15), .B(G2435), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT85), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT84), .B(KEYINPUT14), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n641), .A2(new_n643), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(G14), .B1(new_n652), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n656), .B2(new_n652), .ZN(G401));
  XNOR2_X1  g233(.A(G2072), .B(G2078), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT17), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  OR3_X1    g239(.A1(new_n661), .A2(new_n659), .A3(new_n662), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n661), .A2(new_n659), .A3(new_n662), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT18), .Z(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(new_n637), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2100), .ZN(G227));
  XNOR2_X1  g246(.A(G1961), .B(G1966), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT86), .ZN(new_n673));
  XOR2_X1   g248(.A(G1956), .B(G2474), .Z(new_n674));
  OR2_X1    g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n673), .A2(new_n674), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n679), .A2(new_n677), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n678), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n675), .A2(new_n677), .A3(new_n679), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1981), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n688), .B(new_n690), .ZN(G229));
  INV_X1    g266(.A(G16), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G24), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT89), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(G290), .B2(G16), .ZN(new_n696));
  INV_X1    g271(.A(G1986), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G25), .ZN(new_n700));
  OR2_X1    g275(.A1(G95), .A2(G2105), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n701), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT88), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n481), .B2(G119), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n483), .A2(G131), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n700), .B1(new_n707), .B2(new_n699), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT35), .B(G1991), .Z(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n708), .B(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(KEYINPUT94), .B2(KEYINPUT36), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n696), .A2(new_n697), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n698), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n692), .A2(G23), .ZN(new_n715));
  INV_X1    g290(.A(G288), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n692), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT33), .Z(new_n718));
  INV_X1    g293(.A(G1976), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n692), .A2(G6), .ZN(new_n721));
  INV_X1    g296(.A(G305), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(new_n692), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT90), .Z(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT32), .B(G1981), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n692), .A2(G22), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT91), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G166), .B2(new_n692), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT92), .B(G1971), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n720), .A2(new_n726), .A3(new_n727), .A4(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT34), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n714), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(KEYINPUT93), .B1(new_n733), .B2(KEYINPUT34), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n726), .A2(new_n727), .A3(new_n732), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n718), .B(G1976), .ZN(new_n739));
  OAI211_X1 g314(.A(KEYINPUT93), .B(KEYINPUT34), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n736), .B1(new_n737), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI221_X1 g319(.A(new_n736), .B1(KEYINPUT94), .B2(KEYINPUT36), .C1(new_n737), .C2(new_n741), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n692), .A2(G5), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G171), .B2(new_n692), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT101), .ZN(new_n748));
  INV_X1    g323(.A(G1961), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n692), .A2(G20), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT23), .Z(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G299), .B2(G16), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT102), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(G1956), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n692), .A2(G19), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n555), .B2(new_n692), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT95), .B(G1341), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n699), .A2(G32), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n481), .A2(G129), .ZN(new_n762));
  NAND3_X1  g337(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT26), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n765), .A2(new_n766), .B1(G105), .B2(new_n471), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n762), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n483), .A2(G141), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n761), .B1(new_n771), .B2(new_n699), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT27), .B(G1996), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n699), .A2(G27), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G164), .B2(new_n699), .ZN(new_n777));
  INV_X1    g352(.A(G2078), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n757), .A2(new_n759), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n772), .A2(new_n774), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n750), .A2(new_n755), .A3(new_n760), .A4(new_n783), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n483), .A2(G139), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT25), .Z(new_n787));
  AOI22_X1  g362(.A1(new_n478), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(new_n463), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n790), .A2(new_n699), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n699), .B2(G33), .ZN(new_n792));
  INV_X1    g367(.A(G2072), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT98), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n611), .A2(new_n692), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G4), .B2(new_n692), .ZN(new_n797));
  INV_X1    g372(.A(G1348), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n699), .A2(G26), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT28), .Z(new_n801));
  NAND2_X1  g376(.A1(new_n483), .A2(G140), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n481), .A2(G128), .ZN(new_n803));
  OAI21_X1  g378(.A(KEYINPUT96), .B1(G104), .B2(G2105), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  NOR3_X1   g380(.A1(KEYINPUT96), .A2(G104), .A3(G2105), .ZN(new_n806));
  OAI221_X1 g381(.A(G2104), .B1(G116), .B2(new_n463), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n802), .A2(new_n803), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n801), .B1(new_n808), .B2(G29), .ZN(new_n809));
  INV_X1    g384(.A(G2067), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n795), .A2(new_n799), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n792), .A2(new_n793), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT97), .B(KEYINPUT24), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(G34), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(new_n699), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n473), .B2(new_n699), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G2084), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n636), .A2(new_n699), .ZN(new_n819));
  INV_X1    g394(.A(G28), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n820), .A2(KEYINPUT30), .ZN(new_n821));
  AOI21_X1  g396(.A(G29), .B1(new_n820), .B2(KEYINPUT30), .ZN(new_n822));
  OR2_X1    g397(.A1(KEYINPUT31), .A2(G11), .ZN(new_n823));
  NAND2_X1  g398(.A1(KEYINPUT31), .A2(G11), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n821), .A2(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n813), .A2(new_n818), .A3(new_n819), .A4(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(new_n797), .B2(new_n798), .ZN(new_n827));
  NOR2_X1   g402(.A1(G286), .A2(new_n692), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT99), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(G16), .B2(G21), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT100), .B(G1966), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n830), .B(new_n831), .Z(new_n832));
  NAND3_X1  g407(.A1(new_n812), .A2(new_n827), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n699), .A2(G35), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(G162), .B2(new_n699), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT29), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G2090), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n784), .A2(new_n833), .A3(new_n837), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n744), .A2(new_n745), .A3(new_n838), .ZN(G311));
  NAND3_X1  g414(.A1(new_n744), .A2(new_n745), .A3(new_n838), .ZN(G150));
  AOI22_X1  g415(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(new_n518), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n521), .A2(G55), .ZN(new_n843));
  INV_X1    g418(.A(G93), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n843), .B1(new_n523), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n548), .A2(new_n550), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n554), .A2(G651), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n555), .A2(new_n846), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT38), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n611), .A2(G559), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n856));
  AOI21_X1  g431(.A(G860), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n856), .B2(new_n855), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n847), .A2(G860), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT37), .Z(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(G145));
  INV_X1    g436(.A(KEYINPUT40), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT103), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n770), .A2(new_n808), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n770), .A2(new_n808), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n864), .A2(G164), .A3(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(G164), .B1(new_n864), .B2(new_n865), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n863), .B(new_n790), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n790), .A2(new_n863), .ZN(new_n871));
  OAI21_X1  g446(.A(KEYINPUT103), .B1(new_n785), .B2(new_n789), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .A4(new_n866), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n706), .B(KEYINPUT104), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n875), .A2(new_n629), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n629), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n483), .A2(G142), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n481), .A2(G130), .ZN(new_n880));
  OR2_X1    g455(.A1(G106), .A2(G2105), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n881), .B(G2104), .C1(G118), .C2(new_n463), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n878), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n876), .A2(new_n883), .A3(new_n877), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n874), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n485), .B(new_n473), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n636), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n869), .A2(new_n873), .A3(new_n885), .A4(new_n886), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(G37), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n890), .B1(new_n888), .B2(new_n891), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n862), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n895), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n897), .A2(KEYINPUT40), .A3(new_n893), .A4(new_n892), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n896), .A2(new_n898), .ZN(G395));
  XNOR2_X1  g474(.A(G303), .B(G288), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n595), .A2(G305), .A3(new_n596), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(G305), .B1(new_n595), .B2(new_n596), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n901), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n904), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n906), .A2(new_n900), .A3(new_n902), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT42), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n611), .A2(G299), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n604), .A2(new_n610), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(new_n571), .A3(new_n567), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT41), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT105), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n914), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n910), .A2(KEYINPUT41), .A3(new_n912), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n915), .B1(new_n918), .B2(KEYINPUT105), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n852), .B(new_n624), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n920), .A2(new_n913), .ZN(new_n922));
  OR3_X1    g497(.A1(new_n921), .A2(KEYINPUT106), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT106), .B1(new_n921), .B2(new_n922), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n909), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n909), .A2(new_n924), .ZN(new_n926));
  OAI21_X1  g501(.A(G868), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n927), .B1(G868), .B2(new_n846), .ZN(G295));
  OAI21_X1  g503(.A(new_n927), .B1(G868), .B2(new_n846), .ZN(G331));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n905), .A2(new_n907), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n850), .A2(new_n851), .A3(G301), .ZN(new_n932));
  AOI21_X1  g507(.A(G301), .B1(new_n850), .B2(new_n851), .ZN(new_n933));
  OAI21_X1  g508(.A(G286), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n852), .A2(G171), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n850), .A2(G301), .A3(new_n851), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(G168), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n934), .A2(new_n937), .A3(new_n918), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  AOI22_X1  g514(.A1(new_n934), .A2(new_n937), .B1(new_n910), .B2(new_n912), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n931), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(new_n916), .B2(new_n917), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n937), .B(new_n934), .C1(new_n943), .C2(new_n915), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n934), .A2(new_n937), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n913), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n944), .A2(new_n946), .A3(new_n908), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n941), .A2(new_n947), .A3(new_n893), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n944), .A2(new_n946), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n931), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT43), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n951), .A2(new_n952), .A3(new_n893), .A4(new_n947), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n930), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n951), .A2(new_n893), .A3(new_n947), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n947), .A2(new_n952), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n946), .A2(new_n938), .ZN(new_n957));
  AOI21_X1  g532(.A(G37), .B1(new_n957), .B2(new_n931), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n955), .A2(KEYINPUT43), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n954), .B1(new_n930), .B2(new_n959), .ZN(G397));
  INV_X1    g535(.A(G1384), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n507), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n467), .A2(new_n472), .A3(G40), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(G290), .A2(G1986), .A3(new_n966), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n595), .A2(new_n697), .A3(new_n596), .A4(new_n966), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  XOR2_X1   g544(.A(new_n969), .B(KEYINPUT107), .Z(new_n970));
  NOR2_X1   g545(.A1(new_n707), .A2(new_n709), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n706), .A2(new_n710), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n966), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n808), .B(G2067), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n966), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n975), .B(KEYINPUT108), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n771), .A2(G1996), .ZN(new_n977));
  INV_X1    g552(.A(G1996), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n770), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n977), .A2(new_n966), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n976), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n970), .A2(new_n973), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G1981), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n581), .A2(new_n585), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT111), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n518), .B1(new_n578), .B2(new_n579), .ZN(new_n987));
  OAI21_X1  g562(.A(G1981), .B1(new_n987), .B2(new_n584), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n985), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(G305), .A2(KEYINPUT111), .A3(G1981), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT49), .ZN(new_n992));
  INV_X1    g567(.A(G8), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT109), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n502), .B1(new_n460), .B2(new_n461), .ZN(new_n995));
  INV_X1    g570(.A(new_n503), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n499), .B1(new_n997), .B2(new_n504), .ZN(new_n998));
  AOI211_X1 g573(.A(new_n994), .B(G1384), .C1(new_n998), .C2(new_n495), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT109), .B1(new_n507), .B2(new_n961), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n965), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n993), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT49), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n989), .A2(new_n1004), .A3(new_n990), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n992), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1006), .A2(new_n719), .A3(new_n716), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n985), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n1009));
  AOI21_X1  g584(.A(G1384), .B1(new_n998), .B2(new_n495), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT50), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n962), .A2(KEYINPUT110), .A3(KEYINPUT50), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n962), .A2(new_n994), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n507), .A2(KEYINPUT109), .A3(new_n961), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1015), .A2(new_n1011), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G2090), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1014), .A2(new_n1017), .A3(new_n1018), .A4(new_n1002), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1010), .A2(KEYINPUT45), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n964), .A2(new_n1020), .A3(new_n1002), .ZN(new_n1021));
  INV_X1    g596(.A(G1971), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1019), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT55), .B1(G166), .B2(new_n993), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n1026));
  NAND3_X1  g601(.A1(G303), .A2(new_n1026), .A3(G8), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1024), .A2(new_n1029), .A3(G8), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n716), .A2(G1976), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT52), .B1(G288), .B2(new_n719), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1003), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1015), .A2(new_n1002), .A3(new_n1016), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1035), .A2(G8), .A3(new_n1032), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT52), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1006), .A2(new_n1034), .A3(new_n1037), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1008), .A2(new_n1003), .B1(new_n1031), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1014), .A2(new_n1017), .A3(new_n1002), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n964), .A2(new_n1020), .A3(new_n1002), .A4(new_n778), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n1040), .A2(new_n749), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT125), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT123), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1041), .B1(new_n1045), .B2(G2078), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1046), .B1(new_n1045), .B2(G2078), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1047), .B1(new_n1010), .B2(KEYINPUT45), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT122), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n964), .A2(new_n1049), .A3(new_n1002), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1049), .B1(new_n964), .B2(new_n1002), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1048), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1043), .A2(new_n1044), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1044), .B1(new_n1043), .B2(new_n1052), .ZN(new_n1054));
  OAI21_X1  g629(.A(G171), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT126), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT45), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT112), .B1(new_n1058), .B2(new_n965), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n963), .B1(new_n999), .B2(new_n1000), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT112), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(new_n1061), .A3(new_n1002), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1041), .A2(G2078), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1059), .A2(new_n1020), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n1043), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT124), .B1(new_n1065), .B2(G171), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT124), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1064), .A2(new_n1043), .A3(new_n1067), .A4(G301), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1057), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT126), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1070), .B(G171), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1056), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1062), .A2(new_n1020), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1061), .B1(new_n1060), .B2(new_n1002), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n831), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1040), .A2(G2084), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1075), .A2(G168), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT51), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1079), .A2(new_n993), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(G168), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT51), .B1(new_n1078), .B2(G8), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT50), .B1(new_n999), .B2(new_n1000), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n965), .B1(new_n1011), .B2(new_n1010), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1088), .A2(new_n1018), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1028), .B1(new_n1089), .B2(new_n993), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1090), .A2(new_n1038), .A3(new_n1030), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1065), .A2(G171), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1043), .A2(G301), .A3(new_n1052), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1091), .B1(new_n1094), .B2(new_n1057), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1072), .A2(new_n1085), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT117), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1035), .A2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1015), .A2(new_n1002), .A3(KEYINPUT117), .A4(new_n1016), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1100), .A2(new_n810), .B1(new_n798), .B2(new_n1040), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1101), .A2(new_n911), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n617), .A2(KEYINPUT57), .A3(new_n566), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1103), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1104));
  AOI21_X1  g679(.A(G1956), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1106), .B(new_n793), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1021), .A2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1104), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1102), .A2(new_n1111), .ZN(new_n1112));
  AND2_X1   g687(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1113));
  OAI22_X1  g688(.A1(new_n1113), .A2(new_n1103), .B1(new_n1105), .B2(new_n1109), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT117), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1099), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n810), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1040), .A2(new_n798), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT60), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT121), .B1(new_n1101), .B2(KEYINPUT60), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1120), .B1(new_n1121), .B2(new_n911), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1118), .A2(KEYINPUT60), .A3(new_n1119), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1101), .A2(KEYINPUT121), .A3(KEYINPUT60), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(new_n1126), .A3(new_n611), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT120), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1129), .B1(new_n1104), .B2(new_n1110), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1128), .B1(new_n1130), .B2(KEYINPUT61), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT61), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1111), .A2(new_n1114), .A3(new_n1129), .A4(new_n1132), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1122), .A2(new_n1127), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  XOR2_X1   g709(.A(KEYINPUT58), .B(G1341), .Z(new_n1135));
  NAND3_X1  g710(.A1(new_n1098), .A2(new_n1099), .A3(new_n1135), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n1021), .A2(G1996), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1136), .A2(KEYINPUT118), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(KEYINPUT118), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n555), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n555), .B(new_n1141), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1115), .B1(new_n1134), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1039), .B1(new_n1096), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT115), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1024), .A2(G8), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n1028), .ZN(new_n1150));
  AOI21_X1  g725(.A(KEYINPUT114), .B1(new_n1150), .B2(new_n1038), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1029), .B1(new_n1024), .B2(G8), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1006), .A2(new_n1034), .A3(new_n1037), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT114), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1157));
  NOR2_X1   g732(.A1(G286), .A2(new_n993), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1157), .A2(KEYINPUT63), .A3(new_n1030), .A4(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1148), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1159), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1161), .B(KEYINPUT115), .C1(new_n1151), .C2(new_n1155), .ZN(new_n1162));
  XOR2_X1   g737(.A(KEYINPUT113), .B(KEYINPUT63), .Z(new_n1163));
  NAND2_X1  g738(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1163), .B1(new_n1091), .B2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1160), .A2(new_n1162), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT62), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1167), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1078), .A2(G8), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n1079), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1170), .B(KEYINPUT62), .C1(new_n1082), .C2(new_n1081), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1168), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1166), .A2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n983), .B1(new_n1147), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT46), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n771), .B1(new_n1176), .B2(G1996), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n966), .B1(new_n1177), .B2(new_n974), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n966), .A2(new_n978), .ZN(new_n1179));
  AOI21_X1  g754(.A(KEYINPUT127), .B1(new_n1179), .B2(new_n1176), .ZN(new_n1180));
  AND3_X1   g755(.A1(new_n1179), .A2(KEYINPUT127), .A3(new_n1176), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1178), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n1182), .B(KEYINPUT47), .Z(new_n1183));
  XNOR2_X1  g758(.A(new_n968), .B(KEYINPUT48), .ZN(new_n1184));
  AND3_X1   g759(.A1(new_n982), .A2(new_n973), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(new_n972), .ZN(new_n1186));
  OAI22_X1  g761(.A1(new_n981), .A2(new_n1186), .B1(G2067), .B2(new_n808), .ZN(new_n1187));
  AOI211_X1 g762(.A(new_n1183), .B(new_n1185), .C1(new_n966), .C2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1175), .A2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g764(.A(new_n458), .ZN(new_n1191));
  OR3_X1    g765(.A1(G401), .A2(G227), .A3(new_n1191), .ZN(new_n1192));
  NOR2_X1   g766(.A1(G229), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g767(.A(new_n1193), .B1(new_n894), .B2(new_n895), .ZN(new_n1194));
  NOR2_X1   g768(.A1(new_n1194), .A2(new_n959), .ZN(G308));
  OR2_X1    g769(.A1(new_n1194), .A2(new_n959), .ZN(G225));
endmodule


