//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 0 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G169gat), .ZN(new_n204));
  INV_X1    g003(.A(G176gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n203), .B1(KEYINPUT26), .B2(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT26), .ZN(new_n209));
  AND3_X1   g008(.A1(new_n208), .A2(KEYINPUT70), .A3(new_n209), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT70), .B1(new_n208), .B2(new_n209), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n207), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT27), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n216), .A2(G183gat), .ZN(new_n217));
  INV_X1    g016(.A(G183gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(KEYINPUT27), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT28), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(G190gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT68), .B1(new_n217), .B2(new_n219), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n218), .A2(KEYINPUT27), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT68), .ZN(new_n226));
  AOI21_X1  g025(.A(G190gat), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT28), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT69), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n223), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n216), .A2(G183gat), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n226), .B1(new_n225), .B2(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n226), .B1(new_n216), .B2(G183gat), .ZN(new_n233));
  INV_X1    g032(.A(G190gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n229), .B(new_n221), .C1(new_n232), .C2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n215), .B1(new_n230), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G120gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G113gat), .ZN(new_n240));
  INV_X1    g039(.A(G113gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G120gat), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT1), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G127gat), .B(G134gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  OR2_X1    g045(.A1(KEYINPUT71), .A2(G127gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT72), .ZN(new_n248));
  NAND2_X1  g047(.A1(KEYINPUT71), .A2(G127gat), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n247), .A2(new_n248), .A3(G134gat), .A4(new_n249), .ZN(new_n250));
  AND2_X1   g049(.A1(KEYINPUT71), .A2(G127gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(KEYINPUT71), .A2(G127gat), .ZN(new_n252));
  INV_X1    g051(.A(G134gat), .ZN(new_n253));
  NOR3_X1   g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G127gat), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT72), .B1(new_n255), .B2(G134gat), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n250), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT73), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n243), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  OAI211_X1 g058(.A(KEYINPUT73), .B(new_n250), .C1(new_n254), .C2(new_n256), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n246), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n262), .B1(G183gat), .B2(G190gat), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n264));
  OAI21_X1  g063(.A(KEYINPUT65), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n264), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n218), .A2(new_n234), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT65), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n266), .A2(new_n267), .A3(new_n268), .A4(new_n262), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n203), .B1(KEYINPUT23), .B2(new_n208), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT23), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n206), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n265), .A2(new_n269), .A3(new_n270), .A4(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT25), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT66), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n208), .A2(KEYINPUT23), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n276), .B1(new_n277), .B2(new_n202), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n272), .A2(KEYINPUT25), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT24), .ZN(new_n281));
  INV_X1    g080(.A(new_n213), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n281), .B1(new_n282), .B2(KEYINPUT67), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT67), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n213), .A2(new_n284), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n267), .B(new_n262), .C1(new_n283), .C2(new_n285), .ZN(new_n286));
  AND3_X1   g085(.A1(new_n277), .A2(new_n276), .A3(new_n202), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n280), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n275), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n238), .A2(new_n261), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT74), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n221), .B1(new_n232), .B2(new_n235), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT69), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n294), .A2(new_n236), .A3(new_n223), .ZN(new_n295));
  AOI22_X1  g094(.A1(new_n295), .A2(new_n215), .B1(new_n275), .B2(new_n289), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n296), .A2(new_n297), .A3(new_n261), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT75), .B1(new_n296), .B2(new_n261), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n257), .A2(new_n258), .ZN(new_n300));
  INV_X1    g099(.A(new_n243), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(new_n301), .A3(new_n260), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(new_n245), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT75), .ZN(new_n304));
  AOI22_X1  g103(.A1(new_n293), .A2(KEYINPUT69), .B1(new_n220), .B2(new_n222), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n214), .B1(new_n305), .B2(new_n236), .ZN(new_n306));
  NOR3_X1   g105(.A1(new_n287), .A2(new_n278), .A3(new_n279), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n307), .A2(new_n286), .B1(new_n273), .B2(new_n274), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n303), .B(new_n304), .C1(new_n306), .C2(new_n308), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n292), .A2(new_n298), .B1(new_n299), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G227gat), .A2(G233gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n311), .B(KEYINPUT64), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT32), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT33), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n315), .B1(new_n310), .B2(new_n313), .ZN(new_n316));
  XOR2_X1   g115(.A(G15gat), .B(G43gat), .Z(new_n317));
  XNOR2_X1  g116(.A(G71gat), .B(G99gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n314), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n319), .ZN(new_n321));
  OAI221_X1 g120(.A(KEYINPUT32), .B1(new_n315), .B2(new_n321), .C1(new_n310), .C2(new_n313), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n292), .A2(new_n298), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n299), .A2(new_n309), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT34), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n324), .A2(new_n325), .A3(new_n326), .A4(new_n313), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT77), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n324), .A2(new_n325), .A3(new_n311), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT76), .B(KEYINPUT34), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n327), .A2(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OR2_X1    g130(.A1(new_n327), .A2(new_n328), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n323), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n320), .A2(new_n322), .A3(new_n332), .A4(new_n331), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n334), .A2(KEYINPUT36), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT36), .ZN(new_n337));
  AND4_X1   g136(.A1(new_n320), .A2(new_n322), .A3(new_n332), .A4(new_n331), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n320), .A2(new_n322), .B1(new_n331), .B2(new_n332), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G1gat), .B(G29gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n341), .B(KEYINPUT0), .ZN(new_n342));
  XNOR2_X1  g141(.A(G57gat), .B(G85gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n342), .B(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT82), .B(G162gat), .ZN(new_n345));
  INV_X1    g144(.A(G155gat), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT2), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OR2_X1    g146(.A1(G141gat), .A2(G148gat), .ZN(new_n348));
  INV_X1    g147(.A(G162gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G155gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n346), .A2(G162gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(G141gat), .A2(G148gat), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n348), .A2(new_n350), .A3(new_n351), .A4(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT2), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n348), .A2(new_n355), .A3(new_n352), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n350), .A2(new_n351), .ZN(new_n357));
  AOI22_X1  g156(.A1(new_n347), .A2(new_n354), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n302), .A2(new_n245), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n356), .A2(new_n357), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT3), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n349), .A2(KEYINPUT82), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT82), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(G162gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n355), .B1(new_n367), .B2(G155gat), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n362), .B(new_n363), .C1(new_n368), .C2(new_n353), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n362), .B1(new_n368), .B2(new_n353), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT3), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n303), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n261), .A2(KEYINPUT4), .A3(new_n358), .ZN(new_n373));
  NAND2_X1  g172(.A1(G225gat), .A2(G233gat), .ZN(new_n374));
  AND4_X1   g173(.A1(new_n361), .A2(new_n372), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n374), .ZN(new_n376));
  AOI211_X1 g175(.A(new_n246), .B(new_n370), .C1(new_n259), .C2(new_n260), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n358), .B1(new_n302), .B2(new_n245), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT5), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT5), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n372), .A2(new_n382), .A3(new_n374), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT83), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n359), .A2(new_n360), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT4), .B1(new_n261), .B2(new_n358), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n361), .A2(new_n373), .A3(KEYINPUT83), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n383), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI211_X1 g188(.A(KEYINPUT6), .B(new_n344), .C1(new_n381), .C2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n344), .B1(new_n381), .B2(new_n389), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n303), .A2(new_n370), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n359), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n382), .B1(new_n393), .B2(new_n376), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n361), .A2(new_n372), .A3(new_n373), .A4(new_n374), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n344), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n383), .ZN(new_n397));
  INV_X1    g196(.A(new_n388), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT83), .B1(new_n361), .B2(new_n373), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT6), .B1(new_n396), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n391), .B1(new_n401), .B2(KEYINPUT84), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT6), .ZN(new_n403));
  INV_X1    g202(.A(new_n344), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n404), .B1(new_n375), .B2(new_n380), .ZN(new_n405));
  OAI211_X1 g204(.A(KEYINPUT84), .B(new_n403), .C1(new_n405), .C2(new_n389), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n390), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT81), .ZN(new_n409));
  XNOR2_X1  g208(.A(G8gat), .B(G36gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(G64gat), .B(G92gat), .ZN(new_n411));
  XOR2_X1   g210(.A(new_n410), .B(new_n411), .Z(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(G226gat), .A2(G233gat), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n415), .B1(new_n306), .B2(new_n308), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT29), .B1(new_n238), .B2(new_n290), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n416), .B1(new_n417), .B2(new_n415), .ZN(new_n418));
  XNOR2_X1  g217(.A(G211gat), .B(G218gat), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT22), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT78), .B(G211gat), .ZN(new_n422));
  INV_X1    g221(.A(G218gat), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n421), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G197gat), .B(G204gat), .ZN(new_n425));
  AOI211_X1 g224(.A(KEYINPUT79), .B(new_n420), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(G211gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT78), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT78), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(G211gat), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n423), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n425), .B1(new_n431), .B2(KEYINPUT22), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT79), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n419), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n426), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n414), .B1(new_n296), .B2(KEYINPUT29), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n432), .A2(new_n433), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n420), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n432), .A2(new_n433), .A3(new_n419), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n437), .A2(new_n441), .A3(new_n416), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n413), .B1(new_n436), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n409), .B1(new_n443), .B2(KEYINPUT30), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n437), .A2(new_n441), .A3(new_n416), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n441), .B1(new_n437), .B2(new_n416), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n412), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT30), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(KEYINPUT81), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n443), .A2(KEYINPUT30), .ZN(new_n450));
  XOR2_X1   g249(.A(new_n412), .B(KEYINPUT80), .Z(new_n451));
  NAND3_X1  g250(.A1(new_n436), .A2(new_n442), .A3(new_n451), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n444), .A2(new_n449), .A3(new_n450), .A4(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n408), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT29), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n439), .A2(new_n456), .A3(new_n440), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n358), .B1(new_n457), .B2(new_n363), .ZN(new_n458));
  NAND2_X1  g257(.A1(G228gat), .A2(G233gat), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT29), .B1(new_n358), .B2(new_n363), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n460), .B1(new_n435), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n459), .B(KEYINPUT85), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n432), .A2(new_n419), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n424), .A2(new_n420), .A3(new_n425), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n456), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n363), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n370), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n369), .A2(new_n456), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n441), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n465), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(G22gat), .B1(new_n463), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(G78gat), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n358), .B1(new_n468), .B2(new_n363), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n439), .A2(new_n440), .B1(new_n456), .B2(new_n369), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n464), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(G22gat), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n478), .B(new_n479), .C1(new_n458), .C2(new_n462), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n474), .A2(new_n475), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n475), .B1(new_n474), .B2(new_n480), .ZN(new_n482));
  XNOR2_X1  g281(.A(KEYINPUT31), .B(G50gat), .ZN(new_n483));
  INV_X1    g282(.A(G106gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n481), .A2(new_n482), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n480), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n459), .B1(new_n441), .B2(new_n471), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT3), .B1(new_n435), .B2(new_n456), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n489), .B1(new_n490), .B2(new_n358), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n479), .B1(new_n491), .B2(new_n478), .ZN(new_n492));
  OAI21_X1  g291(.A(G78gat), .B1(new_n488), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n474), .A2(new_n475), .A3(new_n480), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n485), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n487), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n336), .A2(new_n340), .B1(new_n455), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n403), .B1(new_n405), .B2(new_n389), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n394), .A2(new_n395), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n404), .B1(new_n400), .B2(new_n500), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n390), .B(new_n447), .C1(new_n499), .C2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT37), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(new_n445), .B2(new_n446), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n436), .A2(new_n442), .A3(KEYINPUT37), .ZN(new_n506));
  XOR2_X1   g305(.A(KEYINPUT86), .B(KEYINPUT38), .Z(new_n507));
  AND2_X1   g306(.A1(new_n451), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n505), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT87), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT87), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n505), .A2(new_n506), .A3(new_n511), .A4(new_n508), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n505), .A2(new_n413), .A3(new_n506), .ZN(new_n514));
  INV_X1    g313(.A(new_n507), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n503), .A2(new_n513), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n392), .A2(new_n359), .A3(new_n374), .ZN(new_n518));
  INV_X1    g317(.A(new_n372), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n519), .B1(new_n387), .B2(new_n388), .ZN(new_n520));
  OAI211_X1 g319(.A(KEYINPUT39), .B(new_n518), .C1(new_n520), .C2(new_n374), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n372), .B1(new_n398), .B2(new_n399), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT39), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(new_n523), .A3(new_n376), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n521), .A2(new_n524), .A3(new_n404), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT40), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n521), .A2(new_n524), .A3(KEYINPUT40), .A4(new_n404), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n527), .A2(new_n453), .A3(new_n391), .A4(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n517), .A2(new_n529), .A3(new_n496), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n334), .A2(new_n496), .A3(new_n335), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT35), .B1(new_n455), .B2(new_n531), .ZN(new_n532));
  NOR3_X1   g331(.A1(new_n338), .A2(new_n339), .A3(new_n453), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT35), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n390), .B1(new_n499), .B2(new_n501), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n496), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n498), .A2(new_n530), .B1(new_n532), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G15gat), .B(G22gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(KEYINPUT91), .ZN(new_n540));
  INV_X1    g339(.A(G1gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n541), .A2(KEYINPUT16), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n542), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(G8gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(G50gat), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT15), .B1(new_n547), .B2(G43gat), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n548), .B1(G43gat), .B2(new_n547), .ZN(new_n549));
  XOR2_X1   g348(.A(KEYINPUT89), .B(G36gat), .Z(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(G29gat), .ZN(new_n551));
  NOR2_X1   g350(.A1(G29gat), .A2(G36gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT14), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT88), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n551), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n553), .A2(new_n554), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n549), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n549), .A2(new_n553), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n547), .A2(G43gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n547), .A2(G43gat), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n559), .B1(new_n560), .B2(KEYINPUT90), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n561), .B1(KEYINPUT90), .B2(new_n560), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n558), .B(new_n551), .C1(new_n562), .C2(KEYINPUT15), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n557), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT17), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n564), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT17), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n546), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G229gat), .A2(G233gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n544), .B(G8gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(new_n564), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT18), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n569), .A2(new_n572), .A3(KEYINPUT18), .A4(new_n570), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n546), .A2(new_n567), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n570), .B(KEYINPUT13), .Z(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n575), .A2(new_n576), .A3(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G113gat), .B(G141gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(G197gat), .ZN(new_n583));
  XOR2_X1   g382(.A(KEYINPUT11), .B(G169gat), .Z(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n585), .B(KEYINPUT12), .Z(new_n586));
  NAND2_X1  g385(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n586), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n575), .A2(new_n588), .A3(new_n576), .A4(new_n580), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n538), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G183gat), .B(G211gat), .Z(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G127gat), .B(G155gat), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n595), .B(KEYINPUT96), .Z(new_n596));
  INV_X1    g395(.A(G71gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n597), .A2(new_n475), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n475), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n598), .B1(KEYINPUT92), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT9), .ZN(new_n601));
  XNOR2_X1  g400(.A(G57gat), .B(G64gat), .ZN(new_n602));
  OAI221_X1 g401(.A(new_n600), .B1(KEYINPUT92), .B2(new_n599), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(KEYINPUT93), .ZN(new_n604));
  INV_X1    g403(.A(new_n598), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n605), .B1(new_n599), .B2(new_n601), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT94), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT94), .B1(new_n604), .B2(new_n606), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n603), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n612), .A2(KEYINPUT21), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT95), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n613), .A2(new_n614), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n596), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n617), .ZN(new_n619));
  INV_X1    g418(.A(new_n596), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n619), .A2(new_n620), .A3(new_n615), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n594), .B1(new_n618), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT21), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n546), .B1(new_n624), .B2(new_n611), .ZN(new_n625));
  XOR2_X1   g424(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n626));
  NAND2_X1  g425(.A1(G231gat), .A2(G233gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n625), .B(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n618), .A2(new_n621), .A3(new_n594), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n623), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n629), .ZN(new_n632));
  INV_X1    g431(.A(new_n630), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n632), .B1(new_n633), .B2(new_n622), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT97), .ZN(new_n637));
  XNOR2_X1  g436(.A(G134gat), .B(G162gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G99gat), .B(G106gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT98), .ZN(new_n642));
  NAND2_X1  g441(.A1(G85gat), .A2(G92gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT7), .ZN(new_n644));
  NAND2_X1  g443(.A1(G99gat), .A2(G106gat), .ZN(new_n645));
  INV_X1    g444(.A(G85gat), .ZN(new_n646));
  INV_X1    g445(.A(G92gat), .ZN(new_n647));
  AOI22_X1  g446(.A1(KEYINPUT8), .A2(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n642), .B(new_n649), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n650), .A2(KEYINPUT99), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(KEYINPUT99), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n568), .A2(new_n651), .A3(new_n566), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G190gat), .B(G218gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(KEYINPUT100), .ZN(new_n655));
  NAND3_X1  g454(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n650), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n657), .B1(new_n658), .B2(new_n564), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n654), .A2(KEYINPUT100), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n660), .A2(new_n661), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n640), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n660), .A2(new_n661), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n666), .A2(new_n639), .A3(new_n662), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(G230gat), .ZN(new_n670));
  INV_X1    g469(.A(G233gat), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n607), .B(new_n608), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n673), .A2(new_n603), .A3(new_n658), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n611), .A2(new_n650), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT10), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n611), .A2(new_n650), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(KEYINPUT10), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n672), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n672), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n681), .B1(new_n674), .B2(new_n675), .ZN(new_n682));
  XNOR2_X1  g481(.A(G120gat), .B(G148gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(G176gat), .B(G204gat), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n683), .B(new_n684), .Z(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  OR3_X1    g485(.A1(new_n680), .A2(new_n682), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n686), .B1(new_n680), .B2(new_n682), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n635), .A2(new_n669), .A3(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n592), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(new_n408), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT101), .B(G1gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1324gat));
  INV_X1    g495(.A(new_n693), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n545), .B1(new_n697), .B2(new_n453), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT16), .B(G8gat), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n693), .A2(new_n454), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(KEYINPUT42), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(KEYINPUT42), .B2(new_n700), .ZN(G1325gat));
  NAND2_X1  g501(.A1(new_n340), .A2(new_n336), .ZN(new_n703));
  OAI21_X1  g502(.A(G15gat), .B1(new_n693), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n338), .A2(new_n339), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n706), .A2(G15gat), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n704), .B1(new_n693), .B2(new_n707), .ZN(G1326gat));
  NOR2_X1   g507(.A1(new_n693), .A2(new_n496), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT43), .B(G22gat), .Z(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1327gat));
  NOR2_X1   g510(.A1(new_n635), .A2(new_n689), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(new_n669), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n592), .A2(new_n714), .ZN(new_n715));
  OR3_X1    g514(.A1(new_n715), .A2(G29gat), .A3(new_n408), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n716), .A2(KEYINPUT102), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(KEYINPUT102), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT45), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n665), .A2(KEYINPUT104), .A3(new_n667), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT104), .B1(new_n665), .B2(new_n667), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(KEYINPUT44), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(KEYINPUT105), .B1(new_n538), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(KEYINPUT44), .B1(new_n538), .B2(new_n669), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n532), .A2(new_n537), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n455), .A2(new_n497), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n703), .A2(new_n530), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n732), .A2(new_n733), .A3(new_n725), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n727), .A2(new_n728), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n590), .B(KEYINPUT103), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n713), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(G29gat), .B1(new_n738), .B2(new_n408), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n717), .A2(KEYINPUT45), .A3(new_n718), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n721), .A2(new_n739), .A3(new_n740), .ZN(G1328gat));
  NOR3_X1   g540(.A1(new_n715), .A2(new_n454), .A3(new_n550), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT46), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n550), .B1(new_n738), .B2(new_n454), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(G1329gat));
  OAI21_X1  g544(.A(G43gat), .B1(new_n738), .B2(new_n703), .ZN(new_n746));
  INV_X1    g545(.A(new_n715), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n706), .A2(G43gat), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT47), .ZN(new_n749));
  AOI22_X1  g548(.A1(new_n747), .A2(new_n748), .B1(KEYINPUT106), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n749), .A2(KEYINPUT106), .ZN(new_n752));
  XOR2_X1   g551(.A(new_n751), .B(new_n752), .Z(G1330gat));
  OR2_X1    g552(.A1(new_n715), .A2(KEYINPUT107), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n715), .A2(KEYINPUT107), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n754), .A2(new_n547), .A3(new_n497), .A4(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(G50gat), .B1(new_n738), .B2(new_n496), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g558(.A(KEYINPUT103), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n590), .B(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n635), .A2(new_n669), .A3(new_n689), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n538), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n408), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G57gat), .ZN(G1332gat));
  INV_X1    g565(.A(KEYINPUT49), .ZN(new_n767));
  INV_X1    g566(.A(G64gat), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n763), .B(new_n453), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n769), .B(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(KEYINPUT108), .B(KEYINPUT109), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n771), .B(new_n772), .ZN(G1333gat));
  INV_X1    g572(.A(new_n703), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n597), .B1(new_n763), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n706), .A2(G71gat), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n775), .B1(new_n763), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n497), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g579(.A1(new_n761), .A2(new_n635), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n689), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n732), .A2(new_n668), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n726), .B1(new_n729), .B2(new_n731), .ZN(new_n784));
  AOI22_X1  g583(.A1(new_n783), .A2(KEYINPUT44), .B1(new_n784), .B2(new_n733), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n782), .B1(new_n785), .B2(new_n727), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n786), .A2(new_n764), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n788), .A2(KEYINPUT110), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n761), .A2(new_n635), .A3(new_n789), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n703), .A2(new_n530), .A3(new_n730), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT84), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n499), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n793), .A2(new_n391), .A3(new_n406), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n453), .B1(new_n794), .B2(new_n390), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n705), .A2(new_n795), .A3(new_n496), .ZN(new_n796));
  AOI22_X1  g595(.A1(new_n796), .A2(KEYINPUT35), .B1(new_n533), .B2(new_n536), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n668), .B(new_n790), .C1(new_n791), .C2(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n788), .A2(KEYINPUT110), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n799), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n732), .A2(new_n668), .A3(new_n790), .A4(new_n801), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n764), .A2(new_n646), .A3(new_n689), .ZN(new_n805));
  OAI22_X1  g604(.A1(new_n787), .A2(new_n646), .B1(new_n804), .B2(new_n805), .ZN(G1336gat));
  NAND2_X1  g605(.A1(new_n786), .A2(new_n453), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n454), .A2(new_n690), .A3(G92gat), .ZN(new_n808));
  AOI22_X1  g607(.A1(new_n807), .A2(G92gat), .B1(new_n803), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n809), .B(new_n810), .ZN(G1337gat));
  NAND2_X1  g610(.A1(new_n786), .A2(new_n774), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n706), .A2(G99gat), .A3(new_n690), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n812), .A2(G99gat), .B1(new_n803), .B2(new_n813), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(KEYINPUT111), .ZN(G1338gat));
  INV_X1    g614(.A(new_n782), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n735), .A2(new_n497), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(G106gat), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n496), .A2(new_n690), .A3(G106gat), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n800), .A2(new_n802), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n818), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n484), .B1(new_n786), .B2(new_n497), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT112), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n800), .A2(KEYINPUT112), .A3(new_n802), .A4(new_n820), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI211_X1 g626(.A(KEYINPUT113), .B(KEYINPUT53), .C1(new_n823), .C2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n818), .A2(new_n825), .A3(new_n826), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT113), .B1(new_n830), .B2(KEYINPUT53), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n822), .B1(new_n829), .B2(new_n831), .ZN(G1339gat));
  NOR2_X1   g631(.A1(new_n691), .A2(new_n761), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n677), .A2(new_n679), .A3(new_n672), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT114), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n677), .A2(new_n679), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n681), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT114), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n677), .A2(new_n679), .A3(new_n839), .A4(new_n672), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n836), .A2(new_n838), .A3(KEYINPUT54), .A4(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n685), .B1(new_n680), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n841), .A2(KEYINPUT55), .A3(new_n843), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n844), .A2(new_n687), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n570), .B1(new_n569), .B2(new_n572), .ZN(new_n846));
  OAI22_X1  g645(.A1(new_n846), .A2(KEYINPUT115), .B1(new_n578), .B2(new_n579), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n846), .A2(KEYINPUT115), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n585), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n849), .A2(new_n589), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n841), .A2(new_n843), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT55), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n845), .A2(new_n850), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(new_n724), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n849), .A2(new_n689), .A3(new_n589), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n845), .A2(new_n853), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(new_n736), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n855), .B1(new_n858), .B2(new_n724), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n834), .B1(new_n859), .B2(new_n635), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n860), .A2(new_n764), .A3(new_n496), .A4(new_n533), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(new_n241), .A3(new_n761), .ZN(new_n863));
  INV_X1    g662(.A(new_n855), .ZN(new_n864));
  INV_X1    g663(.A(new_n856), .ZN(new_n865));
  INV_X1    g664(.A(new_n857), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n865), .B1(new_n866), .B2(new_n761), .ZN(new_n867));
  INV_X1    g666(.A(new_n724), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n864), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n635), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n833), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(new_n497), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT116), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n872), .A2(new_n873), .A3(new_n764), .A4(new_n533), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n861), .A2(KEYINPUT116), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n591), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n863), .B1(new_n876), .B2(new_n241), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT117), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n879), .B(new_n863), .C1(new_n876), .C2(new_n241), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(G1340gat));
  AOI21_X1  g680(.A(G120gat), .B1(new_n862), .B2(new_n689), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n874), .A2(new_n875), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n690), .A2(new_n239), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(G1341gat));
  NOR2_X1   g684(.A1(new_n251), .A2(new_n252), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n862), .A2(new_n886), .A3(new_n635), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n870), .B1(new_n874), .B2(new_n875), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n887), .B1(new_n888), .B2(new_n886), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT118), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI211_X1 g690(.A(KEYINPUT118), .B(new_n887), .C1(new_n888), .C2(new_n886), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(G1342gat));
  NAND2_X1  g692(.A1(new_n454), .A2(new_n668), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n706), .A2(G134gat), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n872), .A2(new_n764), .A3(new_n895), .ZN(new_n896));
  XOR2_X1   g695(.A(new_n896), .B(KEYINPUT56), .Z(new_n897));
  AOI21_X1  g696(.A(new_n669), .B1(new_n874), .B2(new_n875), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n253), .B2(new_n898), .ZN(G1343gat));
  NOR3_X1   g698(.A1(new_n774), .A2(new_n408), .A3(new_n453), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT57), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n901), .B1(new_n871), .B2(new_n496), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n496), .A2(new_n901), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n853), .A2(new_n590), .A3(new_n687), .A4(new_n844), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT119), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n856), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n849), .A2(new_n689), .A3(KEYINPUT119), .A4(new_n589), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n904), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n669), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n855), .B1(new_n909), .B2(KEYINPUT120), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n908), .A2(new_n911), .A3(new_n669), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n635), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  OAI211_X1 g712(.A(KEYINPUT121), .B(new_n903), .C1(new_n913), .C2(new_n833), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n902), .A2(new_n914), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n908), .A2(new_n911), .A3(new_n669), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n911), .B1(new_n908), .B2(new_n669), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n916), .A2(new_n917), .A3(new_n855), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n834), .B1(new_n918), .B2(new_n635), .ZN(new_n919));
  AOI21_X1  g718(.A(KEYINPUT121), .B1(new_n919), .B2(new_n903), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n590), .B(new_n900), .C1(new_n915), .C2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(G141gat), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n774), .A2(new_n408), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n860), .A2(new_n454), .A3(new_n497), .A4(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n591), .A2(G141gat), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT122), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT122), .ZN(new_n928));
  INV_X1    g727(.A(new_n926), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n924), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n927), .A2(KEYINPUT58), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n922), .A2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT58), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n761), .B(new_n900), .C1(new_n915), .C2(new_n920), .ZN(new_n934));
  AOI22_X1  g733(.A1(new_n934), .A2(G141gat), .B1(new_n925), .B2(new_n926), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n932), .B1(new_n933), .B2(new_n935), .ZN(G1344gat));
  INV_X1    g735(.A(G148gat), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n937), .A2(KEYINPUT59), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n900), .B1(new_n915), .B2(new_n920), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n939), .B2(new_n690), .ZN(new_n940));
  OAI21_X1  g739(.A(KEYINPUT57), .B1(new_n871), .B2(new_n496), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n854), .A2(new_n669), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n635), .B1(new_n942), .B2(new_n909), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n691), .A2(new_n590), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n901), .B(new_n497), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n900), .A2(new_n689), .ZN(new_n947));
  OAI21_X1  g746(.A(G148gat), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  XOR2_X1   g747(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n940), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n925), .A2(new_n937), .A3(new_n689), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1345gat));
  OAI21_X1  g752(.A(G155gat), .B1(new_n939), .B2(new_n870), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n925), .A2(new_n346), .A3(new_n635), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1346gat));
  OAI21_X1  g755(.A(new_n367), .B1(new_n939), .B2(new_n724), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n894), .A2(new_n367), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n860), .A2(new_n497), .A3(new_n923), .A4(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n959), .ZN(G1347gat));
  NAND2_X1  g759(.A1(new_n408), .A2(new_n453), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n706), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n872), .A2(new_n962), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n963), .A2(new_n204), .A3(new_n591), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n871), .A2(new_n764), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n531), .A2(new_n454), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT124), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n967), .B(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(new_n761), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n964), .B1(new_n970), .B2(new_n204), .ZN(G1348gat));
  NAND3_X1  g770(.A1(new_n969), .A2(new_n205), .A3(new_n689), .ZN(new_n972));
  OAI21_X1  g771(.A(G176gat), .B1(new_n963), .B2(new_n690), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(G1349gat));
  OAI21_X1  g773(.A(G183gat), .B1(new_n963), .B2(new_n870), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n635), .A2(new_n220), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n975), .B1(new_n967), .B2(new_n976), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n977), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g777(.A1(new_n969), .A2(new_n234), .A3(new_n868), .ZN(new_n979));
  OAI21_X1  g778(.A(G190gat), .B1(new_n963), .B2(new_n669), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n980), .A2(KEYINPUT61), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n980), .A2(KEYINPUT61), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(G1351gat));
  NOR2_X1   g782(.A1(new_n774), .A2(new_n961), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n941), .A2(new_n945), .A3(new_n984), .ZN(new_n985));
  INV_X1    g784(.A(G197gat), .ZN(new_n986));
  NOR3_X1   g785(.A1(new_n985), .A2(new_n986), .A3(new_n591), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n703), .A2(new_n453), .A3(new_n497), .ZN(new_n988));
  NOR3_X1   g787(.A1(new_n871), .A2(new_n764), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g788(.A(G197gat), .B1(new_n989), .B2(new_n761), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n987), .A2(new_n990), .ZN(G1352gat));
  INV_X1    g790(.A(G204gat), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n989), .A2(new_n992), .A3(new_n689), .ZN(new_n993));
  XOR2_X1   g792(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n994));
  XNOR2_X1  g793(.A(new_n993), .B(new_n994), .ZN(new_n995));
  OAI21_X1  g794(.A(G204gat), .B1(new_n985), .B2(new_n690), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(G1353gat));
  NAND3_X1  g796(.A1(new_n989), .A2(new_n422), .A3(new_n635), .ZN(new_n998));
  XOR2_X1   g797(.A(new_n998), .B(KEYINPUT126), .Z(new_n999));
  OAI21_X1  g798(.A(G211gat), .B1(new_n985), .B2(new_n870), .ZN(new_n1000));
  OR2_X1    g799(.A1(new_n1000), .A2(KEYINPUT63), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(KEYINPUT63), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n999), .A2(new_n1001), .A3(new_n1002), .ZN(G1354gat));
  INV_X1    g802(.A(KEYINPUT127), .ZN(new_n1004));
  AND2_X1   g803(.A1(new_n985), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g804(.A(new_n668), .B1(new_n985), .B2(new_n1004), .ZN(new_n1006));
  OAI21_X1  g805(.A(G218gat), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n989), .A2(new_n423), .A3(new_n868), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1007), .A2(new_n1008), .ZN(G1355gat));
endmodule


