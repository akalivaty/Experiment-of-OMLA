//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944;
  INV_X1    g000(.A(KEYINPUT83), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  INV_X1    g002(.A(G211gat), .ZN(new_n204));
  INV_X1    g003(.A(G218gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(KEYINPUT22), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n207), .B(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT29), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT3), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  INV_X1    g012(.A(G155gat), .ZN(new_n214));
  INV_X1    g013(.A(G162gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G141gat), .B(G148gat), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n213), .B(new_n216), .C1(new_n217), .C2(KEYINPUT2), .ZN(new_n218));
  INV_X1    g017(.A(G141gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G148gat), .ZN(new_n220));
  INV_X1    g019(.A(G148gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G141gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n220), .A2(new_n222), .A3(KEYINPUT78), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n216), .A2(new_n213), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT78), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(new_n219), .A3(G148gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n223), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  AND3_X1   g026(.A1(new_n213), .A2(KEYINPUT79), .A3(KEYINPUT2), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT79), .B1(new_n213), .B2(KEYINPUT2), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n218), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n202), .B1(new_n212), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n207), .B(new_n208), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n234), .B1(new_n235), .B2(KEYINPUT29), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n236), .A2(KEYINPUT83), .A3(new_n231), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n211), .B1(new_n231), .B2(KEYINPUT3), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n235), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n233), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G228gat), .ZN(new_n241));
  INV_X1    g040(.A(G233gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n231), .A2(KEYINPUT80), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT80), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n218), .B(new_n246), .C1(new_n227), .C2(new_n230), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  OAI221_X1 g047(.A(new_n239), .B1(new_n241), .B2(new_n242), .C1(new_n248), .C2(new_n212), .ZN(new_n249));
  AND3_X1   g048(.A1(new_n244), .A2(G22gat), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(G22gat), .B1(new_n244), .B2(new_n249), .ZN(new_n251));
  XNOR2_X1  g050(.A(G78gat), .B(G106gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT31), .B(G50gat), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n252), .B(new_n253), .Z(new_n254));
  OAI22_X1  g053(.A1(new_n250), .A2(new_n251), .B1(KEYINPUT84), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n244), .A2(new_n249), .ZN(new_n256));
  INV_X1    g055(.A(G22gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n254), .B(KEYINPUT84), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n244), .A2(G22gat), .A3(new_n249), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n255), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT28), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT27), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(G183gat), .ZN(new_n265));
  INV_X1    g064(.A(G183gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT27), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT70), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT70), .B1(new_n266), .B2(KEYINPUT27), .ZN(new_n269));
  INV_X1    g068(.A(G190gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n263), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n266), .A2(KEYINPUT27), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n264), .A2(G183gat), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n265), .A2(new_n267), .A3(KEYINPUT71), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n263), .A2(G190gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n272), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT26), .ZN(new_n281));
  INV_X1    g080(.A(G169gat), .ZN(new_n282));
  INV_X1    g081(.A(G176gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n285));
  AND3_X1   g084(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n284), .B(new_n285), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT72), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n288), .A2(new_n292), .A3(new_n289), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n280), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  AND2_X1   g093(.A1(KEYINPUT68), .A2(KEYINPUT24), .ZN(new_n295));
  NOR2_X1   g094(.A1(KEYINPUT68), .A2(KEYINPUT24), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n289), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n300), .A2(new_n301), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n297), .B(new_n299), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT23), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n305), .B1(new_n286), .B2(new_n287), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT67), .ZN(new_n307));
  NAND2_X1  g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT65), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT67), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n312), .A2(new_n313), .A3(new_n305), .ZN(new_n314));
  AND2_X1   g113(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n315));
  NOR2_X1   g114(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n316));
  OAI22_X1  g115(.A1(new_n315), .A2(new_n316), .B1(G169gat), .B2(G176gat), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n304), .A2(new_n307), .A3(new_n314), .A4(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT25), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n317), .A2(new_n312), .A3(new_n305), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT66), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT66), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n317), .A2(new_n312), .A3(new_n322), .A4(new_n305), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT24), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n289), .B1(new_n298), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT25), .B1(new_n325), .B2(new_n300), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n321), .A2(new_n323), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n294), .A2(new_n319), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G120gat), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT74), .B1(new_n329), .B2(G113gat), .ZN(new_n330));
  OR3_X1    g129(.A1(new_n329), .A2(KEYINPUT74), .A3(G113gat), .ZN(new_n331));
  XOR2_X1   g130(.A(KEYINPUT73), .B(G120gat), .Z(new_n332));
  INV_X1    g131(.A(G113gat), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n330), .B(new_n331), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G127gat), .B(G134gat), .ZN(new_n335));
  OR2_X1    g134(.A1(KEYINPUT75), .A2(KEYINPUT1), .ZN(new_n336));
  NAND2_X1  g135(.A1(KEYINPUT75), .A2(KEYINPUT1), .ZN(new_n337));
  AND3_X1   g136(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G113gat), .B(G120gat), .ZN(new_n339));
  OR2_X1    g138(.A1(new_n339), .A2(KEYINPUT1), .ZN(new_n340));
  INV_X1    g139(.A(new_n335), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n334), .A2(new_n338), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n328), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(G227gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n344), .A2(new_n242), .ZN(new_n345));
  INV_X1    g144(.A(new_n342), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n346), .A2(new_n294), .A3(new_n319), .A4(new_n327), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n343), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT32), .ZN(new_n349));
  XOR2_X1   g148(.A(G15gat), .B(G43gat), .Z(new_n350));
  XNOR2_X1  g149(.A(G71gat), .B(G99gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT33), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n353), .B1(new_n348), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT34), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n343), .A2(new_n347), .ZN(new_n357));
  INV_X1    g156(.A(new_n345), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AOI211_X1 g158(.A(KEYINPUT34), .B(new_n345), .C1(new_n343), .C2(new_n347), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n355), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n355), .A2(new_n359), .A3(new_n360), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n349), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT35), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n359), .A2(new_n360), .ZN(new_n366));
  INV_X1    g165(.A(new_n355), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n349), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(new_n369), .A3(new_n361), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n262), .A2(new_n364), .A3(new_n365), .A4(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G225gat), .A2(G233gat), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n346), .A2(new_n231), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n342), .A2(new_n232), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT5), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n245), .A2(new_n342), .A3(new_n247), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT81), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n379), .A2(new_n380), .A3(KEYINPUT4), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n380), .B1(new_n379), .B2(KEYINPUT4), .ZN(new_n382));
  NOR3_X1   g181(.A1(new_n346), .A2(KEYINPUT4), .A3(new_n231), .ZN(new_n383));
  NOR3_X1   g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n342), .B1(KEYINPUT3), .B2(new_n231), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n232), .A2(new_n234), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n373), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n378), .B1(new_n384), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT5), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT4), .B1(new_n346), .B2(new_n231), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT4), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n245), .A2(new_n342), .A3(new_n393), .A4(new_n247), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n389), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G1gat), .B(G29gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(KEYINPUT0), .ZN(new_n401));
  XNOR2_X1  g200(.A(G57gat), .B(G85gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n399), .A2(KEYINPUT82), .A3(KEYINPUT6), .A4(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n379), .A2(KEYINPUT4), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT81), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n379), .A2(new_n380), .A3(KEYINPUT4), .ZN(new_n407));
  INV_X1    g206(.A(new_n383), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n377), .B1(new_n409), .B2(new_n387), .ZN(new_n410));
  OAI211_X1 g209(.A(KEYINPUT6), .B(new_n403), .C1(new_n410), .C2(new_n397), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT82), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AND2_X1   g212(.A1(new_n404), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n403), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n415), .B1(new_n389), .B2(new_n398), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT6), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n415), .B1(new_n391), .B2(new_n396), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n417), .B1(new_n410), .B2(new_n418), .ZN(new_n419));
  NOR3_X1   g218(.A1(new_n416), .A2(new_n419), .A3(KEYINPUT87), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT87), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n387), .A2(new_n390), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n403), .B1(new_n422), .B2(new_n395), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT6), .B1(new_n389), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n403), .B1(new_n410), .B2(new_n397), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n421), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n371), .B1(new_n414), .B2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G8gat), .B(G36gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(G64gat), .B(G92gat), .ZN(new_n430));
  XOR2_X1   g229(.A(new_n429), .B(new_n430), .Z(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT76), .ZN(new_n433));
  NAND2_X1  g232(.A1(G226gat), .A2(G233gat), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n435), .A2(KEYINPUT29), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n323), .A2(new_n326), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n321), .A2(new_n437), .B1(new_n318), .B2(KEYINPUT25), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n436), .B1(new_n438), .B2(new_n294), .ZN(new_n439));
  AND4_X1   g238(.A1(new_n434), .A2(new_n294), .A3(new_n319), .A4(new_n327), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n433), .B(new_n235), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n328), .B1(KEYINPUT29), .B2(new_n435), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n438), .A2(new_n434), .A3(new_n294), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(new_n210), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n442), .A2(new_n443), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n433), .B1(new_n446), .B2(new_n235), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n432), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n235), .B1(new_n439), .B2(new_n440), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT76), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n450), .A2(new_n441), .A3(new_n444), .A4(new_n431), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n448), .A2(KEYINPUT77), .A3(KEYINPUT30), .A4(new_n451), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n445), .A2(new_n447), .ZN(new_n453));
  XOR2_X1   g252(.A(KEYINPUT77), .B(KEYINPUT30), .Z(new_n454));
  NAND3_X1  g253(.A1(new_n453), .A2(new_n431), .A3(new_n454), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n452), .A2(KEYINPUT85), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT85), .B1(new_n452), .B2(new_n455), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n362), .A2(new_n363), .A3(new_n349), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n369), .B1(new_n368), .B2(new_n361), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n424), .A2(new_n425), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n462), .A2(new_n404), .A3(new_n413), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n452), .A2(new_n455), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n461), .A2(new_n463), .A3(new_n262), .A4(new_n464), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n428), .A2(new_n458), .B1(KEYINPUT35), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT90), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT87), .B1(new_n416), .B2(new_n419), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n424), .A2(new_n421), .A3(new_n425), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n468), .A2(new_n469), .A3(new_n404), .A4(new_n413), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n431), .A2(KEYINPUT38), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n449), .A2(new_n444), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n471), .B1(new_n472), .B2(KEYINPUT37), .ZN(new_n473));
  XOR2_X1   g272(.A(KEYINPUT88), .B(KEYINPUT37), .Z(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n450), .A2(new_n441), .A3(new_n444), .A4(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT89), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n473), .A2(new_n476), .A3(KEYINPUT89), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n451), .A3(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n467), .B1(new_n470), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n451), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n482), .A2(new_n477), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n427), .A2(new_n483), .A3(KEYINPUT90), .A4(new_n414), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT37), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n476), .B(new_n432), .C1(new_n453), .C2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT91), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n486), .A2(new_n487), .A3(KEYINPUT38), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n487), .B1(new_n486), .B2(KEYINPUT38), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n481), .A2(new_n484), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n262), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n456), .A2(new_n457), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n392), .A2(new_n394), .B1(new_n385), .B2(new_n386), .ZN(new_n494));
  OR3_X1    g293(.A1(new_n494), .A2(KEYINPUT39), .A3(new_n372), .ZN(new_n495));
  OR3_X1    g294(.A1(new_n374), .A2(new_n373), .A3(new_n375), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n496), .B(KEYINPUT39), .C1(new_n494), .C2(new_n372), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n495), .A2(new_n497), .A3(KEYINPUT40), .A4(new_n415), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n498), .B(KEYINPUT86), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n495), .A2(new_n415), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT40), .B1(new_n500), .B2(new_n497), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n499), .A2(new_n416), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n492), .B1(new_n493), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n491), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n463), .A2(new_n464), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n492), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT36), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n507), .B1(new_n459), .B2(new_n460), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n364), .A2(KEYINPUT36), .A3(new_n370), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n466), .B1(new_n504), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(G113gat), .B(G141gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G169gat), .B(G197gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(KEYINPUT12), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G43gat), .B(G50gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT15), .ZN(new_n522));
  NAND2_X1  g321(.A1(G29gat), .A2(G36gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT93), .ZN(new_n525));
  OR3_X1    g324(.A1(new_n521), .A2(new_n525), .A3(KEYINPUT15), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n525), .B1(new_n521), .B2(KEYINPUT15), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT14), .ZN(new_n531));
  INV_X1    g330(.A(G29gat), .ZN(new_n532));
  INV_X1    g331(.A(G36gat), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT94), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n531), .A2(new_n532), .A3(new_n533), .A4(KEYINPUT94), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n530), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n538), .A2(KEYINPUT95), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n538), .A2(KEYINPUT95), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n528), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n522), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n534), .A2(new_n529), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(new_n523), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G15gat), .B(G22gat), .ZN(new_n548));
  INV_X1    g347(.A(G1gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT16), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n551), .B1(G1gat), .B2(new_n548), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n552), .B(G8gat), .Z(new_n553));
  NAND2_X1  g352(.A1(new_n547), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n553), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n546), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G229gat), .A2(G233gat), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n558), .B(KEYINPUT97), .Z(new_n559));
  XOR2_X1   g358(.A(new_n559), .B(KEYINPUT13), .Z(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT17), .B1(new_n541), .B2(new_n545), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT96), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n553), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT17), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n566), .B1(new_n553), .B2(new_n564), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(new_n547), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n559), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n562), .B1(new_n569), .B2(KEYINPUT18), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT18), .ZN(new_n571));
  AOI211_X1 g370(.A(new_n571), .B(new_n559), .C1(new_n565), .C2(new_n568), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n520), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n565), .A2(new_n568), .ZN(new_n574));
  INV_X1    g373(.A(new_n559), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n571), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n569), .A2(KEYINPUT18), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n577), .A2(new_n578), .A3(new_n562), .A4(new_n519), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n573), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT98), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n573), .A2(new_n579), .A3(KEYINPUT98), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n513), .A2(new_n585), .ZN(new_n586));
  OR2_X1    g385(.A1(G71gat), .A2(G78gat), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT99), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n588), .A2(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n589));
  AND2_X1   g388(.A1(G57gat), .A2(G64gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(G57gat), .A2(G64gat), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n587), .B(new_n589), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  NOR3_X1   g393(.A1(new_n593), .A2(new_n590), .A3(new_n591), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n589), .A2(new_n587), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT21), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(G127gat), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n553), .B1(new_n599), .B2(new_n598), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(new_n214), .ZN(new_n607));
  XOR2_X1   g406(.A(G183gat), .B(G211gat), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n605), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G85gat), .A2(G92gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT7), .ZN(new_n612));
  NAND2_X1  g411(.A1(G99gat), .A2(G106gat), .ZN(new_n613));
  INV_X1    g412(.A(G85gat), .ZN(new_n614));
  INV_X1    g413(.A(G92gat), .ZN(new_n615));
  AOI22_X1  g414(.A1(KEYINPUT8), .A2(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G99gat), .B(G106gat), .Z(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n618), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n620), .A2(new_n612), .A3(new_n616), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(new_n566), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n546), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n546), .A2(new_n623), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n628));
  XNOR2_X1  g427(.A(G190gat), .B(G218gat), .ZN(new_n629));
  OAI22_X1  g428(.A1(new_n626), .A2(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n628), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(G134gat), .B(G162gat), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n630), .B(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT102), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n619), .A2(new_n594), .A3(new_n597), .A4(new_n621), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT10), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n622), .A2(new_n598), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n642), .A2(KEYINPUT101), .A3(new_n638), .ZN(new_n643));
  OR3_X1    g442(.A1(new_n622), .A2(KEYINPUT101), .A3(new_n598), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n637), .B(new_n641), .C1(new_n645), .C2(KEYINPUT10), .ZN(new_n646));
  NAND2_X1  g445(.A1(G230gat), .A2(G233gat), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT10), .B1(new_n643), .B2(new_n644), .ZN(new_n648));
  OAI21_X1  g447(.A(KEYINPUT102), .B1(new_n648), .B2(new_n640), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n646), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n647), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n645), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G120gat), .B(G148gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(G176gat), .B(G204gat), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n653), .B(new_n654), .Z(new_n655));
  NAND3_X1  g454(.A1(new_n650), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n648), .A2(new_n640), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n652), .B1(new_n657), .B2(new_n651), .ZN(new_n658));
  INV_X1    g457(.A(new_n655), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n610), .A2(new_n636), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n586), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(new_n463), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(new_n549), .ZN(G1324gat));
  INV_X1    g464(.A(KEYINPUT42), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n663), .A2(new_n458), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n666), .B1(new_n668), .B2(G8gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT16), .B(G8gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT103), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n673));
  MUX2_X1   g472(.A(KEYINPUT104), .B(new_n673), .S(new_n671), .Z(new_n674));
  AOI22_X1  g473(.A1(new_n669), .A2(new_n672), .B1(new_n667), .B2(new_n674), .ZN(G1325gat));
  OAI21_X1  g474(.A(G15gat), .B1(new_n663), .B2(new_n510), .ZN(new_n676));
  INV_X1    g475(.A(new_n461), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n677), .A2(G15gat), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n676), .B1(new_n663), .B2(new_n678), .ZN(G1326gat));
  OR3_X1    g478(.A1(new_n663), .A2(KEYINPUT105), .A3(new_n262), .ZN(new_n680));
  OAI21_X1  g479(.A(KEYINPUT105), .B1(new_n663), .B2(new_n262), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT43), .B(G22gat), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n682), .B(new_n683), .Z(G1327gat));
  XNOR2_X1  g483(.A(new_n636), .B(KEYINPUT108), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(KEYINPUT109), .B1(new_n513), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n636), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT44), .B1(new_n513), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT109), .ZN(new_n691));
  INV_X1    g490(.A(new_n687), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n511), .B1(new_n491), .B2(new_n503), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n691), .B(new_n692), .C1(new_n693), .C2(new_n466), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n688), .A2(new_n690), .A3(new_n694), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n573), .A2(new_n579), .A3(KEYINPUT107), .ZN(new_n696));
  AOI21_X1  g495(.A(KEYINPUT107), .B1(new_n573), .B2(new_n579), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n610), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n698), .A2(new_n699), .A3(new_n661), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n463), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n532), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n705));
  INV_X1    g504(.A(new_n661), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n610), .A2(new_n636), .A3(new_n706), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT106), .Z(new_n708));
  NAND4_X1  g507(.A1(new_n586), .A2(new_n532), .A3(new_n702), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT45), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n704), .A2(new_n705), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n710), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT110), .B1(new_n712), .B2(new_n703), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(G1328gat));
  NAND2_X1  g513(.A1(new_n586), .A2(new_n708), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n715), .A2(G36gat), .A3(new_n458), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT46), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n701), .A2(new_n493), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n717), .B1(new_n533), .B2(new_n718), .ZN(G1329gat));
  INV_X1    g518(.A(new_n510), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n701), .A2(G43gat), .A3(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(G43gat), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(new_n715), .B2(new_n677), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g524(.A1(new_n715), .A2(G50gat), .A3(new_n262), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n695), .A2(new_n492), .A3(new_n700), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT112), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(G50gat), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n727), .A2(new_n728), .ZN(new_n731));
  OAI211_X1 g530(.A(KEYINPUT48), .B(new_n726), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n727), .A2(G50gat), .ZN(new_n733));
  AOI21_X1  g532(.A(KEYINPUT48), .B1(new_n733), .B2(new_n726), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT111), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI211_X1 g535(.A(KEYINPUT111), .B(KEYINPUT48), .C1(new_n733), .C2(new_n726), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n732), .B1(new_n736), .B2(new_n737), .ZN(G1331gat));
  INV_X1    g537(.A(new_n698), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n699), .A2(new_n689), .A3(new_n661), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n513), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n702), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n493), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT49), .B(G64gat), .Z(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n744), .B2(new_n746), .ZN(G1333gat));
  NAND2_X1  g546(.A1(new_n741), .A2(new_n720), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n677), .A2(G71gat), .ZN(new_n749));
  AOI22_X1  g548(.A1(new_n748), .A2(G71gat), .B1(new_n741), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g550(.A1(new_n741), .A2(new_n492), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g552(.A1(new_n739), .A2(new_n699), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n636), .B(new_n754), .C1(new_n693), .C2(new_n466), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT51), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n755), .B(new_n756), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n757), .A2(KEYINPUT113), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(KEYINPUT113), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n758), .A2(new_n759), .A3(new_n706), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n760), .A2(new_n614), .A3(new_n702), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n739), .A2(new_n699), .A3(new_n706), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n695), .A2(new_n762), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n763), .A2(new_n702), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n761), .B1(new_n614), .B2(new_n764), .ZN(G1336gat));
  AOI21_X1  g564(.A(new_n615), .B1(new_n763), .B2(new_n493), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n458), .A2(G92gat), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n757), .A2(new_n661), .A3(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OR3_X1    g569(.A1(new_n766), .A2(new_n770), .A3(KEYINPUT52), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT52), .B1(new_n766), .B2(new_n770), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(G1337gat));
  INV_X1    g572(.A(G99gat), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n760), .A2(new_n774), .A3(new_n461), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n763), .A2(new_n720), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n775), .B1(new_n774), .B2(new_n776), .ZN(G1338gat));
  NAND3_X1  g576(.A1(new_n695), .A2(new_n492), .A3(new_n762), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT115), .ZN(new_n779));
  AOI22_X1  g578(.A1(new_n778), .A2(G106gat), .B1(new_n779), .B2(KEYINPUT53), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n262), .A2(G106gat), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n755), .A2(new_n756), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n755), .A2(new_n756), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n661), .B(new_n781), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT116), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n757), .A2(KEYINPUT116), .A3(new_n661), .A4(new_n781), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n778), .A2(new_n779), .A3(G106gat), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n789), .A2(new_n790), .A3(new_n780), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n785), .B1(new_n791), .B2(new_n792), .ZN(G1339gat));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n794), .B(new_n647), .C1(new_n648), .C2(new_n640), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n659), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n794), .B1(new_n657), .B2(new_n651), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n796), .B1(new_n650), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n656), .B1(new_n798), .B2(KEYINPUT55), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  AOI211_X1 g599(.A(new_n800), .B(new_n796), .C1(new_n650), .C2(new_n797), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n802), .B1(new_n696), .B2(new_n697), .ZN(new_n803));
  OAI22_X1  g602(.A1(new_n574), .A2(new_n575), .B1(new_n557), .B2(new_n561), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n518), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n579), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n661), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n685), .B1(new_n803), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n802), .A2(new_n685), .A3(new_n806), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n610), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n662), .A2(new_n698), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n262), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT117), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n813), .A2(new_n816), .A3(new_n262), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n493), .A2(new_n463), .A3(new_n677), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(G113gat), .B1(new_n820), .B2(new_n585), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n463), .B1(new_n811), .B2(new_n812), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n677), .A2(new_n492), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n458), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n739), .A2(new_n333), .ZN(new_n829));
  OAI22_X1  g628(.A1(new_n823), .A2(new_n824), .B1(new_n828), .B2(new_n829), .ZN(G1340gat));
  OAI21_X1  g629(.A(G120gat), .B1(new_n820), .B2(new_n706), .ZN(new_n831));
  OR2_X1    g630(.A1(new_n706), .A2(new_n332), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n831), .B1(new_n828), .B2(new_n832), .ZN(G1341gat));
  INV_X1    g632(.A(G127gat), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n820), .A2(new_n834), .A3(new_n610), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n828), .A2(new_n610), .ZN(new_n836));
  OR2_X1    g635(.A1(new_n836), .A2(KEYINPUT119), .ZN(new_n837));
  AOI21_X1  g636(.A(G127gat), .B1(new_n836), .B2(KEYINPUT119), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n835), .B1(new_n837), .B2(new_n838), .ZN(G1342gat));
  INV_X1    g638(.A(G134gat), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n493), .A2(new_n689), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT120), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n827), .A2(new_n840), .A3(new_n843), .ZN(new_n844));
  XOR2_X1   g643(.A(new_n844), .B(KEYINPUT56), .Z(new_n845));
  OAI21_X1  g644(.A(G134gat), .B1(new_n820), .B2(new_n689), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1343gat));
  AOI22_X1  g646(.A1(new_n584), .A2(new_n802), .B1(new_n661), .B2(new_n806), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n809), .B1(new_n848), .B2(new_n636), .ZN(new_n849));
  AOI22_X1  g648(.A1(new_n849), .A2(new_n610), .B1(new_n662), .B2(new_n698), .ZN(new_n850));
  OAI21_X1  g649(.A(KEYINPUT57), .B1(new_n850), .B2(new_n262), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n813), .A2(new_n852), .A3(new_n492), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n720), .A2(new_n463), .A3(new_n493), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n851), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(G141gat), .B1(new_n855), .B2(new_n585), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n720), .A2(new_n262), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n825), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n859), .A2(new_n219), .A3(new_n458), .A4(new_n584), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n856), .A2(new_n857), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(G141gat), .B1(new_n855), .B2(new_n698), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n862), .A2(new_n860), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n861), .B1(new_n863), .B2(new_n857), .ZN(G1344gat));
  NAND4_X1  g663(.A1(new_n859), .A2(new_n221), .A3(new_n458), .A4(new_n661), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n865), .B(KEYINPUT121), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n854), .A2(new_n661), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n585), .A2(new_n662), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n802), .A2(new_n806), .A3(new_n636), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n870), .B1(new_n848), .B2(new_n636), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n869), .B1(new_n871), .B2(new_n610), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n852), .B1(new_n872), .B2(new_n262), .ZN(new_n873));
  AOI211_X1 g672(.A(new_n852), .B(new_n262), .C1(new_n811), .C2(new_n812), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(new_n874), .B2(KEYINPUT122), .ZN(new_n875));
  AND4_X1   g674(.A1(KEYINPUT122), .A2(new_n813), .A3(KEYINPUT57), .A4(new_n492), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n868), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n867), .B1(new_n877), .B2(G148gat), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n867), .A2(G148gat), .ZN(new_n879));
  INV_X1    g678(.A(new_n855), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(new_n880), .B2(new_n661), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n866), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT123), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n866), .B(KEYINPUT123), .C1(new_n878), .C2(new_n881), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(G1345gat));
  OAI21_X1  g685(.A(G155gat), .B1(new_n855), .B2(new_n610), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n859), .A2(new_n458), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n699), .A2(new_n214), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(G1346gat));
  NAND3_X1  g689(.A1(new_n859), .A2(new_n215), .A3(new_n843), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n880), .A2(new_n685), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(new_n892), .B2(new_n215), .ZN(G1347gat));
  NOR2_X1   g692(.A1(new_n458), .A2(new_n702), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n895), .B1(new_n811), .B2(new_n812), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n826), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(G169gat), .B1(new_n898), .B2(new_n739), .ZN(new_n899));
  AOI211_X1 g698(.A(new_n677), .B(new_n895), .C1(new_n815), .C2(new_n817), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n585), .A2(new_n282), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(G1348gat));
  AOI21_X1  g701(.A(new_n283), .B1(new_n900), .B2(new_n661), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT124), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n897), .A2(G176gat), .A3(new_n706), .ZN(new_n905));
  OR3_X1    g704(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n904), .B1(new_n903), .B2(new_n905), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1349gat));
  AOI21_X1  g707(.A(new_n266), .B1(new_n900), .B2(new_n699), .ZN(new_n909));
  AND2_X1   g708(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n910));
  AND4_X1   g709(.A1(new_n276), .A2(new_n898), .A3(new_n277), .A4(new_n699), .ZN(new_n911));
  OR3_X1    g710(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n910), .B1(new_n909), .B2(new_n911), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(G1350gat));
  NAND3_X1  g713(.A1(new_n898), .A2(new_n270), .A3(new_n685), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n270), .B1(new_n900), .B2(new_n636), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT61), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n915), .B1(new_n918), .B2(new_n919), .ZN(G1351gat));
  OR2_X1    g719(.A1(new_n875), .A2(new_n876), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n895), .A2(new_n720), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(G197gat), .B1(new_n923), .B2(new_n585), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n896), .A2(new_n858), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT126), .ZN(new_n926));
  INV_X1    g725(.A(G197gat), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n926), .A2(new_n927), .A3(new_n739), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n924), .B1(new_n930), .B2(new_n931), .ZN(G1352gat));
  OAI21_X1  g731(.A(G204gat), .B1(new_n923), .B2(new_n706), .ZN(new_n933));
  INV_X1    g732(.A(G204gat), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n925), .A2(new_n934), .A3(new_n661), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT62), .Z(new_n936));
  NAND2_X1  g735(.A1(new_n933), .A2(new_n936), .ZN(G1353gat));
  NAND3_X1  g736(.A1(new_n926), .A2(new_n204), .A3(new_n699), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n921), .A2(new_n699), .A3(new_n922), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n939), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT63), .B1(new_n939), .B2(G211gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n938), .B1(new_n940), .B2(new_n941), .ZN(G1354gat));
  OAI21_X1  g741(.A(G218gat), .B1(new_n923), .B2(new_n689), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n926), .A2(new_n205), .A3(new_n685), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1355gat));
endmodule


