//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1269, new_n1270, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1342, new_n1343, new_n1344;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(new_n206));
  INV_X1    g0006(.A(KEYINPUT67), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G68), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(KEYINPUT67), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G58), .A2(G232), .ZN(new_n217));
  NAND4_X1  g0017(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n206), .B1(new_n213), .B2(new_n218), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT68), .Z(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT69), .Z(new_n222));
  NOR2_X1   g0022(.A1(new_n206), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT0), .Z(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(G50), .ZN(new_n229));
  INV_X1    g0029(.A(KEYINPUT65), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n229), .B1(new_n202), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n231), .B1(new_n230), .B2(new_n202), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT66), .Z(new_n233));
  AOI21_X1  g0033(.A(new_n225), .B1(new_n228), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n220), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n222), .A2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  INV_X1    g0046(.A(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT70), .B(G50), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n248), .B(new_n249), .Z(new_n250));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XOR2_X1   g0051(.A(G107), .B(G116), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  AOI21_X1  g0054(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT71), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  OAI211_X1 g0058(.A(G1), .B(G13), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT71), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AND2_X1   g0061(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G33), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G223), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G1698), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n268), .B1(G222), .B2(G1698), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n262), .B(new_n270), .C1(G77), .C2(new_n266), .ZN(new_n271));
  INV_X1    g0071(.A(G45), .ZN(new_n272));
  AOI21_X1  g0072(.A(G1), .B1(new_n258), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n259), .A2(G274), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G1), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n276), .B1(G41), .B2(G45), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n259), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n275), .B1(G226), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n271), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G169), .ZN(new_n283));
  OAI21_X1  g0083(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT8), .B(G58), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n227), .A2(G33), .ZN(new_n286));
  OR3_X1    g0086(.A1(KEYINPUT72), .A2(G20), .A3(G33), .ZN(new_n287));
  OAI21_X1  g0087(.A(KEYINPUT72), .B1(G20), .B2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G150), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n284), .B1(new_n285), .B2(new_n286), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n226), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n276), .A2(G13), .A3(G20), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(new_n294), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n229), .B1(new_n276), .B2(G20), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n298), .A2(new_n299), .B1(new_n229), .B2(new_n297), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n295), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n281), .A2(G179), .ZN(new_n303));
  NOR3_X1   g0103(.A1(new_n283), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n282), .A2(G190), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT9), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n295), .A2(KEYINPUT9), .A3(new_n300), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n281), .A2(G200), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n305), .A2(new_n307), .A3(new_n308), .A4(new_n309), .ZN(new_n310));
  OR2_X1    g0110(.A1(new_n310), .A2(KEYINPUT10), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(KEYINPUT10), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n304), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n276), .A2(G20), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n298), .A2(G68), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G13), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n316), .A2(G1), .ZN(new_n317));
  AND4_X1   g0117(.A1(KEYINPUT12), .A2(new_n211), .A3(G20), .A4(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(KEYINPUT12), .B1(new_n297), .B2(new_n209), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n290), .A2(new_n229), .ZN(new_n321));
  XOR2_X1   g0121(.A(KEYINPUT67), .B(G68), .Z(new_n322));
  INV_X1    g0122(.A(G77), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n322), .A2(new_n227), .B1(new_n323), .B2(new_n286), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n294), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT11), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n315), .B(new_n320), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n325), .A2(new_n326), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(G226), .A2(G1698), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(new_n238), .B2(G1698), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n266), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(G33), .A2(G97), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT77), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT77), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(G33), .A3(G97), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n262), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n274), .B1(new_n278), .B2(new_n212), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT13), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT13), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n340), .A2(new_n345), .A3(new_n342), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n344), .A2(G179), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G169), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n348), .A2(KEYINPUT78), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n350), .B1(new_n344), .B2(new_n346), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT14), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n347), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n346), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n345), .B1(new_n340), .B2(new_n342), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n349), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n356), .A2(KEYINPUT14), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n330), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(G200), .B1(new_n354), .B2(new_n355), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n344), .A2(G190), .A3(new_n346), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n329), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n298), .A2(G77), .A3(new_n314), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT75), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n298), .A2(KEYINPUT75), .A3(G77), .A4(new_n314), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n297), .A2(new_n323), .ZN(new_n367));
  INV_X1    g0167(.A(new_n294), .ZN(new_n368));
  XNOR2_X1  g0168(.A(KEYINPUT15), .B(G87), .ZN(new_n369));
  OAI22_X1  g0169(.A1(new_n369), .A2(new_n286), .B1(new_n227), .B2(new_n323), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT74), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n285), .B(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n370), .B1(new_n372), .B2(new_n289), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n366), .B(new_n367), .C1(new_n368), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n263), .A2(new_n265), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G107), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n263), .A2(new_n265), .A3(G238), .A4(G1698), .ZN(new_n377));
  INV_X1    g0177(.A(G1698), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(G232), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n376), .B(new_n377), .C1(new_n375), .C2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n262), .ZN(new_n381));
  INV_X1    g0181(.A(G244), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n274), .B1(new_n278), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT73), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n274), .B(KEYINPUT73), .C1(new_n278), .C2(new_n382), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n381), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n374), .B1(G200), .B2(new_n387), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n262), .A2(new_n380), .B1(new_n383), .B2(new_n384), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n389), .A2(G190), .A3(new_n386), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT76), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n387), .B2(G179), .ZN(new_n392));
  INV_X1    g0192(.A(G179), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n389), .A2(KEYINPUT76), .A3(new_n393), .A4(new_n386), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n370), .ZN(new_n396));
  XNOR2_X1  g0196(.A(new_n285), .B(KEYINPUT74), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n396), .B1(new_n397), .B2(new_n290), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n398), .A2(new_n294), .B1(new_n323), .B2(new_n297), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n399), .A2(new_n366), .B1(new_n348), .B2(new_n387), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n388), .A2(new_n390), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n313), .A2(new_n358), .A3(new_n361), .A4(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT83), .ZN(new_n403));
  INV_X1    g0203(.A(new_n285), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n314), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n406), .A2(new_n298), .B1(new_n297), .B2(new_n285), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT79), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n264), .ZN(new_n410));
  NAND2_X1  g0210(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(G33), .A3(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(KEYINPUT80), .B1(new_n264), .B2(G33), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT7), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT80), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n410), .A2(new_n417), .A3(G33), .A4(new_n411), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n415), .A2(new_n416), .A3(new_n227), .A4(new_n418), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n419), .A2(G68), .ZN(new_n420));
  AND2_X1   g0220(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n421));
  NOR2_X1   g0221(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n421), .A2(new_n422), .A3(new_n257), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n227), .B(new_n418), .C1(new_n423), .C2(new_n413), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT7), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT81), .ZN(new_n426));
  OAI21_X1  g0226(.A(G58), .B1(new_n208), .B2(new_n210), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n227), .B1(new_n427), .B2(new_n202), .ZN(new_n428));
  INV_X1    g0228(.A(G159), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n287), .B2(new_n288), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n426), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n430), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n201), .B1(new_n322), .B2(G58), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n432), .B(KEYINPUT81), .C1(new_n433), .C2(new_n227), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n420), .A2(new_n425), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n368), .B1(new_n435), .B2(KEYINPUT16), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT16), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n257), .B1(new_n421), .B2(new_n422), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT82), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT82), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n440), .B(new_n257), .C1(new_n421), .C2(new_n422), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n439), .A2(new_n265), .A3(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n416), .A2(G20), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT7), .B1(new_n375), .B2(new_n227), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n211), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n428), .A2(new_n430), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n437), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n408), .B1(new_n436), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n267), .A2(new_n378), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(G226), .B2(new_n378), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n453), .B1(new_n415), .B2(new_n418), .ZN(new_n454));
  INV_X1    g0254(.A(G87), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n257), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n262), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n275), .B1(G232), .B2(new_n279), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n457), .A2(G179), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n348), .B1(new_n457), .B2(new_n458), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(KEYINPUT18), .B1(new_n451), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n431), .A2(new_n434), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n425), .A2(G68), .A3(new_n419), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(KEYINPUT16), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n294), .ZN(new_n466));
  INV_X1    g0266(.A(new_n443), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n438), .A2(KEYINPUT82), .B1(new_n264), .B2(G33), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n467), .B1(new_n468), .B2(new_n441), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n322), .B1(new_n469), .B2(new_n445), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT16), .B1(new_n470), .B2(new_n448), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n407), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n461), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT18), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n450), .A2(new_n294), .A3(new_n465), .ZN(new_n476));
  INV_X1    g0276(.A(G200), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n477), .B1(new_n457), .B2(new_n458), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n457), .A2(new_n458), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n478), .B1(G190), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n476), .A2(new_n407), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT17), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n476), .A2(KEYINPUT17), .A3(new_n480), .A4(new_n407), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n462), .A2(new_n475), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  OR3_X1    g0285(.A1(new_n402), .A2(new_n403), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n403), .B1(new_n402), .B2(new_n485), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n369), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n490), .A2(new_n296), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n415), .A2(new_n418), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(new_n227), .A3(G68), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT19), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n227), .B1(new_n338), .B2(new_n494), .ZN(new_n495));
  NOR3_X1   g0295(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(G97), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n494), .B1(new_n286), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n493), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n491), .B1(new_n501), .B2(new_n294), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n257), .A2(G1), .ZN(new_n503));
  NOR3_X1   g0303(.A1(new_n297), .A2(new_n294), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G87), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n256), .A2(new_n261), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n382), .A2(G1698), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(G238), .B2(G1698), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n421), .A2(new_n422), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n413), .B1(new_n510), .B2(G33), .ZN(new_n511));
  INV_X1    g0311(.A(new_n418), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(G116), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n257), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n506), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n259), .A2(G274), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n272), .A2(G1), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n521), .A2(G250), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n519), .A2(new_n520), .B1(new_n522), .B2(new_n259), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(G200), .B1(new_n517), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n508), .B1(new_n415), .B2(new_n418), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n262), .B1(new_n526), .B2(new_n515), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n527), .A2(G190), .A3(new_n523), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n502), .A2(new_n505), .A3(new_n525), .A4(new_n528), .ZN(new_n529));
  AOI211_X1 g0329(.A(G20), .B(new_n209), .C1(new_n415), .C2(new_n418), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n335), .A2(new_n337), .ZN(new_n531));
  AOI21_X1  g0331(.A(G20), .B1(new_n531), .B2(KEYINPUT19), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n500), .B1(new_n532), .B2(new_n496), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n294), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n491), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n504), .A2(new_n490), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n527), .A2(new_n523), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n348), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n527), .A2(new_n393), .A3(new_n523), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n537), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n529), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(G107), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n543), .A2(KEYINPUT6), .A3(G97), .ZN(new_n544));
  XOR2_X1   g0344(.A(G97), .B(G107), .Z(new_n545));
  OAI21_X1  g0345(.A(new_n544), .B1(new_n545), .B2(KEYINPUT6), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n546), .A2(G20), .B1(G77), .B2(new_n289), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n445), .B1(new_n442), .B2(new_n443), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n547), .B1(new_n548), .B2(new_n543), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n294), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n296), .A2(G97), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(new_n504), .B2(G97), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g0353(.A(KEYINPUT5), .B(G41), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n520), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n555), .A2(new_n518), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n259), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n556), .B1(new_n558), .B2(G257), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n266), .A2(G250), .A3(G1698), .ZN(new_n560));
  NAND2_X1  g0360(.A1(G33), .A2(G283), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT85), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT4), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n378), .A2(G244), .ZN(new_n564));
  NOR4_X1   g0364(.A1(new_n375), .A2(new_n562), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n564), .A2(new_n563), .ZN(new_n566));
  AOI21_X1  g0366(.A(KEYINPUT85), .B1(new_n266), .B2(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n560), .B(new_n561), .C1(new_n565), .C2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n564), .B1(new_n415), .B2(new_n418), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT84), .ZN(new_n570));
  AOI21_X1  g0370(.A(KEYINPUT4), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n564), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(new_n511), .B2(new_n512), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT84), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n568), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n393), .B(new_n559), .C1(new_n575), .C2(new_n506), .ZN(new_n576));
  INV_X1    g0376(.A(new_n559), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n560), .A2(new_n561), .ZN(new_n578));
  INV_X1    g0378(.A(new_n565), .ZN(new_n579));
  INV_X1    g0379(.A(new_n567), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n570), .B(new_n572), .C1(new_n511), .C2(new_n512), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n563), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n569), .A2(new_n570), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n577), .B1(new_n585), .B2(new_n262), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n553), .B(new_n576), .C1(new_n586), .C2(G169), .ZN(new_n587));
  OAI211_X1 g0387(.A(G190), .B(new_n559), .C1(new_n575), .C2(new_n506), .ZN(new_n588));
  INV_X1    g0388(.A(new_n552), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(new_n549), .B2(new_n294), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n588), .B(new_n590), .C1(new_n586), .C2(new_n477), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n542), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n504), .A2(G107), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT87), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT25), .ZN(new_n595));
  AOI21_X1  g0395(.A(G107), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n297), .A2(new_n596), .B1(KEYINPUT87), .B2(KEYINPUT25), .ZN(new_n597));
  NOR4_X1   g0397(.A1(new_n296), .A2(new_n594), .A3(new_n595), .A4(G107), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n593), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(KEYINPUT22), .A2(G87), .ZN(new_n600));
  AOI211_X1 g0400(.A(G20), .B(new_n600), .C1(new_n415), .C2(new_n418), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n515), .A2(new_n227), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT23), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n227), .B2(G107), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n543), .A2(KEYINPUT23), .A3(G20), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR3_X1   g0406(.A1(new_n375), .A2(G20), .A3(new_n455), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n602), .B(new_n606), .C1(new_n607), .C2(KEYINPUT22), .ZN(new_n608));
  OAI21_X1  g0408(.A(KEYINPUT24), .B1(new_n601), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT24), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n455), .A2(G20), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT22), .B1(new_n266), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n606), .A2(new_n602), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n492), .A2(new_n227), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n610), .B(new_n614), .C1(new_n615), .C2(new_n600), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n609), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n599), .B1(new_n617), .B2(new_n294), .ZN(new_n618));
  OR2_X1    g0418(.A1(G250), .A2(G1698), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(G257), .B2(new_n378), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n620), .B1(new_n415), .B2(new_n418), .ZN(new_n621));
  INV_X1    g0421(.A(G294), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n257), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n262), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n556), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n558), .A2(G264), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n348), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n624), .A2(new_n393), .A3(new_n625), .A4(new_n626), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n618), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n627), .A2(new_n477), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(G190), .B2(new_n627), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n631), .B1(new_n618), .B2(new_n633), .ZN(new_n634));
  OR2_X1    g0434(.A1(G257), .A2(G1698), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(G264), .B2(new_n378), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n636), .B1(new_n415), .B2(new_n418), .ZN(new_n637));
  INV_X1    g0437(.A(G303), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n266), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n262), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n556), .B1(new_n558), .B2(G270), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n297), .A2(KEYINPUT86), .A3(new_n514), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT86), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n644), .B1(new_n296), .B2(G116), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n504), .A2(G116), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n561), .B(new_n227), .C1(G33), .C2(new_n499), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n514), .A2(G20), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(new_n294), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT20), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n647), .A2(KEYINPUT20), .A3(new_n294), .A4(new_n648), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n348), .B1(new_n646), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n642), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT21), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n640), .A2(new_n641), .A3(G179), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n646), .A2(new_n653), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n642), .A2(KEYINPUT21), .A3(new_n654), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n657), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n642), .A2(G200), .ZN(new_n663));
  INV_X1    g0463(.A(new_n659), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n640), .A2(new_n641), .A3(G190), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n634), .A2(new_n667), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n489), .A2(new_n592), .A3(new_n668), .ZN(G372));
  AND2_X1   g0469(.A1(new_n483), .A2(new_n484), .ZN(new_n670));
  INV_X1    g0470(.A(new_n361), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n395), .A2(new_n400), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n671), .B1(new_n358), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  AOI211_X1 g0474(.A(KEYINPUT18), .B(new_n461), .C1(new_n476), .C2(new_n407), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n474), .B1(new_n472), .B2(new_n473), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n310), .B(KEYINPUT10), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n304), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n559), .B1(new_n575), .B2(new_n506), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n590), .B1(new_n681), .B2(new_n348), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n542), .A2(KEYINPUT26), .A3(new_n576), .A4(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT26), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n529), .A2(new_n541), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n684), .B1(new_n587), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n633), .A2(new_n618), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n631), .B2(new_n662), .ZN(new_n689));
  OAI211_X1 g0489(.A(new_n687), .B(new_n541), .C1(new_n592), .C2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n680), .B1(new_n489), .B2(new_n691), .ZN(G369));
  NAND2_X1  g0492(.A1(new_n317), .A2(new_n227), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n694), .A2(G213), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G343), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n634), .B1(new_n618), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n697), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n631), .A2(new_n699), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n698), .A2(KEYINPUT88), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(KEYINPUT88), .B1(new_n698), .B2(new_n700), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n662), .A2(new_n697), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n631), .A2(new_n697), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n703), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n699), .A2(new_n659), .ZN(new_n710));
  MUX2_X1   g0510(.A(new_n662), .B(new_n667), .S(new_n710), .Z(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(G330), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n708), .A2(new_n714), .ZN(G399));
  INV_X1    g0515(.A(new_n223), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G41), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n497), .A2(G116), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(G1), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n232), .B2(new_n718), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT28), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT29), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n690), .A2(new_n723), .A3(new_n697), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n541), .B1(new_n592), .B2(new_n689), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT89), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n683), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n683), .A2(new_n686), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n726), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n699), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n724), .B1(new_n731), .B2(new_n723), .ZN(new_n732));
  INV_X1    g0532(.A(new_n538), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n624), .A2(new_n626), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n658), .A2(new_n733), .A3(KEYINPUT30), .A4(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT30), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n527), .A2(new_n624), .A3(new_n523), .A4(new_n626), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n640), .A2(new_n641), .A3(G179), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n735), .A2(new_n739), .A3(new_n586), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n627), .A2(new_n642), .A3(new_n538), .A4(new_n393), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n681), .A2(new_n741), .A3(KEYINPUT30), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n740), .A2(new_n699), .A3(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT31), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n740), .A2(KEYINPUT31), .A3(new_n742), .A4(new_n699), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n618), .A2(new_n630), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n667), .A2(new_n747), .A3(new_n688), .A4(new_n697), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n745), .B(new_n746), .C1(new_n748), .C2(new_n592), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G330), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n732), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n722), .B1(new_n752), .B2(G1), .ZN(G364));
  INV_X1    g0553(.A(new_n712), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n316), .A2(G20), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G45), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n756), .A2(KEYINPUT90), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(KEYINPUT90), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n757), .A2(G1), .A3(new_n758), .ZN(new_n759));
  OR3_X1    g0559(.A1(new_n717), .A2(KEYINPUT91), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(KEYINPUT91), .B1(new_n717), .B2(new_n759), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n754), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n764), .B1(G330), .B2(new_n711), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n226), .B1(G20), .B2(new_n348), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OR3_X1    g0567(.A1(new_n477), .A2(KEYINPUT96), .A3(G179), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n227), .A2(G190), .ZN(new_n769));
  OAI21_X1  g0569(.A(KEYINPUT96), .B1(new_n477), .B2(G179), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n543), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n393), .A2(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G190), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n227), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n773), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n266), .B1(new_n774), .B2(new_n323), .C1(new_n247), .C2(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n768), .A2(new_n770), .A3(new_n776), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n772), .B(new_n778), .C1(G87), .C2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G179), .A2(G200), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n769), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n429), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT95), .ZN(new_n785));
  XNOR2_X1  g0585(.A(KEYINPUT94), .B(KEYINPUT32), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n785), .A2(new_n787), .ZN(new_n789));
  NAND3_X1  g0589(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(G190), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n227), .B1(new_n782), .B2(G190), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n792), .A2(new_n209), .B1(new_n793), .B2(new_n499), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n790), .A2(new_n775), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n794), .B1(G50), .B2(new_n795), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n781), .A2(new_n788), .A3(new_n789), .A4(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n793), .A2(new_n622), .ZN(new_n798));
  OR2_X1    g0598(.A1(KEYINPUT33), .A2(G317), .ZN(new_n799));
  NAND2_X1  g0599(.A1(KEYINPUT33), .A2(G317), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n792), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n798), .B(new_n801), .C1(G326), .C2(new_n795), .ZN(new_n802));
  INV_X1    g0602(.A(new_n771), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G283), .ZN(new_n804));
  INV_X1    g0604(.A(G311), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n774), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G322), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n375), .B1(new_n777), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n783), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n806), .B(new_n808), .C1(G329), .C2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n780), .A2(G303), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n802), .A2(new_n804), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n767), .B1(new_n797), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(G13), .A2(G33), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(G20), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n766), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n716), .A2(new_n492), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(new_n233), .B2(new_n272), .ZN(new_n820));
  INV_X1    g0620(.A(new_n250), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n820), .B1(new_n821), .B2(new_n272), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n223), .A2(new_n266), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT92), .ZN(new_n824));
  XOR2_X1   g0624(.A(G355), .B(KEYINPUT93), .Z(new_n825));
  AOI22_X1  g0625(.A1(new_n824), .A2(new_n825), .B1(new_n514), .B2(new_n716), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n762), .B(new_n813), .C1(new_n817), .C2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n816), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n828), .B1(new_n711), .B2(new_n829), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n765), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(G396));
  AOI21_X1  g0632(.A(new_n697), .B1(new_n399), .B2(new_n366), .ZN(new_n833));
  AND3_X1   g0633(.A1(new_n395), .A2(new_n400), .A3(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n833), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n834), .B1(new_n401), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(new_n690), .B2(new_n697), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT99), .Z(new_n839));
  AND2_X1   g0639(.A1(new_n401), .A2(new_n697), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n839), .B1(new_n690), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n841), .A2(new_n751), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n842), .A2(new_n763), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n841), .A2(new_n751), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n774), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n846), .A2(G116), .B1(G283), .B2(new_n791), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT97), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n375), .B1(new_n783), .B2(new_n805), .C1(new_n622), .C2(new_n777), .ZN(new_n849));
  INV_X1    g0649(.A(new_n795), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n850), .A2(new_n638), .B1(new_n793), .B2(new_n499), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n543), .A2(new_n779), .B1(new_n771), .B2(new_n455), .ZN(new_n852));
  NOR4_X1   g0652(.A1(new_n848), .A2(new_n849), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT98), .ZN(new_n855));
  INV_X1    g0655(.A(new_n777), .ZN(new_n856));
  AOI22_X1  g0656(.A1(G143), .A2(new_n856), .B1(new_n846), .B2(G159), .ZN(new_n857));
  INV_X1    g0657(.A(G137), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n857), .B1(new_n850), .B2(new_n858), .C1(new_n291), .C2(new_n792), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT34), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n859), .A2(new_n860), .ZN(new_n862));
  INV_X1    g0662(.A(new_n793), .ZN(new_n863));
  AOI22_X1  g0663(.A1(G132), .A2(new_n809), .B1(new_n863), .B2(G58), .ZN(new_n864));
  AOI22_X1  g0664(.A1(G50), .A2(new_n780), .B1(new_n803), .B2(G68), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n862), .A2(new_n492), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n855), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n854), .A2(KEYINPUT98), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n766), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n766), .A2(new_n814), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n762), .B1(new_n323), .B2(new_n870), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n869), .B(new_n871), .C1(new_n837), .C2(new_n815), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n845), .A2(new_n872), .ZN(G384));
  AOI21_X1  g0673(.A(KEYINPUT16), .B1(new_n463), .B2(new_n464), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n407), .B1(new_n466), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n473), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n696), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(new_n877), .A3(new_n481), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT37), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n472), .A2(new_n473), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n472), .A2(new_n696), .ZN(new_n881));
  XNOR2_X1  g0681(.A(KEYINPUT100), .B(KEYINPUT37), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n880), .A2(new_n881), .A3(new_n481), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n877), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n485), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n884), .A2(new_n886), .A3(KEYINPUT38), .ZN(new_n887));
  INV_X1    g0687(.A(new_n882), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n481), .B1(new_n451), .B2(new_n461), .ZN(new_n889));
  INV_X1    g0689(.A(new_n696), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n451), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n888), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n883), .A2(new_n892), .B1(new_n485), .B2(new_n891), .ZN(new_n893));
  XOR2_X1   g0693(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n887), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n330), .A2(new_n699), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n358), .A2(new_n361), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n356), .A2(KEYINPUT14), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n351), .A2(new_n352), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n899), .A2(new_n900), .A3(new_n347), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n330), .B(new_n699), .C1(new_n901), .C2(new_n671), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n836), .B1(new_n898), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n749), .A2(new_n903), .A3(KEYINPUT40), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n896), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT102), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT102), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n896), .A2(new_n908), .A3(new_n905), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n749), .A2(new_n903), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n884), .A2(new_n886), .A3(KEYINPUT38), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT38), .B1(new_n884), .B2(new_n886), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT40), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n910), .A2(new_n917), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n488), .A2(new_n749), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n918), .A2(new_n919), .ZN(new_n921));
  INV_X1    g0721(.A(G330), .ZN(new_n922));
  NOR3_X1   g0722(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT39), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n913), .A2(new_n914), .A3(new_n924), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n892), .A2(new_n883), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n881), .B1(new_n670), .B2(new_n677), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n894), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT39), .B1(new_n928), .B2(new_n887), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n901), .A2(new_n330), .A3(new_n697), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n677), .A2(new_n696), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n913), .A2(new_n914), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n898), .A2(new_n902), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n840), .B1(new_n729), .B2(new_n725), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n672), .A2(new_n699), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n936), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n933), .B1(new_n934), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n932), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n680), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n732), .B2(new_n488), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n942), .B(new_n944), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n923), .A2(new_n945), .B1(new_n276), .B2(new_n755), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n945), .B2(new_n923), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n546), .A2(KEYINPUT35), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n546), .A2(KEYINPUT35), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n948), .A2(G116), .A3(new_n228), .A4(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT36), .Z(new_n951));
  INV_X1    g0751(.A(new_n232), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n952), .A2(G77), .A3(new_n427), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n229), .A2(G68), .ZN(new_n954));
  AOI211_X1 g0754(.A(new_n276), .B(G13), .C1(new_n953), .C2(new_n954), .ZN(new_n955));
  OR3_X1    g0755(.A1(new_n947), .A2(new_n951), .A3(new_n955), .ZN(G367));
  OAI221_X1 g0756(.A(new_n817), .B1(new_n223), .B2(new_n369), .C1(new_n819), .C2(new_n244), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n763), .A2(new_n957), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n777), .A2(new_n291), .B1(new_n774), .B2(new_n229), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n375), .B(new_n959), .C1(G137), .C2(new_n809), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n793), .A2(new_n209), .ZN(new_n961));
  INV_X1    g0761(.A(G143), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n850), .A2(new_n962), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n961), .B(new_n963), .C1(G159), .C2(new_n791), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n780), .A2(G58), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n803), .A2(G77), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n960), .A2(new_n964), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n779), .A2(new_n514), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT46), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n850), .A2(new_n805), .B1(new_n793), .B2(new_n543), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(G294), .B2(new_n791), .ZN(new_n971));
  INV_X1    g0771(.A(G317), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n777), .A2(new_n638), .B1(new_n783), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(G283), .B2(new_n846), .ZN(new_n974));
  INV_X1    g0774(.A(new_n492), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n771), .A2(new_n499), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n971), .A2(new_n974), .A3(new_n975), .A4(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n967), .B1(new_n969), .B2(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT47), .Z(new_n980));
  NAND2_X1  g0780(.A1(new_n502), .A2(new_n505), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n699), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n542), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n541), .B2(new_n982), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n958), .B1(new_n980), .B2(new_n767), .C1(new_n984), .C2(new_n829), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT44), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n587), .B(new_n591), .C1(new_n590), .C2(new_n697), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n682), .A2(new_n576), .A3(new_n699), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n986), .B1(new_n708), .B2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n989), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n707), .A2(KEYINPUT44), .A3(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n705), .A2(new_n706), .A3(new_n989), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT45), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n993), .A2(new_n994), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n990), .A2(new_n992), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n714), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n703), .B(new_n704), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(new_n754), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n752), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n714), .A2(KEYINPUT104), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n998), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  NOR3_X1   g0804(.A1(new_n997), .A2(KEYINPUT104), .A3(new_n714), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n752), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n717), .B(KEYINPUT41), .Z(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n759), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n987), .A2(new_n747), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n699), .B1(new_n1010), .B2(new_n587), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n703), .A2(new_n704), .A3(new_n989), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1013), .A2(KEYINPUT42), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(KEYINPUT42), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1011), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n984), .A2(KEYINPUT103), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n984), .A2(KEYINPUT103), .ZN(new_n1019));
  NOR3_X1   g0819(.A1(new_n1018), .A2(new_n1019), .A3(KEYINPUT43), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1021), .B1(new_n1016), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n713), .A2(new_n989), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1024), .B(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n985), .B1(new_n1009), .B2(new_n1026), .ZN(G387));
  NAND2_X1  g0827(.A1(new_n1000), .A2(new_n759), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n492), .B1(G326), .B2(new_n809), .ZN(new_n1029));
  INV_X1    g0829(.A(G283), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n779), .A2(new_n622), .B1(new_n1030), .B2(new_n793), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G317), .A2(new_n856), .B1(new_n846), .B2(G303), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n850), .B2(new_n807), .C1(new_n805), .C2(new_n792), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT48), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1031), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n1034), .B2(new_n1033), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT49), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1029), .B1(new_n514), .B2(new_n771), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  AND2_X1   g0838(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n780), .A2(G77), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n977), .A2(new_n492), .A3(new_n1040), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G68), .A2(new_n846), .B1(new_n809), .B2(G150), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n850), .B2(new_n429), .C1(new_n285), .C2(new_n792), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT105), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n777), .A2(new_n229), .B1(new_n793), .B2(new_n369), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n1038), .A2(new_n1039), .B1(new_n1041), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n766), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n241), .A2(new_n272), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n719), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1050), .A2(new_n818), .B1(new_n824), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n397), .A2(G50), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT50), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n719), .B(new_n1053), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n1055), .B2(new_n1054), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n1052), .A2(new_n1057), .B1(G107), .B2(new_n223), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n762), .B1(new_n1058), .B2(new_n817), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1049), .B(new_n1059), .C1(new_n703), .C2(new_n829), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1001), .A2(new_n717), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1000), .A2(new_n752), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1028), .B(new_n1060), .C1(new_n1061), .C2(new_n1062), .ZN(G393));
  NAND2_X1  g0863(.A1(new_n818), .A2(new_n253), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1064), .B(new_n817), .C1(new_n499), .C2(new_n223), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n763), .A2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT106), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n779), .A2(new_n211), .B1(new_n962), .B2(new_n783), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT107), .Z(new_n1069));
  NOR2_X1   g0869(.A1(new_n793), .A2(new_n323), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1070), .B(new_n975), .C1(G50), .C2(new_n791), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n850), .A2(new_n291), .B1(new_n777), .B2(new_n429), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT51), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n372), .A2(new_n846), .B1(new_n803), .B2(G87), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1069), .A2(new_n1071), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n850), .A2(new_n972), .B1(new_n777), .B2(new_n805), .ZN(new_n1076));
  XOR2_X1   g0876(.A(KEYINPUT108), .B(KEYINPUT52), .Z(new_n1077));
  XNOR2_X1  g0877(.A(new_n1076), .B(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n375), .B1(new_n774), .B2(new_n622), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(G322), .B2(new_n809), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n863), .A2(G116), .B1(G303), .B2(new_n791), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n772), .B1(G283), .B2(new_n780), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1078), .A2(new_n1080), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1075), .A2(new_n1083), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1067), .B1(new_n767), .B2(new_n1084), .C1(new_n989), .C2(new_n829), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n997), .B(new_n714), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n759), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1086), .ZN(new_n1089));
  OAI21_X1  g0889(.A(KEYINPUT109), .B1(new_n1089), .B2(new_n1002), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT109), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1086), .A2(new_n1091), .A3(new_n1001), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1004), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1005), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n718), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1088), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(G390));
  NAND2_X1  g0898(.A1(new_n488), .A2(new_n751), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n944), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n938), .B1(new_n690), .B2(new_n840), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n936), .B1(new_n750), .B2(new_n836), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n749), .A2(G330), .A3(new_n837), .A4(new_n935), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n938), .B1(new_n731), .B2(new_n837), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1104), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1100), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n931), .ZN(new_n1110));
  OAI21_X1  g0910(.A(KEYINPUT110), .B1(new_n940), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT110), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1112), .B(new_n931), .C1(new_n1101), .C2(new_n936), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1111), .B(new_n1113), .C1(new_n925), .C2(new_n929), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n931), .B(new_n896), .C1(new_n1105), .C2(new_n936), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1114), .A2(new_n1103), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1103), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1109), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1103), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n944), .A2(new_n1099), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1123), .A2(new_n1107), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1122), .A2(new_n1116), .A3(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1119), .A2(new_n1125), .A3(new_n717), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n930), .A2(new_n814), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n774), .A2(new_n499), .B1(new_n783), .B2(new_n622), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n266), .B(new_n1128), .C1(G116), .C2(new_n856), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n850), .A2(new_n1030), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1070), .B(new_n1130), .C1(G107), .C2(new_n791), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n780), .A2(G87), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n803), .A2(G68), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1129), .A2(new_n1131), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n792), .A2(new_n858), .B1(new_n793), .B2(new_n429), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G128), .B2(new_n795), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n803), .A2(G50), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT54), .B(G143), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n375), .B1(new_n846), .B2(new_n1139), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(G132), .A2(new_n856), .B1(new_n809), .B2(G125), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1136), .A2(new_n1137), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n780), .A2(G150), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT53), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1134), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT112), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n767), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n1146), .B2(new_n1145), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n870), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1148), .B(new_n763), .C1(new_n404), .C2(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT113), .ZN(new_n1151));
  OR2_X1    g0951(.A1(new_n1127), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT111), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1153), .B1(new_n1154), .B2(new_n759), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1122), .A2(new_n759), .A3(new_n1116), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1156), .A2(KEYINPUT111), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1126), .B(new_n1152), .C1(new_n1155), .C2(new_n1157), .ZN(G378));
  INV_X1    g0958(.A(KEYINPUT57), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n1125), .B2(new_n1100), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT116), .ZN(new_n1161));
  AOI211_X1 g0961(.A(KEYINPUT102), .B(new_n904), .C1(new_n928), .C2(new_n887), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n908), .B1(new_n896), .B2(new_n905), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n917), .A2(G330), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1161), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n922), .B1(new_n915), .B2(new_n916), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1167), .B(KEYINPUT116), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1168));
  XOR2_X1   g0968(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n302), .A2(new_n890), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n313), .A2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n313), .A2(new_n1172), .ZN(new_n1174));
  OAI21_X1  g0974(.A(KEYINPUT115), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NOR3_X1   g0976(.A1(new_n1173), .A2(new_n1174), .A3(KEYINPUT115), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1170), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1177), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1179), .A2(new_n1169), .A3(new_n1175), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1166), .A2(new_n1168), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1181), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1183), .B(new_n1161), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1182), .A2(new_n942), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n942), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1160), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n717), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n932), .A2(new_n941), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1168), .A2(new_n1181), .ZN(new_n1190));
  AOI21_X1  g0990(.A(KEYINPUT116), .B1(new_n910), .B2(new_n1167), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1184), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1189), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT117), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1182), .A2(new_n942), .A3(new_n1184), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1125), .A2(new_n1100), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1182), .A2(new_n942), .A3(KEYINPUT117), .A4(new_n1184), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1188), .B1(new_n1159), .B2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1197), .A2(new_n759), .A3(new_n1199), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1181), .A2(new_n814), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n777), .A2(new_n543), .B1(new_n783), .B2(new_n1030), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n961), .B(new_n1204), .C1(G116), .C2(new_n795), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n492), .A2(G41), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n803), .A2(G58), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1205), .A2(new_n1040), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n846), .A2(new_n490), .B1(G97), .B2(new_n791), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT114), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n780), .A2(new_n1139), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G128), .A2(new_n856), .B1(new_n846), .B2(G137), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n791), .A2(G132), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n863), .A2(G150), .B1(G125), .B2(new_n795), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n1216), .A2(KEYINPUT59), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(KEYINPUT59), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n803), .A2(G159), .ZN(new_n1219));
  AOI211_X1 g1019(.A(G33), .B(G41), .C1(new_n809), .C2(G124), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1211), .A2(KEYINPUT58), .B1(new_n1217), .B2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1222), .B1(KEYINPUT58), .B2(new_n1211), .C1(new_n1206), .C2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n766), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n870), .A2(new_n229), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1203), .A2(new_n763), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1202), .A2(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1201), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(G375));
  NAND2_X1  g1030(.A1(new_n1123), .A2(new_n1107), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1109), .A2(new_n1008), .A3(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n936), .A2(new_n814), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n763), .B1(G68), .B2(new_n1149), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n266), .B1(new_n809), .B2(G303), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n966), .B(new_n1235), .C1(new_n622), .C2(new_n850), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n792), .A2(new_n514), .B1(new_n774), .B2(new_n543), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT118), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n856), .A2(G283), .B1(new_n863), .B2(new_n490), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1239), .B1(KEYINPUT119), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(KEYINPUT119), .C2(new_n1240), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n1236), .B(new_n1243), .C1(G97), .C2(new_n780), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT120), .ZN(new_n1245));
  OR2_X1    g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n795), .A2(G132), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n1248), .B1(new_n793), .B2(new_n229), .C1(new_n792), .C2(new_n1138), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(G159), .A2(new_n780), .B1(new_n803), .B2(G58), .ZN(new_n1250));
  INV_X1    g1050(.A(G128), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n777), .A2(new_n858), .B1(new_n783), .B2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(G150), .B2(new_n846), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1250), .A2(new_n492), .A3(new_n1253), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1246), .B(new_n1247), .C1(new_n1249), .C2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1234), .B1(new_n1255), .B2(new_n766), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1108), .A2(new_n759), .B1(new_n1233), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1232), .A2(new_n1257), .ZN(G381));
  OR3_X1    g1058(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1259));
  NOR4_X1   g1059(.A1(G390), .A2(G387), .A3(G381), .A4(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(G378), .A2(KEYINPUT121), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1156), .B(KEYINPUT111), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT121), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1262), .A2(new_n1263), .A3(new_n1126), .A4(new_n1152), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1261), .A2(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(G375), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1260), .A2(new_n1266), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(KEYINPUT122), .ZN(G407));
  INV_X1    g1068(.A(new_n1265), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1229), .A2(new_n1269), .ZN(new_n1270));
  OAI211_X1 g1070(.A(G407), .B(G213), .C1(G343), .C2(new_n1270), .ZN(G409));
  XNOR2_X1  g1071(.A(G393), .B(new_n831), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1097), .A2(G387), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1097), .A2(G387), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1273), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  OR2_X1    g1077(.A1(new_n1097), .A2(G387), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1278), .A2(new_n1272), .A3(new_n1274), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1277), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1231), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n718), .B1(new_n1281), .B2(KEYINPUT60), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n1123), .B2(new_n1107), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT124), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1284), .A2(new_n1285), .A3(new_n1231), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1285), .B1(new_n1284), .B2(new_n1231), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1282), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(KEYINPUT125), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT125), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1282), .B(new_n1290), .C1(new_n1286), .C2(new_n1287), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1292), .A2(G384), .A3(new_n1257), .ZN(new_n1293));
  AOI21_X1  g1093(.A(G384), .B1(new_n1292), .B2(new_n1257), .ZN(new_n1294));
  OR2_X1    g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(G213), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1296), .A2(G343), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(G2897), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(new_n1295), .B(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1200), .A2(new_n1159), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1188), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1228), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1302), .A2(G378), .A3(new_n1303), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1197), .A2(new_n1008), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1227), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1306), .B1(new_n1307), .B2(new_n759), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1305), .A2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1269), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1304), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1297), .ZN(new_n1312));
  AOI21_X1  g1112(.A(KEYINPUT126), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT126), .ZN(new_n1314));
  AOI211_X1 g1114(.A(new_n1314), .B(new_n1297), .C1(new_n1304), .C2(new_n1310), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1299), .B1(new_n1313), .B2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(G378), .ZN(new_n1317));
  NOR3_X1   g1117(.A1(new_n1201), .A2(new_n1317), .A3(new_n1228), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1265), .B1(new_n1305), .B2(new_n1308), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1312), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1314), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1311), .A2(KEYINPUT126), .A3(new_n1312), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT127), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT62), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1295), .A2(new_n1324), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1321), .A2(new_n1322), .A3(new_n1323), .A4(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT61), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1316), .A2(new_n1326), .A3(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1321), .A2(new_n1322), .A3(new_n1325), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1311), .A2(new_n1312), .A3(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1323), .B1(new_n1331), .B2(new_n1324), .ZN(new_n1332));
  AND2_X1   g1132(.A1(new_n1329), .A2(new_n1332), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1280), .B1(new_n1328), .B2(new_n1333), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1280), .A2(KEYINPUT61), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1321), .A2(KEYINPUT63), .A3(new_n1322), .A4(new_n1330), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT63), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1331), .A2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1299), .A2(new_n1320), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1335), .A2(new_n1336), .A3(new_n1338), .A4(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1334), .A2(new_n1340), .ZN(G405));
  NAND2_X1  g1141(.A1(G375), .A2(new_n1269), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(new_n1304), .ZN(new_n1343));
  XNOR2_X1  g1143(.A(new_n1343), .B(new_n1330), .ZN(new_n1344));
  XNOR2_X1  g1144(.A(new_n1344), .B(new_n1280), .ZN(G402));
endmodule


