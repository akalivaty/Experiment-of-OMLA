//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 0 1 0 0 1 1 1 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 1 1 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003;
  INV_X1    g000(.A(G64gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(G57gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(G57gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT9), .ZN(new_n205));
  NAND2_X1  g004(.A1(G71gat), .A2(G78gat), .ZN(new_n206));
  AOI22_X1  g005(.A1(new_n203), .A2(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G71gat), .ZN(new_n208));
  INV_X1    g007(.A(G78gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AND3_X1   g009(.A1(new_n207), .A2(new_n206), .A3(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT89), .B1(new_n208), .B2(new_n209), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(KEYINPUT90), .A2(G71gat), .A3(G78gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT90), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n206), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n213), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n214), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(new_n212), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n207), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n211), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT21), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n223), .B(KEYINPUT91), .ZN(new_n224));
  XNOR2_X1  g023(.A(G127gat), .B(G155gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n225), .B(KEYINPUT20), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n224), .B(new_n226), .ZN(new_n227));
  XOR2_X1   g026(.A(G183gat), .B(G211gat), .Z(new_n228));
  XNOR2_X1  g027(.A(new_n228), .B(KEYINPUT93), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G15gat), .B(G22gat), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n231), .A2(G1gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT86), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT16), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n231), .B1(new_n234), .B2(G1gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n232), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G8gat), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n236), .A2(G8gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(new_n222), .B2(new_n221), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n242));
  NAND2_X1  g041(.A1(G231gat), .A2(G233gat), .ZN(new_n243));
  XOR2_X1   g042(.A(new_n242), .B(new_n243), .Z(new_n244));
  XNOR2_X1  g043(.A(new_n241), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n229), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n230), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n245), .B1(new_n230), .B2(new_n246), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(G232gat), .A2(G233gat), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n251), .A2(KEYINPUT41), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT94), .ZN(new_n253));
  XNOR2_X1  g052(.A(G190gat), .B(G218gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n251), .A2(KEYINPUT41), .ZN(new_n257));
  NOR2_X1   g056(.A1(G29gat), .A2(G36gat), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT14), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G29gat), .A2(G36gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT84), .ZN(new_n262));
  XNOR2_X1  g061(.A(G43gat), .B(G50gat), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n260), .A2(KEYINPUT15), .A3(new_n262), .A4(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n260), .A2(KEYINPUT15), .A3(new_n262), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(new_n263), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT15), .B1(new_n260), .B2(new_n262), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n265), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT85), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI211_X1 g070(.A(KEYINPUT85), .B(new_n265), .C1(new_n267), .C2(new_n268), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G99gat), .A2(G106gat), .ZN(new_n274));
  INV_X1    g073(.A(G85gat), .ZN(new_n275));
  INV_X1    g074(.A(G92gat), .ZN(new_n276));
  AOI22_X1  g075(.A1(KEYINPUT8), .A2(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT7), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(new_n275), .B2(new_n276), .ZN(new_n279));
  NAND3_X1  g078(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G99gat), .B(G106gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n277), .A2(new_n282), .A3(new_n279), .A4(new_n280), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n284), .A2(KEYINPUT95), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT95), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n281), .A2(new_n287), .A3(new_n283), .ZN(new_n288));
  AND2_X1   g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n257), .B1(new_n273), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT96), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT17), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n271), .A2(new_n293), .A3(new_n272), .ZN(new_n294));
  OAI211_X1 g093(.A(KEYINPUT17), .B(new_n265), .C1(new_n267), .C2(new_n268), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n291), .A2(new_n292), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n297), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT96), .B1(new_n299), .B2(new_n290), .ZN(new_n300));
  XNOR2_X1  g099(.A(G134gat), .B(G162gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  AND3_X1   g101(.A1(new_n298), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n302), .B1(new_n298), .B2(new_n300), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n256), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n298), .A2(new_n300), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(new_n301), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n298), .A2(new_n300), .A3(new_n302), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n255), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G230gat), .A2(G233gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n311), .B(KEYINPUT98), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n286), .A2(new_n288), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(new_n221), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n284), .A2(KEYINPUT97), .A3(new_n285), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT97), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n281), .A2(new_n317), .A3(new_n283), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n316), .B(new_n318), .C1(new_n220), .C2(new_n211), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT10), .B1(new_n315), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT10), .ZN(new_n321));
  NOR3_X1   g120(.A1(new_n289), .A2(new_n321), .A3(new_n221), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n313), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  AND2_X1   g122(.A1(new_n315), .A2(new_n319), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n324), .A2(G230gat), .A3(G233gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G120gat), .B(G148gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(G176gat), .B(G204gat), .ZN(new_n328));
  XOR2_X1   g127(.A(new_n327), .B(new_n328), .Z(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT99), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n326), .A2(KEYINPUT99), .A3(new_n330), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n311), .B1(new_n320), .B2(new_n322), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n336), .A2(new_n325), .A3(new_n329), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n249), .A2(new_n310), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G229gat), .A2(G233gat), .ZN(new_n341));
  INV_X1    g140(.A(new_n240), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(new_n271), .A3(new_n272), .ZN(new_n343));
  INV_X1    g142(.A(new_n294), .ZN(new_n344));
  OAI21_X1  g143(.A(KEYINPUT87), .B1(new_n238), .B2(new_n239), .ZN(new_n345));
  INV_X1    g144(.A(new_n239), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT87), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n346), .A2(new_n347), .A3(new_n237), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n345), .A2(new_n348), .A3(new_n295), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n341), .B(new_n343), .C1(new_n344), .C2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT18), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  XOR2_X1   g151(.A(new_n341), .B(KEYINPUT13), .Z(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n273), .A2(new_n240), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n354), .B1(new_n343), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G113gat), .B(G141gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(G197gat), .ZN(new_n359));
  XOR2_X1   g158(.A(KEYINPUT11), .B(G169gat), .Z(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(KEYINPUT12), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n294), .A2(new_n295), .A3(new_n348), .A4(new_n345), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n363), .A2(KEYINPUT18), .A3(new_n341), .A4(new_n343), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n352), .A2(new_n357), .A3(new_n362), .A4(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n356), .B1(new_n350), .B2(new_n351), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n362), .B1(new_n367), .B2(new_n364), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G169gat), .A2(G176gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(G169gat), .A2(G176gat), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT26), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AND2_X1   g172(.A1(KEYINPUT67), .A2(KEYINPUT26), .ZN(new_n374));
  NOR2_X1   g173(.A1(KEYINPUT67), .A2(KEYINPUT26), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n371), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT68), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI211_X1 g177(.A(KEYINPUT68), .B(new_n371), .C1(new_n374), .C2(new_n375), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n373), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT27), .B(G183gat), .ZN(new_n381));
  INV_X1    g180(.A(G190gat), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT28), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT66), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT66), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT28), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n381), .A2(new_n382), .A3(new_n384), .A4(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(G183gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT27), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT27), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(G183gat), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(new_n391), .A3(new_n382), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n384), .A2(new_n386), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G183gat), .A2(G190gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n387), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n380), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(G169gat), .ZN(new_n399));
  INV_X1    g198(.A(G176gat), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(new_n400), .A3(KEYINPUT23), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT23), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n402), .B1(G169gat), .B2(G176gat), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT24), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n404), .A2(G183gat), .A3(G190gat), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n401), .A2(new_n403), .A3(new_n405), .A4(new_n370), .ZN(new_n406));
  AND2_X1   g205(.A1(G183gat), .A2(G190gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(G183gat), .A2(G190gat), .ZN(new_n408));
  NOR3_X1   g207(.A1(new_n407), .A2(new_n408), .A3(new_n404), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT64), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT25), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI211_X1 g211(.A(KEYINPUT64), .B(KEYINPUT25), .C1(new_n406), .C2(new_n409), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n412), .A2(KEYINPUT65), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT65), .B1(new_n412), .B2(new_n413), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n398), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(G134gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(G127gat), .ZN(new_n418));
  INV_X1    g217(.A(G127gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(G134gat), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT1), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n418), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(G113gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT71), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT71), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(G113gat), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n424), .A2(new_n426), .A3(G120gat), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT70), .B1(new_n423), .B2(G120gat), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT70), .ZN(new_n429));
  INV_X1    g228(.A(G120gat), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(new_n430), .A3(G113gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n422), .B1(new_n427), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT69), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n420), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n417), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(G113gat), .B(G120gat), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n435), .B(new_n436), .C1(KEYINPUT1), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n416), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(G227gat), .ZN(new_n442));
  INV_X1    g241(.A(G233gat), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n398), .B(new_n439), .C1(new_n414), .C2(new_n415), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n441), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT32), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT33), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g248(.A(G15gat), .B(G43gat), .Z(new_n450));
  XNOR2_X1  g249(.A(G71gat), .B(G99gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n447), .A2(new_n449), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n452), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n446), .B(KEYINPUT32), .C1(new_n448), .C2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT72), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n445), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n458), .B1(new_n442), .B2(new_n443), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT34), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT34), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n458), .B(new_n461), .C1(new_n442), .C2(new_n443), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n457), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g264(.A1(G155gat), .A2(G162gat), .ZN(new_n466));
  NOR2_X1   g265(.A1(G155gat), .A2(G162gat), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OR2_X1    g267(.A1(G141gat), .A2(G148gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(G141gat), .A2(G148gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(KEYINPUT76), .B(KEYINPUT2), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n468), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(G155gat), .B(G162gat), .ZN(new_n474));
  INV_X1    g273(.A(G155gat), .ZN(new_n475));
  INV_X1    g274(.A(G162gat), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT2), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n474), .A2(new_n469), .A3(new_n477), .A4(new_n470), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(G197gat), .B(G204gat), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT22), .ZN(new_n481));
  INV_X1    g280(.A(G211gat), .ZN(new_n482));
  INV_X1    g281(.A(G218gat), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G211gat), .B(G218gat), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n486), .A2(new_n480), .A3(new_n484), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT29), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n479), .B1(new_n490), .B2(KEYINPUT3), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n488), .A2(new_n489), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT73), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n492), .B(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT3), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n473), .A2(new_n495), .A3(new_n478), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT29), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n491), .B1(new_n494), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(G228gat), .A3(G233gat), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n491), .A2(KEYINPUT81), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n491), .A2(KEYINPUT81), .ZN(new_n503));
  INV_X1    g302(.A(new_n492), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n498), .A2(new_n504), .B1(G228gat), .B2(G233gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n502), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G78gat), .B(G106gat), .ZN(new_n510));
  INV_X1    g309(.A(G50gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(G22gat), .ZN(new_n513));
  INV_X1    g312(.A(new_n508), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n501), .A2(new_n506), .A3(new_n514), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n509), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n513), .B1(new_n509), .B2(new_n515), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n456), .A2(KEYINPUT72), .A3(new_n463), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n465), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n494), .ZN(new_n522));
  NAND2_X1  g321(.A1(G226gat), .A2(G233gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(KEYINPUT74), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n524), .B1(new_n416), .B2(new_n497), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n412), .A2(new_n413), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n524), .B1(new_n526), .B2(new_n397), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n522), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n497), .B1(new_n526), .B2(new_n397), .ZN(new_n530));
  INV_X1    g329(.A(new_n524), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT65), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n403), .A2(new_n370), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n388), .A2(new_n382), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n535), .A2(KEYINPUT24), .A3(new_n395), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n534), .A2(new_n536), .A3(new_n405), .A4(new_n401), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT25), .B1(new_n537), .B2(KEYINPUT64), .ZN(new_n538));
  INV_X1    g337(.A(new_n413), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n533), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n412), .A2(KEYINPUT65), .A3(new_n413), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n397), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n532), .B(new_n492), .C1(new_n542), .C2(new_n531), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT75), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n416), .A2(new_n524), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n546), .A2(KEYINPUT75), .A3(new_n492), .A4(new_n532), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n529), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G8gat), .B(G36gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(G64gat), .B(G92gat), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n549), .B(new_n550), .Z(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n529), .A2(new_n545), .A3(new_n551), .A4(new_n547), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(KEYINPUT30), .A3(new_n554), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n529), .A2(new_n547), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT30), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n556), .A2(new_n557), .A3(new_n551), .A4(new_n545), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n433), .A2(new_n473), .A3(new_n438), .A4(new_n478), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT4), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n473), .A2(new_n478), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n563), .A2(KEYINPUT4), .A3(new_n438), .A4(new_n433), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT5), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT77), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n567), .B1(new_n479), .B2(KEYINPUT3), .ZN(new_n568));
  AOI211_X1 g367(.A(KEYINPUT77), .B(new_n495), .C1(new_n473), .C2(new_n478), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n496), .B(new_n439), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(G225gat), .A2(G233gat), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n565), .A2(new_n566), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n438), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n418), .A2(new_n420), .A3(new_n421), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n428), .A2(new_n431), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n424), .A2(new_n426), .A3(G120gat), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n479), .B1(new_n573), .B2(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n571), .B1(new_n578), .B2(new_n560), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n566), .B1(new_n579), .B2(KEYINPUT78), .ZN(new_n580));
  INV_X1    g379(.A(new_n571), .ZN(new_n581));
  INV_X1    g380(.A(new_n560), .ZN(new_n582));
  AOI22_X1  g381(.A1(new_n433), .A2(new_n438), .B1(new_n473), .B2(new_n478), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT78), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n580), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n439), .A2(new_n496), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n479), .A2(KEYINPUT3), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT77), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n479), .A2(new_n567), .A3(KEYINPUT3), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n588), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n562), .A2(new_n564), .ZN(new_n593));
  NOR3_X1   g392(.A1(new_n592), .A2(new_n593), .A3(new_n581), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n572), .B1(new_n587), .B2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G1gat), .B(G29gat), .Z(new_n596));
  XNOR2_X1  g395(.A(G57gat), .B(G85gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT6), .ZN(new_n602));
  INV_X1    g401(.A(new_n600), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n603), .B(new_n572), .C1(new_n587), .C2(new_n594), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n601), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n595), .A2(KEYINPUT6), .A3(new_n600), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n559), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(KEYINPUT35), .B1(new_n521), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n464), .A2(new_n456), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n463), .A2(new_n453), .A3(new_n455), .ZN(new_n611));
  AOI22_X1  g410(.A1(new_n610), .A2(new_n611), .B1(new_n555), .B2(new_n558), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n605), .A2(new_n606), .ZN(new_n613));
  NOR3_X1   g412(.A1(new_n613), .A2(new_n518), .A3(KEYINPUT35), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n609), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n531), .B1(new_n542), .B2(KEYINPUT29), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n617), .A2(new_n494), .A3(new_n527), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n542), .A2(new_n531), .ZN(new_n619));
  INV_X1    g418(.A(new_n532), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n504), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT38), .B1(new_n622), .B2(KEYINPUT37), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n623), .B(new_n552), .C1(KEYINPUT37), .C2(new_n548), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n605), .A2(new_n554), .A3(new_n606), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n552), .A2(KEYINPUT37), .ZN(new_n626));
  AOI22_X1  g425(.A1(new_n553), .A2(new_n626), .B1(KEYINPUT37), .B2(new_n548), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT38), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n624), .B(new_n625), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT82), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n565), .A2(new_n570), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n631), .B1(new_n632), .B2(new_n581), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n631), .B(new_n581), .C1(new_n592), .C2(new_n593), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n630), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n581), .B1(new_n592), .B2(new_n593), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(KEYINPUT82), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n582), .A2(new_n583), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n630), .B1(new_n639), .B2(new_n571), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n638), .A2(new_n634), .A3(new_n640), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n636), .A2(KEYINPUT40), .A3(new_n603), .A4(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT83), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n638), .A2(new_n634), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n600), .B1(new_n645), .B2(new_n630), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n646), .A2(KEYINPUT83), .A3(KEYINPUT40), .A4(new_n641), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n636), .A2(new_n603), .A3(new_n641), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT40), .ZN(new_n650));
  AOI22_X1  g449(.A1(new_n649), .A2(new_n650), .B1(new_n600), .B2(new_n595), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n648), .A2(new_n558), .A3(new_n555), .A4(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n629), .A2(new_n652), .A3(new_n519), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n465), .A2(KEYINPUT36), .A3(new_n520), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT36), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n610), .A2(new_n655), .A3(new_n611), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n608), .A2(new_n518), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n653), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n369), .B1(new_n616), .B2(new_n659), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n660), .A2(KEYINPUT88), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(KEYINPUT88), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n340), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n607), .B(KEYINPUT100), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  INV_X1    g465(.A(new_n663), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT101), .B(KEYINPUT16), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(G8gat), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n667), .A2(new_n559), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(G8gat), .ZN(new_n671));
  INV_X1    g470(.A(new_n559), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n671), .B1(new_n663), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT42), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(KEYINPUT42), .B2(new_n670), .ZN(G1325gat));
  NAND2_X1  g474(.A1(new_n610), .A2(new_n611), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  OR3_X1    g476(.A1(new_n667), .A2(G15gat), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(G15gat), .B1(new_n667), .B2(new_n657), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(G1326gat));
  NAND2_X1  g479(.A1(new_n663), .A2(new_n518), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT43), .B(G22gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  NOR2_X1   g482(.A1(new_n249), .A2(new_n338), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n305), .A2(new_n309), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n686), .B1(new_n661), .B2(new_n662), .ZN(new_n687));
  INV_X1    g486(.A(G29gat), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n687), .A2(new_n688), .A3(new_n664), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT45), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n616), .A2(new_n659), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n691), .B1(new_n692), .B2(new_n685), .ZN(new_n693));
  AND3_X1   g492(.A1(new_n456), .A2(KEYINPUT72), .A3(new_n463), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n463), .B1(new_n456), .B2(KEYINPUT72), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n694), .A2(new_n695), .A3(new_n655), .ZN(new_n696));
  AND3_X1   g495(.A1(new_n610), .A2(new_n655), .A3(new_n611), .ZN(new_n697));
  AOI22_X1  g496(.A1(new_n555), .A2(new_n558), .B1(new_n606), .B2(new_n605), .ZN(new_n698));
  OAI22_X1  g497(.A1(new_n696), .A2(new_n697), .B1(new_n519), .B2(new_n698), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n629), .A2(new_n652), .A3(new_n519), .ZN(new_n700));
  OAI21_X1  g499(.A(KEYINPUT102), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  AOI22_X1  g500(.A1(new_n654), .A2(new_n656), .B1(new_n608), .B2(new_n518), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT102), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n702), .A2(new_n703), .A3(new_n653), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n698), .A2(new_n519), .A3(new_n465), .A4(new_n520), .ZN(new_n705));
  AOI221_X4 g504(.A(KEYINPUT103), .B1(new_n612), .B2(new_n614), .C1(new_n705), .C2(KEYINPUT35), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n707), .B1(new_n609), .B2(new_n615), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n701), .B(new_n704), .C1(new_n706), .C2(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n310), .A2(KEYINPUT44), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n693), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n684), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n369), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(KEYINPUT104), .B1(new_n711), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT104), .ZN(new_n716));
  INV_X1    g515(.A(new_n710), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n702), .A2(new_n703), .A3(new_n653), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n703), .B1(new_n702), .B2(new_n653), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n616), .A2(KEYINPUT103), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n609), .A2(new_n707), .A3(new_n615), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n717), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n716), .B(new_n713), .C1(new_n724), .C2(new_n693), .ZN(new_n725));
  AND3_X1   g524(.A1(new_n715), .A2(new_n664), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n690), .B1(new_n688), .B2(new_n726), .ZN(G1328gat));
  INV_X1    g526(.A(KEYINPUT46), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(KEYINPUT105), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n559), .A2(G36gat), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n687), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n728), .A2(KEYINPUT105), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n731), .B(new_n732), .Z(new_n733));
  NAND3_X1  g532(.A1(new_n715), .A2(new_n672), .A3(new_n725), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(G36gat), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(G1329gat));
  NAND2_X1  g535(.A1(new_n709), .A2(new_n710), .ZN(new_n737));
  INV_X1    g536(.A(new_n693), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n713), .ZN(new_n740));
  OAI21_X1  g539(.A(G43gat), .B1(new_n740), .B2(new_n657), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n677), .A2(G43gat), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n687), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n741), .A2(KEYINPUT47), .A3(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n743), .ZN(new_n745));
  INV_X1    g544(.A(new_n657), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n715), .A2(new_n746), .A3(new_n725), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n745), .B1(new_n747), .B2(G43gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n744), .B1(new_n748), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI211_X1 g548(.A(KEYINPUT48), .B(G50gat), .C1(new_n740), .C2(new_n519), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n518), .A2(new_n511), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT106), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT48), .ZN(new_n753));
  AOI22_X1  g552(.A1(new_n687), .A2(new_n752), .B1(KEYINPUT107), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n687), .A2(KEYINPUT107), .A3(new_n752), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n715), .A2(new_n518), .A3(new_n725), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n756), .B1(new_n757), .B2(G50gat), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n755), .B1(new_n758), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g558(.A(new_n369), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(new_n339), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n709), .A2(new_n249), .A3(new_n310), .A4(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n664), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n764), .B(G57gat), .Z(G1332gat));
  AOI21_X1  g564(.A(new_n559), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT108), .ZN(new_n767));
  OR3_X1    g566(.A1(new_n762), .A2(KEYINPUT109), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(KEYINPUT109), .B1(new_n762), .B2(new_n767), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1333gat));
  OAI21_X1  g571(.A(G71gat), .B1(new_n762), .B2(new_n657), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n676), .A2(new_n208), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n762), .B2(new_n774), .ZN(new_n775));
  XOR2_X1   g574(.A(new_n775), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g575(.A1(new_n762), .A2(new_n519), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(new_n209), .ZN(G1335gat));
  INV_X1    g577(.A(new_n761), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n711), .A2(new_n249), .A3(new_n779), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n780), .A2(new_n664), .ZN(new_n781));
  NOR2_X1   g580(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n249), .A2(new_n760), .A3(new_n310), .ZN(new_n785));
  AND3_X1   g584(.A1(new_n709), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n784), .B1(new_n709), .B2(new_n785), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n783), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n338), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n664), .A2(new_n275), .ZN(new_n790));
  OAI22_X1  g589(.A1(new_n781), .A2(new_n275), .B1(new_n789), .B2(new_n790), .ZN(G1336gat));
  NOR2_X1   g590(.A1(new_n559), .A2(G92gat), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n788), .A2(new_n338), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n779), .A2(new_n249), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n739), .A2(new_n672), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(G92gat), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT52), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n793), .A2(new_n799), .A3(new_n796), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(G1337gat));
  NAND2_X1  g600(.A1(new_n780), .A2(new_n746), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(G99gat), .ZN(new_n803));
  OR2_X1    g602(.A1(new_n677), .A2(G99gat), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n803), .B1(new_n789), .B2(new_n804), .ZN(G1338gat));
  NOR2_X1   g604(.A1(new_n519), .A2(G106gat), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n788), .A2(new_n338), .A3(new_n806), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n518), .B(new_n794), .C1(new_n724), .C2(new_n693), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(G106gat), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT53), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n808), .A2(KEYINPUT111), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT111), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n739), .A2(new_n813), .A3(new_n518), .A4(new_n794), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n812), .A2(G106gat), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n815), .A2(new_n816), .A3(new_n807), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n811), .A2(new_n817), .ZN(G1339gat));
  INV_X1    g617(.A(new_n249), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n314), .B(KEYINPUT10), .C1(new_n220), .C2(new_n211), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n820), .B(new_n312), .C1(new_n324), .C2(KEYINPUT10), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(KEYINPUT54), .A3(new_n336), .ZN(new_n822));
  XNOR2_X1  g621(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n313), .B(new_n823), .C1(new_n320), .C2(new_n322), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n824), .A2(KEYINPUT113), .A3(new_n330), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT113), .B1(new_n824), .B2(new_n330), .ZN(new_n827));
  OAI211_X1 g626(.A(KEYINPUT55), .B(new_n822), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n821), .A2(new_n336), .A3(KEYINPUT54), .ZN(new_n829));
  INV_X1    g628(.A(new_n827), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n829), .B1(new_n830), .B2(new_n825), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n828), .B(new_n337), .C1(new_n831), .C2(KEYINPUT55), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT114), .ZN(new_n833));
  INV_X1    g632(.A(new_n337), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n830), .A2(new_n825), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n829), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n834), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n826), .A2(new_n827), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n836), .B1(new_n839), .B2(new_n829), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT114), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n838), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n833), .A2(new_n760), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n341), .B1(new_n363), .B2(new_n343), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n343), .A2(new_n355), .A3(new_n354), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n361), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n365), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n338), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n685), .B1(new_n843), .B2(new_n848), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n685), .A2(new_n833), .A3(new_n847), .A4(new_n842), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n819), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n340), .A2(new_n760), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n518), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n855), .A2(new_n664), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n694), .A2(new_n695), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n856), .A2(new_n559), .A3(new_n857), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n858), .A2(new_n424), .A3(new_n426), .A4(new_n760), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n856), .A2(new_n612), .ZN(new_n860));
  OAI21_X1  g659(.A(G113gat), .B1(new_n860), .B2(new_n369), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(G1340gat));
  NOR3_X1   g661(.A1(new_n860), .A2(new_n430), .A3(new_n339), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n858), .A2(new_n338), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n863), .B1(new_n864), .B2(new_n430), .ZN(G1341gat));
  OAI21_X1  g664(.A(G127gat), .B1(new_n860), .B2(new_n819), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n819), .A2(G127gat), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n856), .A2(new_n559), .A3(new_n857), .A4(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT115), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n866), .A2(KEYINPUT115), .A3(new_n868), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(G1342gat));
  NOR2_X1   g672(.A1(new_n672), .A2(new_n310), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n856), .A2(new_n417), .A3(new_n857), .A4(new_n874), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n875), .A2(KEYINPUT56), .ZN(new_n876));
  OAI21_X1  g675(.A(G134gat), .B1(new_n860), .B2(new_n310), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(KEYINPUT56), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(G1343gat));
  INV_X1    g678(.A(KEYINPUT58), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n519), .B1(new_n852), .B2(new_n854), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n746), .A2(new_n763), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n369), .A2(G141gat), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n883), .A2(new_n559), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n852), .A2(new_n854), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT57), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n887), .A3(new_n518), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n882), .A2(new_n559), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n848), .B1(new_n832), .B2(new_n369), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n310), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n249), .B1(new_n891), .B2(new_n850), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n518), .B1(new_n892), .B2(new_n853), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n889), .B1(new_n893), .B2(KEYINPUT57), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n888), .A2(new_n894), .A3(new_n760), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT117), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(G141gat), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n895), .A2(new_n896), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n880), .B(new_n885), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n895), .A2(G141gat), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n885), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT116), .B1(new_n902), .B2(KEYINPUT58), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT116), .ZN(new_n904));
  AOI211_X1 g703(.A(new_n904), .B(new_n880), .C1(new_n901), .C2(new_n885), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n900), .B1(new_n903), .B2(new_n905), .ZN(G1344gat));
  INV_X1    g705(.A(G148gat), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n883), .A2(new_n907), .A3(new_n559), .A4(new_n338), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n888), .A2(new_n894), .A3(new_n338), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n907), .A2(KEYINPUT59), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n685), .A2(new_n847), .A3(new_n840), .A4(new_n838), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n249), .B1(new_n891), .B2(new_n913), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n887), .B(new_n518), .C1(new_n914), .C2(new_n853), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n657), .A2(new_n664), .A3(KEYINPUT118), .A4(new_n559), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n338), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(new_n889), .B2(new_n918), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n915), .B(new_n919), .C1(new_n881), .C2(new_n887), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n912), .B1(new_n920), .B2(G148gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n908), .B1(new_n911), .B2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g723(.A(KEYINPUT119), .B(new_n908), .C1(new_n911), .C2(new_n921), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1345gat));
  NAND3_X1  g725(.A1(new_n883), .A2(new_n559), .A3(new_n249), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n888), .A2(new_n894), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n249), .A2(G155gat), .ZN(new_n929));
  XOR2_X1   g728(.A(new_n929), .B(KEYINPUT120), .Z(new_n930));
  AOI22_X1  g729(.A1(new_n927), .A2(new_n475), .B1(new_n928), .B2(new_n930), .ZN(G1346gat));
  NAND3_X1  g730(.A1(new_n883), .A2(new_n476), .A3(new_n874), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n928), .A2(new_n685), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n933), .B2(new_n476), .ZN(G1347gat));
  NAND2_X1  g733(.A1(new_n763), .A2(new_n672), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n935), .A2(new_n677), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n855), .A2(new_n936), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n937), .A2(new_n399), .A3(new_n369), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n664), .B1(new_n852), .B2(new_n854), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n521), .A2(new_n559), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT121), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(new_n760), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n938), .B1(new_n399), .B2(new_n944), .ZN(G1348gat));
  INV_X1    g744(.A(new_n937), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n946), .A2(G176gat), .A3(new_n338), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n947), .A2(KEYINPUT122), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n947), .A2(KEYINPUT122), .ZN(new_n949));
  AOI21_X1  g748(.A(G176gat), .B1(new_n943), .B2(new_n338), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(G1349gat));
  INV_X1    g750(.A(KEYINPUT123), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(KEYINPUT60), .ZN(new_n953));
  XOR2_X1   g752(.A(new_n953), .B(KEYINPUT124), .Z(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n388), .B1(new_n946), .B2(new_n249), .ZN(new_n956));
  INV_X1    g755(.A(new_n381), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n942), .A2(new_n957), .A3(new_n819), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n952), .A2(KEYINPUT60), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n955), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI221_X1 g760(.A(new_n954), .B1(new_n952), .B2(KEYINPUT60), .C1(new_n956), .C2(new_n958), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1350gat));
  NAND3_X1  g762(.A1(new_n943), .A2(new_n382), .A3(new_n685), .ZN(new_n964));
  OAI21_X1  g763(.A(G190gat), .B1(new_n937), .B2(new_n310), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n965), .A2(KEYINPUT61), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n965), .A2(KEYINPUT61), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n964), .B1(new_n966), .B2(new_n967), .ZN(G1351gat));
  OR2_X1    g767(.A1(new_n881), .A2(new_n887), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n746), .A2(new_n935), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n969), .A2(new_n915), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n760), .A2(G197gat), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n746), .A2(new_n519), .A3(new_n559), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n939), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n974), .A2(new_n369), .ZN(new_n975));
  OAI22_X1  g774(.A1(new_n971), .A2(new_n972), .B1(new_n975), .B2(G197gat), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(G1352gat));
  NOR2_X1   g776(.A1(new_n339), .A2(G204gat), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n886), .A2(new_n763), .A3(new_n973), .A4(new_n978), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT125), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n979), .B(new_n980), .ZN(new_n981));
  OAI21_X1  g780(.A(KEYINPUT126), .B1(new_n981), .B2(KEYINPUT62), .ZN(new_n982));
  OR2_X1    g781(.A1(new_n979), .A2(new_n980), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT62), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n979), .A2(new_n980), .ZN(new_n986));
  NAND4_X1  g785(.A1(new_n983), .A2(new_n984), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n982), .A2(new_n987), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n969), .A2(new_n338), .A3(new_n915), .A4(new_n970), .ZN(new_n989));
  AOI22_X1  g788(.A1(new_n981), .A2(KEYINPUT62), .B1(new_n989), .B2(G204gat), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n988), .A2(new_n990), .ZN(G1353gat));
  INV_X1    g790(.A(new_n974), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n992), .A2(new_n482), .A3(new_n249), .ZN(new_n993));
  NAND4_X1  g792(.A1(new_n969), .A2(new_n249), .A3(new_n915), .A4(new_n970), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT63), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n995), .A2(KEYINPUT127), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n482), .B1(KEYINPUT127), .B2(new_n995), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n994), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  INV_X1    g797(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g798(.A(new_n996), .B1(new_n994), .B2(new_n997), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n993), .B1(new_n999), .B2(new_n1000), .ZN(G1354gat));
  OAI21_X1  g800(.A(G218gat), .B1(new_n971), .B2(new_n310), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n992), .A2(new_n483), .A3(new_n685), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1002), .A2(new_n1003), .ZN(G1355gat));
endmodule


