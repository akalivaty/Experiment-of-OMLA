//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 1 1 0 1 0 1 0 0 1 1 1 0 1 1 0 0 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n864, new_n865, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984, new_n985;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  AND2_X1   g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  NOR3_X1   g005(.A1(new_n205), .A2(new_n206), .A3(KEYINPUT26), .ZN(new_n207));
  AOI211_X1 g006(.A(new_n204), .B(new_n207), .C1(KEYINPUT26), .C2(new_n206), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT27), .B(G183gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT69), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT28), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT70), .ZN(new_n215));
  INV_X1    g014(.A(G183gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT27), .ZN(new_n217));
  AOI211_X1 g016(.A(KEYINPUT28), .B(G190gat), .C1(new_n217), .C2(KEYINPUT68), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(KEYINPUT68), .B2(new_n209), .ZN(new_n219));
  AND3_X1   g018(.A1(new_n214), .A2(new_n215), .A3(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n215), .B1(new_n214), .B2(new_n219), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n208), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G113gat), .B(G120gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  XNOR2_X1  g023(.A(G127gat), .B(G134gat), .ZN(new_n225));
  XOR2_X1   g024(.A(new_n224), .B(new_n225), .Z(new_n226));
  NAND3_X1  g025(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(G183gat), .B2(G190gat), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n204), .A2(KEYINPUT66), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT24), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n204), .A2(KEYINPUT66), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n228), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(new_n233), .B2(new_n232), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n206), .A2(KEYINPUT23), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n206), .A2(KEYINPUT23), .ZN(new_n237));
  NOR3_X1   g036(.A1(new_n236), .A2(new_n237), .A3(new_n205), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n235), .A2(KEYINPUT25), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n228), .B1(new_n230), .B2(new_n203), .ZN(new_n240));
  OR2_X1    g039(.A1(new_n240), .A2(KEYINPUT65), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(KEYINPUT65), .ZN(new_n242));
  AND3_X1   g041(.A1(new_n241), .A2(new_n242), .A3(new_n238), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n239), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n222), .A2(new_n226), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT71), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n222), .A2(KEYINPUT71), .A3(new_n226), .A4(new_n245), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n222), .A2(new_n245), .ZN(new_n250));
  INV_X1    g049(.A(new_n226), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n248), .A2(new_n249), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G227gat), .A2(G233gat), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  OR3_X1    g054(.A1(new_n253), .A2(KEYINPUT34), .A3(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(KEYINPUT34), .B1(new_n253), .B2(new_n255), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT33), .B1(new_n253), .B2(new_n255), .ZN(new_n259));
  XNOR2_X1  g058(.A(G15gat), .B(G43gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(G71gat), .B(G99gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n253), .A2(new_n255), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT32), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n256), .B(new_n257), .C1(new_n259), .C2(new_n262), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n264), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n267), .B1(new_n264), .B2(new_n268), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n202), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n264), .A2(new_n268), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(new_n266), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n264), .A2(new_n267), .A3(new_n268), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(KEYINPUT36), .A3(new_n274), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT29), .ZN(new_n277));
  INV_X1    g076(.A(G141gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(G148gat), .ZN(new_n279));
  XOR2_X1   g078(.A(KEYINPUT75), .B(G148gat), .Z(new_n280));
  OAI21_X1  g079(.A(new_n279), .B1(new_n280), .B2(new_n278), .ZN(new_n281));
  XNOR2_X1  g080(.A(G155gat), .B(G162gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT2), .ZN(new_n284));
  AND2_X1   g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT77), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n281), .A2(KEYINPUT77), .A3(new_n285), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(G141gat), .B(G148gat), .Z(new_n291));
  XOR2_X1   g090(.A(KEYINPUT74), .B(KEYINPUT2), .Z(new_n292));
  AOI21_X1  g091(.A(new_n282), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n277), .B1(new_n295), .B2(KEYINPUT3), .ZN(new_n296));
  XNOR2_X1  g095(.A(G197gat), .B(G204gat), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT22), .ZN(new_n298));
  INV_X1    g097(.A(G211gat), .ZN(new_n299));
  INV_X1    g098(.A(G218gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G211gat), .B(G218gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n296), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT3), .ZN(new_n306));
  INV_X1    g105(.A(new_n304), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n307), .A2(KEYINPUT84), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n303), .A2(new_n297), .A3(new_n301), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT84), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n277), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n306), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n295), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n305), .A2(new_n313), .B1(G228gat), .B2(G233gat), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n306), .B1(new_n304), .B2(KEYINPUT29), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n295), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n316), .A2(G228gat), .A3(G233gat), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n317), .B1(new_n304), .B2(new_n296), .ZN(new_n318));
  OAI21_X1  g117(.A(G22gat), .B1(new_n314), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT85), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(G78gat), .B(G106gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT31), .B(G50gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n322), .B(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  OR3_X1    g124(.A1(new_n314), .A2(new_n318), .A3(G22gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(new_n319), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n325), .A2(new_n327), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G226gat), .A2(G233gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n250), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n333), .B(KEYINPUT73), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT72), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n250), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n222), .A2(KEYINPUT72), .A3(new_n245), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n331), .B1(new_n338), .B2(KEYINPUT29), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(new_n304), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n338), .A2(new_n332), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n250), .A2(new_n277), .A3(new_n331), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n304), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G8gat), .B(G36gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(G64gat), .B(G92gat), .ZN(new_n347));
  XOR2_X1   g146(.A(new_n346), .B(new_n347), .Z(new_n348));
  NAND3_X1  g147(.A1(new_n341), .A2(new_n345), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n348), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n307), .B1(new_n334), .B2(new_n339), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n350), .B1(new_n351), .B2(new_n344), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n349), .A2(KEYINPUT30), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT30), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n341), .A2(new_n354), .A3(new_n345), .A4(new_n348), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT88), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n293), .B1(new_n288), .B2(new_n289), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n226), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT79), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n358), .A2(new_n361), .A3(new_n226), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n360), .A2(KEYINPUT4), .A3(new_n362), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n363), .B(KEYINPUT83), .C1(KEYINPUT4), .C2(new_n359), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n226), .B1(new_n295), .B2(KEYINPUT3), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n365), .B1(KEYINPUT3), .B2(new_n295), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT83), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n360), .A2(new_n367), .A3(KEYINPUT4), .A4(new_n362), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n364), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G225gat), .A2(G233gat), .ZN(new_n370));
  XOR2_X1   g169(.A(new_n370), .B(KEYINPUT78), .Z(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n371), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n295), .A2(new_n251), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n360), .A2(new_n373), .A3(new_n362), .A4(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT39), .B1(new_n375), .B2(KEYINPUT87), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n376), .B1(KEYINPUT87), .B2(new_n375), .ZN(new_n377));
  AND2_X1   g176(.A1(new_n372), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT39), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n369), .A2(new_n379), .A3(new_n371), .ZN(new_n380));
  XNOR2_X1  g179(.A(G1gat), .B(G29gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(KEYINPUT0), .ZN(new_n382));
  XNOR2_X1  g181(.A(G57gat), .B(G85gat), .ZN(new_n383));
  XOR2_X1   g182(.A(new_n382), .B(new_n383), .Z(new_n384));
  XOR2_X1   g183(.A(new_n384), .B(KEYINPUT86), .Z(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n357), .B(KEYINPUT40), .C1(new_n378), .C2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n377), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(new_n386), .A3(new_n380), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT40), .B1(new_n391), .B2(new_n357), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n356), .A2(new_n393), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n366), .A2(new_n373), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT4), .B1(new_n360), .B2(new_n362), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT80), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n359), .A2(KEYINPUT4), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n399), .B1(new_n396), .B2(new_n397), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n395), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT81), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI211_X1 g202(.A(KEYINPUT81), .B(new_n395), .C1(new_n398), .C2(new_n400), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n360), .A2(new_n362), .A3(new_n374), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n371), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT5), .ZN(new_n407));
  OR2_X1    g206(.A1(new_n407), .A2(KEYINPUT82), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(KEYINPUT82), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n403), .A2(new_n404), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT5), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n364), .A2(new_n395), .A3(new_n411), .A4(new_n368), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n410), .A2(KEYINPUT89), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT89), .B1(new_n410), .B2(new_n412), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n385), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n330), .B1(new_n394), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n410), .A2(new_n384), .A3(new_n412), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT6), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n384), .B1(new_n410), .B2(new_n412), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT6), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n350), .A2(KEYINPUT37), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n352), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT37), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n428), .B1(new_n341), .B2(new_n345), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT38), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n349), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n340), .A2(new_n307), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n342), .A2(new_n343), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n428), .B1(new_n433), .B2(new_n304), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT38), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n431), .B1(new_n426), .B2(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n422), .A2(new_n424), .A3(new_n430), .A4(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n276), .B1(new_n417), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n410), .A2(new_n412), .ZN(new_n439));
  INV_X1    g238(.A(new_n384), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n441), .A2(new_n419), .A3(new_n418), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n424), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n356), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n330), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n438), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n330), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n273), .A2(new_n447), .A3(new_n274), .ZN(new_n448));
  INV_X1    g247(.A(new_n356), .ZN(new_n449));
  NOR3_X1   g248(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT35), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT89), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n439), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n386), .B1(new_n452), .B2(new_n413), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n424), .B1(new_n453), .B2(new_n420), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n269), .A2(new_n270), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n456), .A2(KEYINPUT90), .A3(new_n447), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT90), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n448), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n444), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT35), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n455), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(G57gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(G64gat), .ZN(new_n465));
  INV_X1    g264(.A(G64gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(G57gat), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT9), .ZN(new_n468));
  NAND2_X1  g267(.A1(G71gat), .A2(G78gat), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n465), .A2(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n469), .ZN(new_n471));
  NOR2_X1   g270(.A1(G71gat), .A2(G78gat), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT97), .ZN(new_n473));
  NOR3_X1   g272(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(G71gat), .ZN(new_n475));
  INV_X1    g274(.A(G78gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT97), .B1(new_n477), .B2(new_n469), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n470), .B1(new_n474), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT96), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n472), .B1(new_n480), .B2(new_n469), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n471), .A2(KEYINPUT96), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n471), .A2(KEYINPUT9), .ZN(new_n483));
  XNOR2_X1  g282(.A(G57gat), .B(G64gat), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n481), .B(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT21), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(G231gat), .A2(G233gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(G127gat), .ZN(new_n491));
  XOR2_X1   g290(.A(G183gat), .B(G211gat), .Z(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  OR2_X1    g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n491), .A2(new_n493), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G15gat), .B(G22gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(KEYINPUT93), .ZN(new_n498));
  INV_X1    g297(.A(G1gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT16), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n501), .A2(G1gat), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n500), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(G8gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n486), .A2(new_n487), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT98), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT98), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n505), .B(new_n509), .C1(new_n487), .C2(new_n486), .ZN(new_n510));
  XNOR2_X1  g309(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n511));
  XOR2_X1   g310(.A(new_n511), .B(G155gat), .Z(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n508), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n513), .B1(new_n508), .B2(new_n510), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n496), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n516), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n518), .A2(new_n494), .A3(new_n495), .A4(new_n514), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(G43gat), .B(G50gat), .Z(new_n522));
  INV_X1    g321(.A(KEYINPUT15), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(G29gat), .A2(G36gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT14), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n526), .A2(KEYINPUT91), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT92), .B(G29gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(G36gat), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(new_n526), .B2(KEYINPUT91), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n524), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n524), .A2(new_n526), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n522), .A2(new_n523), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(new_n529), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT17), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT99), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n537), .A2(G85gat), .A3(G92gat), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT100), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n539), .A2(KEYINPUT7), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT7), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n541), .A2(KEYINPUT100), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n538), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(G85gat), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n544), .A2(KEYINPUT99), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n541), .A2(KEYINPUT100), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n539), .A2(KEYINPUT7), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n545), .A2(new_n546), .A3(new_n547), .A4(G92gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  AND2_X1   g348(.A1(G99gat), .A2(G106gat), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT8), .ZN(new_n551));
  OAI22_X1  g350(.A1(new_n550), .A2(new_n551), .B1(G85gat), .B2(G92gat), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  OR2_X1    g353(.A1(G99gat), .A2(G106gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(G99gat), .A2(G106gat), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n555), .A2(KEYINPUT101), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT101), .ZN(new_n558));
  NOR2_X1   g357(.A1(G99gat), .A2(G106gat), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n558), .B1(new_n550), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n554), .A2(new_n562), .ZN(new_n563));
  AND4_X1   g362(.A1(KEYINPUT102), .A2(new_n549), .A3(new_n561), .A4(new_n553), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n552), .B1(new_n543), .B2(new_n548), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT102), .B1(new_n565), .B2(new_n561), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n563), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n536), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n549), .A2(new_n561), .A3(new_n553), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT102), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n565), .A2(KEYINPUT102), .A3(new_n561), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n571), .A2(new_n572), .B1(new_n562), .B2(new_n554), .ZN(new_n573));
  AND2_X1   g372(.A1(G232gat), .A2(G233gat), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n573), .A2(new_n535), .B1(KEYINPUT41), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n568), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G190gat), .B(G218gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT103), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n576), .A2(new_n578), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n574), .A2(KEYINPUT41), .ZN(new_n581));
  XNOR2_X1  g380(.A(G134gat), .B(G162gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  OR3_X1    g383(.A1(new_n579), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n584), .B1(new_n579), .B2(new_n580), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT104), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n521), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n588), .B1(new_n521), .B2(new_n587), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n571), .A2(new_n572), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT105), .ZN(new_n592));
  AOI22_X1  g391(.A1(new_n549), .A2(new_n553), .B1(new_n561), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n557), .A2(new_n560), .A3(KEYINPUT105), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n486), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n567), .A2(new_n486), .B1(new_n591), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G230gat), .A2(G233gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G120gat), .B(G148gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(G176gat), .B(G204gat), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n599), .B(new_n600), .Z(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n486), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n561), .A2(new_n592), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n554), .A2(new_n594), .A3(new_n605), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n604), .B(new_n606), .C1(new_n564), .C2(new_n566), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT10), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n607), .B(new_n608), .C1(new_n573), .C2(new_n604), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT106), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT106), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n596), .A2(new_n611), .A3(new_n608), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n486), .A2(new_n608), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n573), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT107), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n573), .A2(KEYINPUT107), .A3(new_n613), .ZN(new_n617));
  AOI22_X1  g416(.A1(new_n610), .A2(new_n612), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT108), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n597), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n616), .A2(new_n617), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n609), .A2(KEYINPUT106), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n611), .B1(new_n596), .B2(new_n608), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n624), .A2(KEYINPUT108), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n603), .B1(new_n620), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT109), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT109), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n628), .B(new_n603), .C1(new_n620), .C2(new_n625), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n601), .B(KEYINPUT110), .Z(new_n631));
  INV_X1    g430(.A(new_n597), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n618), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n631), .B1(new_n633), .B2(new_n598), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n506), .A2(new_n535), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n505), .A2(new_n531), .A3(new_n534), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT95), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n506), .A2(KEYINPUT95), .A3(new_n535), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(G229gat), .A2(G233gat), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n642), .B(KEYINPUT13), .Z(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n506), .A2(KEYINPUT94), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT94), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n505), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n645), .A2(new_n647), .A3(new_n536), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n648), .A2(KEYINPUT18), .A3(new_n642), .A4(new_n636), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n648), .A2(new_n642), .A3(new_n636), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT18), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n644), .A2(new_n649), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G113gat), .B(G141gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G197gat), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT11), .B(G169gat), .Z(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n657), .B(KEYINPUT12), .Z(new_n658));
  NAND2_X1  g457(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n658), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n644), .A2(new_n660), .A3(new_n652), .A4(new_n649), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NOR4_X1   g462(.A1(new_n589), .A2(new_n590), .A3(new_n635), .A4(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n463), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(new_n443), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(new_n499), .ZN(G1324gat));
  INV_X1    g466(.A(new_n665), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(new_n449), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n501), .A2(new_n504), .ZN(new_n670));
  NOR2_X1   g469(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n504), .B1(new_n668), .B2(new_n449), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT42), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n675), .B1(KEYINPUT42), .B2(new_n673), .ZN(G1325gat));
  AOI21_X1  g475(.A(G15gat), .B1(new_n668), .B2(new_n456), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n276), .A2(G15gat), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n678), .B(KEYINPUT111), .Z(new_n679));
  AOI21_X1  g478(.A(new_n677), .B1(new_n668), .B2(new_n679), .ZN(G1326gat));
  XNOR2_X1  g479(.A(KEYINPUT43), .B(G22gat), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n668), .A2(new_n330), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT112), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n683), .A2(KEYINPUT112), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n682), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n683), .A2(KEYINPUT112), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n688), .A2(new_n684), .A3(new_n681), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(new_n689), .ZN(G1327gat));
  AOI22_X1  g489(.A1(new_n442), .A2(new_n424), .B1(new_n355), .B2(new_n353), .ZN(new_n691));
  AOI21_X1  g490(.A(KEYINPUT90), .B1(new_n456), .B2(new_n447), .ZN(new_n692));
  NOR4_X1   g491(.A1(new_n269), .A2(new_n270), .A3(new_n458), .A4(new_n330), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT35), .ZN(new_n695));
  AOI22_X1  g494(.A1(new_n695), .A2(new_n455), .B1(new_n438), .B2(new_n445), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT44), .B1(new_n696), .B2(new_n587), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n391), .A2(new_n357), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT40), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n388), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n416), .A2(new_n355), .A3(new_n701), .A4(new_n353), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n426), .A2(new_n435), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n429), .B1(new_n352), .B2(new_n425), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT38), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n349), .B(new_n703), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n447), .B(new_n702), .C1(new_n454), .C2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n276), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT113), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n444), .A2(new_n709), .A3(new_n330), .ZN(new_n710));
  OAI21_X1  g509(.A(KEYINPUT113), .B1(new_n691), .B2(new_n447), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n707), .A2(new_n708), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n587), .B1(new_n462), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(KEYINPUT114), .B(KEYINPUT44), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n697), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n443), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n663), .A2(new_n521), .A3(new_n635), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n528), .ZN(new_n720));
  INV_X1    g519(.A(new_n587), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n463), .A2(new_n721), .A3(new_n718), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n722), .A2(new_n443), .A3(new_n528), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n723), .A2(KEYINPUT45), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(KEYINPUT45), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n720), .A2(new_n724), .A3(new_n725), .ZN(G1328gat));
  NOR3_X1   g525(.A1(new_n722), .A2(G36gat), .A3(new_n356), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT46), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n716), .A2(new_n449), .A3(new_n718), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(G36gat), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(G1329gat));
  NAND4_X1  g530(.A1(new_n716), .A2(G43gat), .A3(new_n276), .A4(new_n718), .ZN(new_n732));
  INV_X1    g531(.A(G43gat), .ZN(new_n733));
  INV_X1    g532(.A(new_n456), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n722), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT47), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT47), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n732), .A2(new_n738), .A3(new_n735), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(G1330gat));
  INV_X1    g539(.A(G50gat), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n447), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n716), .A2(new_n718), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT115), .ZN(new_n744));
  OR2_X1    g543(.A1(new_n744), .A2(KEYINPUT48), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n463), .A2(new_n330), .A3(new_n721), .A4(new_n718), .ZN(new_n746));
  AOI22_X1  g545(.A1(new_n746), .A2(new_n741), .B1(new_n744), .B2(KEYINPUT48), .ZN(new_n747));
  AND3_X1   g546(.A1(new_n743), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n745), .B1(new_n743), .B2(new_n747), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n748), .A2(new_n749), .ZN(G1331gat));
  INV_X1    g549(.A(new_n635), .ZN(new_n751));
  NOR4_X1   g550(.A1(new_n751), .A2(new_n589), .A3(new_n590), .A4(new_n662), .ZN(new_n752));
  AND4_X1   g551(.A1(new_n707), .A2(new_n708), .A3(new_n710), .A4(new_n711), .ZN(new_n753));
  AOI22_X1  g552(.A1(new_n694), .A2(KEYINPUT35), .B1(new_n454), .B2(new_n450), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(new_n443), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(new_n464), .ZN(G1332gat));
  NOR2_X1   g556(.A1(new_n755), .A2(new_n356), .ZN(new_n758));
  NOR2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  AND2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n758), .B2(new_n759), .ZN(G1333gat));
  OAI21_X1  g561(.A(G71gat), .B1(new_n755), .B2(new_n708), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n456), .A2(new_n475), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n763), .B1(new_n755), .B2(new_n764), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g565(.A1(new_n755), .A2(new_n447), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(new_n476), .ZN(G1335gat));
  NOR2_X1   g567(.A1(new_n662), .A2(new_n521), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n770), .A2(new_n751), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n713), .A2(new_n714), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n773), .B1(new_n463), .B2(new_n721), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n717), .B(new_n771), .C1(new_n772), .C2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT116), .ZN(new_n776));
  INV_X1    g575(.A(new_n771), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n777), .B1(new_n697), .B2(new_n715), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n778), .A2(new_n779), .A3(new_n717), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n776), .A2(G85gat), .A3(new_n780), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n721), .B(new_n769), .C1(new_n753), .C2(new_n754), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n713), .A2(KEYINPUT51), .A3(new_n769), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n786), .A2(new_n544), .A3(new_n717), .A4(new_n635), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n781), .A2(new_n787), .ZN(G1336gat));
  INV_X1    g587(.A(G92gat), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n789), .B1(new_n778), .B2(new_n449), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n356), .A2(G92gat), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  AOI211_X1 g591(.A(new_n751), .B(new_n792), .C1(new_n784), .C2(new_n785), .ZN(new_n793));
  OAI21_X1  g592(.A(KEYINPUT52), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n449), .B(new_n771), .C1(new_n772), .C2(new_n774), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(G92gat), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n786), .A2(new_n635), .A3(new_n791), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n794), .A2(new_n799), .ZN(G1337gat));
  NAND2_X1  g599(.A1(new_n778), .A2(new_n276), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(G99gat), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n734), .A2(G99gat), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n786), .A2(new_n635), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(G1338gat));
  INV_X1    g604(.A(G106gat), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n778), .B2(new_n330), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n447), .A2(new_n751), .A3(G106gat), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(KEYINPUT117), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n810), .B1(new_n784), .B2(new_n785), .ZN(new_n811));
  OAI21_X1  g610(.A(KEYINPUT53), .B1(new_n807), .B2(new_n811), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n330), .B(new_n771), .C1(new_n772), .C2(new_n774), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(G106gat), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n815));
  INV_X1    g614(.A(new_n811), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n812), .A2(new_n817), .ZN(G1339gat));
  NOR2_X1   g617(.A1(new_n641), .A2(new_n643), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n642), .B1(new_n648), .B2(new_n636), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n657), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n635), .A2(new_n661), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(new_n618), .B2(new_n632), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n824), .B1(new_n620), .B2(new_n625), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n601), .B1(new_n633), .B2(new_n823), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT55), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(KEYINPUT120), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT119), .B1(new_n827), .B2(new_n828), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n825), .A2(new_n832), .A3(KEYINPUT55), .A4(new_n826), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n662), .A2(new_n831), .A3(new_n630), .A4(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n822), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT121), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT121), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n837), .B(new_n822), .C1(new_n830), .C2(new_n834), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n836), .A2(new_n587), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n821), .A2(new_n661), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n830), .A2(new_n587), .A3(new_n840), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n831), .A2(new_n630), .A3(new_n833), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n521), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n589), .A2(new_n590), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n845), .A2(new_n663), .A3(new_n751), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n846), .B(new_n847), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n692), .A2(new_n693), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(new_n449), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n849), .A2(new_n717), .A3(new_n851), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT122), .ZN(new_n853));
  INV_X1    g652(.A(G113gat), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n853), .A2(new_n854), .A3(new_n662), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n448), .A2(new_n449), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n849), .A2(new_n717), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(G113gat), .B1(new_n857), .B2(new_n663), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n855), .A2(new_n858), .ZN(G1340gat));
  INV_X1    g658(.A(G120gat), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n853), .A2(new_n860), .A3(new_n635), .ZN(new_n861));
  OAI21_X1  g660(.A(G120gat), .B1(new_n857), .B2(new_n751), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(G1341gat));
  OAI21_X1  g662(.A(G127gat), .B1(new_n857), .B2(new_n520), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n520), .A2(G127gat), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(new_n852), .B2(new_n865), .ZN(G1342gat));
  INV_X1    g665(.A(new_n852), .ZN(new_n867));
  INV_X1    g666(.A(G134gat), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n868), .A3(new_n721), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n869), .A2(KEYINPUT56), .ZN(new_n870));
  OAI21_X1  g669(.A(G134gat), .B1(new_n857), .B2(new_n587), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(KEYINPUT56), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(G1343gat));
  OAI211_X1 g672(.A(new_n621), .B(new_n632), .C1(new_n622), .C2(new_n623), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT54), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n632), .B1(new_n624), .B2(KEYINPUT108), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n618), .A2(new_n619), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n624), .A2(new_n597), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n602), .B1(new_n879), .B2(KEYINPUT54), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT123), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT123), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n825), .A2(new_n882), .A3(new_n826), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n881), .A2(new_n828), .A3(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT124), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n881), .A2(KEYINPUT124), .A3(new_n883), .A4(new_n828), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI211_X1 g687(.A(KEYINPUT125), .B(new_n822), .C1(new_n888), .C2(new_n834), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n587), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n842), .A2(new_n886), .A3(new_n662), .A4(new_n887), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT125), .B1(new_n891), .B2(new_n822), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n843), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n848), .B1(new_n893), .B2(new_n520), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT57), .B1(new_n894), .B2(new_n447), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT57), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n896), .B(new_n330), .C1(new_n844), .C2(new_n848), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n276), .A2(new_n443), .A3(new_n449), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n895), .A2(new_n662), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(G141gat), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT126), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n844), .A2(new_n848), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n902), .A2(new_n447), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n903), .A2(new_n278), .A3(new_n662), .A4(new_n898), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n900), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n901), .A2(new_n905), .A3(KEYINPUT58), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT58), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n900), .B(new_n904), .C1(KEYINPUT126), .C2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(G1344gat));
  NAND2_X1  g708(.A1(new_n903), .A2(new_n898), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n280), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(new_n912), .A3(new_n635), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n895), .A2(new_n897), .A3(new_n898), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n914), .A2(new_n751), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n915), .A2(KEYINPUT59), .A3(new_n912), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT57), .B1(new_n902), .B2(new_n447), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n893), .A2(new_n520), .ZN(new_n919));
  INV_X1    g718(.A(new_n846), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n896), .B(new_n330), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n918), .A2(new_n921), .A3(new_n635), .A4(new_n898), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n917), .B1(new_n922), .B2(G148gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n913), .B1(new_n916), .B2(new_n923), .ZN(G1345gat));
  OAI21_X1  g723(.A(G155gat), .B1(new_n914), .B2(new_n520), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n520), .A2(G155gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n910), .B2(new_n926), .ZN(G1346gat));
  XOR2_X1   g726(.A(KEYINPUT76), .B(G162gat), .Z(new_n928));
  NAND3_X1  g727(.A1(new_n911), .A2(new_n721), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n914), .A2(new_n587), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n929), .B1(new_n928), .B2(new_n930), .ZN(G1347gat));
  NOR3_X1   g730(.A1(new_n717), .A2(new_n448), .A3(new_n356), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n849), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(G169gat), .B1(new_n933), .B2(new_n663), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n902), .A2(new_n717), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n850), .A2(new_n356), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n663), .A2(G169gat), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n935), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NOR4_X1   g740(.A1(new_n938), .A2(KEYINPUT127), .A3(G169gat), .A4(new_n663), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n934), .B1(new_n941), .B2(new_n942), .ZN(G1348gat));
  INV_X1    g742(.A(G176gat), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n939), .A2(new_n944), .A3(new_n635), .ZN(new_n945));
  INV_X1    g744(.A(new_n933), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(new_n635), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n945), .B1(new_n948), .B2(new_n944), .ZN(G1349gat));
  OAI21_X1  g748(.A(G183gat), .B1(new_n933), .B2(new_n520), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n521), .A2(new_n211), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n950), .B1(new_n938), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(KEYINPUT60), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT60), .ZN(new_n954));
  OAI211_X1 g753(.A(new_n950), .B(new_n954), .C1(new_n938), .C2(new_n951), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n953), .A2(new_n955), .ZN(G1350gat));
  NAND3_X1  g755(.A1(new_n939), .A2(new_n212), .A3(new_n721), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT61), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n946), .A2(new_n721), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n958), .B1(new_n959), .B2(G190gat), .ZN(new_n960));
  AOI211_X1 g759(.A(KEYINPUT61), .B(new_n212), .C1(new_n946), .C2(new_n721), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(G1351gat));
  NOR3_X1   g761(.A1(new_n276), .A2(new_n356), .A3(new_n447), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n936), .A2(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(G197gat), .B1(new_n965), .B2(new_n662), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n918), .A2(new_n921), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n276), .A2(new_n717), .A3(new_n356), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n662), .A2(G197gat), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n966), .B1(new_n969), .B2(new_n970), .ZN(G1352gat));
  NOR2_X1   g770(.A1(new_n751), .A2(G204gat), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n936), .A2(new_n963), .A3(new_n972), .ZN(new_n973));
  XOR2_X1   g772(.A(new_n973), .B(KEYINPUT62), .Z(new_n974));
  NAND3_X1  g773(.A1(new_n967), .A2(new_n635), .A3(new_n968), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(G204gat), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n974), .A2(new_n976), .ZN(G1353gat));
  NAND3_X1  g776(.A1(new_n965), .A2(new_n299), .A3(new_n521), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n918), .A2(new_n921), .A3(new_n521), .A4(new_n968), .ZN(new_n979));
  AND3_X1   g778(.A1(new_n979), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n980));
  AOI21_X1  g779(.A(KEYINPUT63), .B1(new_n979), .B2(G211gat), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n978), .B1(new_n980), .B2(new_n981), .ZN(G1354gat));
  NAND3_X1  g781(.A1(new_n967), .A2(new_n721), .A3(new_n968), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(G218gat), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n965), .A2(new_n300), .A3(new_n721), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(new_n985), .ZN(G1355gat));
endmodule


