//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 1 1 0 1 0 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n573, new_n574,
    new_n575, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n626, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1237, new_n1238,
    new_n1239;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G217));
  OR4_X1    g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OR3_X1    g034(.A1(new_n455), .A2(KEYINPUT67), .A3(new_n459), .ZN(new_n460));
  OAI21_X1  g035(.A(KEYINPUT67), .B1(new_n455), .B2(new_n459), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OR2_X1    g046(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n471), .A2(G2105), .B1(G101), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n472), .A2(KEYINPUT3), .A3(new_n473), .ZN(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n476), .A2(G137), .A3(new_n477), .A4(new_n466), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NAND2_X1  g055(.A1(new_n476), .A2(new_n466), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(new_n477), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n477), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n481), .A2(G2105), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(G136), .B2(new_n487), .ZN(G162));
  NAND4_X1  g063(.A1(new_n476), .A2(G138), .A3(new_n477), .A4(new_n466), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n477), .A2(G138), .ZN(new_n491));
  NOR3_X1   g066(.A1(new_n469), .A2(KEYINPUT4), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n496), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n477), .A2(G114), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT69), .B1(new_n501), .B2(new_n495), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n476), .A2(G126), .A3(G2105), .A4(new_n466), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n494), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n508), .A2(G651), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(KEYINPUT6), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n508), .A2(KEYINPUT70), .A3(G651), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT5), .B(G543), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n515), .A2(G88), .ZN(new_n516));
  AND2_X1   g091(.A1(G50), .A2(G543), .ZN(new_n517));
  OAI211_X1 g092(.A(KEYINPUT71), .B(new_n514), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n517), .B1(new_n515), .B2(G88), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n511), .A2(KEYINPUT6), .ZN(new_n521));
  AND3_X1   g096(.A1(new_n508), .A2(KEYINPUT70), .A3(G651), .ZN(new_n522));
  AOI21_X1  g097(.A(KEYINPUT70), .B1(new_n508), .B2(G651), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n519), .B1(new_n520), .B2(new_n524), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n518), .B(new_n525), .C1(new_n511), .C2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  AND2_X1   g103(.A1(KEYINPUT5), .A2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(KEYINPUT5), .A2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n524), .A2(new_n531), .ZN(new_n532));
  XOR2_X1   g107(.A(KEYINPUT74), .B(G89), .Z(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT75), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g114(.A(G543), .B1(new_n514), .B2(KEYINPUT73), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT73), .ZN(new_n541));
  AOI211_X1 g116(.A(new_n541), .B(new_n509), .C1(new_n512), .C2(new_n513), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G51), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n545));
  XOR2_X1   g120(.A(new_n545), .B(KEYINPUT72), .Z(new_n546));
  NAND3_X1  g121(.A1(new_n534), .A2(KEYINPUT75), .A3(new_n536), .ZN(new_n547));
  NAND4_X1  g122(.A1(new_n539), .A2(new_n544), .A3(new_n546), .A4(new_n547), .ZN(G286));
  INV_X1    g123(.A(G286), .ZN(G168));
  NAND2_X1  g124(.A1(G77), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G64), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n531), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT76), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n511), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n554), .B1(new_n553), .B2(new_n552), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n524), .A2(new_n541), .ZN(new_n556));
  OAI211_X1 g131(.A(KEYINPUT73), .B(new_n521), .C1(new_n522), .C2(new_n523), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n556), .A2(G52), .A3(G543), .A4(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT77), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n532), .A2(G90), .ZN(new_n560));
  AND3_X1   g135(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n559), .B1(new_n558), .B2(new_n560), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n555), .B1(new_n561), .B2(new_n562), .ZN(G301));
  INV_X1    g138(.A(G301), .ZN(G171));
  AOI22_X1  g139(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n565), .A2(new_n511), .ZN(new_n566));
  INV_X1    g141(.A(G81), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n514), .A2(new_n515), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(G43), .B2(new_n543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G860), .ZN(G153));
  NAND4_X1  g146(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND4_X1  g149(.A1(G319), .A2(G483), .A3(G661), .A4(new_n574), .ZN(new_n575));
  XOR2_X1   g150(.A(new_n575), .B(KEYINPUT78), .Z(G188));
  XOR2_X1   g151(.A(KEYINPUT79), .B(G65), .Z(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(new_n515), .B1(G78), .B2(G543), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT80), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n511), .B1(new_n578), .B2(new_n579), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n580), .A2(new_n581), .B1(G91), .B2(new_n532), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n556), .A2(G543), .A3(new_n557), .ZN(new_n583));
  INV_X1    g158(.A(G53), .ZN(new_n584));
  NOR3_X1   g159(.A1(new_n583), .A2(KEYINPUT9), .A3(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT9), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(new_n543), .B2(G53), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n582), .B1(new_n585), .B2(new_n587), .ZN(G299));
  NAND2_X1  g163(.A1(new_n543), .A2(G49), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n515), .A2(G74), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n532), .A2(G87), .B1(G651), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n591), .ZN(G288));
  OAI21_X1  g167(.A(G61), .B1(new_n529), .B2(new_n530), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT81), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n593), .A2(new_n594), .B1(G73), .B2(G543), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n515), .A2(KEYINPUT81), .A3(G61), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n511), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n515), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(new_n524), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G305));
  NAND2_X1  g176(.A1(new_n532), .A2(G85), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G47), .ZN(new_n604));
  OAI221_X1 g179(.A(new_n602), .B1(new_n511), .B2(new_n603), .C1(new_n583), .C2(new_n604), .ZN(G290));
  NAND3_X1  g180(.A1(new_n514), .A2(G92), .A3(new_n515), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g183(.A1(new_n514), .A2(KEYINPUT10), .A3(G92), .A4(new_n515), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g185(.A1(new_n556), .A2(G54), .A3(G543), .A4(new_n557), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n531), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G651), .ZN(new_n615));
  AND3_X1   g190(.A1(new_n610), .A2(new_n611), .A3(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G171), .B2(new_n618), .ZN(G284));
  OAI21_X1  g195(.A(new_n619), .B1(G171), .B2(new_n618), .ZN(G321));
  NAND2_X1  g196(.A1(G286), .A2(G868), .ZN(new_n622));
  INV_X1    g197(.A(G299), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G868), .ZN(G297));
  XNOR2_X1  g199(.A(G297), .B(KEYINPUT82), .ZN(G280));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n616), .B1(new_n626), .B2(G860), .ZN(G148));
  NAND2_X1  g202(.A1(new_n616), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G868), .B2(new_n570), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g206(.A1(new_n474), .A2(new_n466), .A3(new_n468), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT83), .B(KEYINPUT12), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(KEYINPUT13), .B(G2100), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n487), .A2(G135), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n482), .A2(G123), .ZN(new_n638));
  OR2_X1    g213(.A1(G99), .A2(G2105), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n639), .B(G2104), .C1(G111), .C2(new_n477), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n637), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(G2096), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(G2096), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n636), .A2(new_n642), .A3(new_n643), .ZN(G156));
  XOR2_X1   g219(.A(G2451), .B(G2454), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(KEYINPUT14), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2430), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2435), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n652), .B2(new_n651), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n648), .B(new_n654), .Z(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(new_n658), .A3(G14), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(G401));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT84), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2072), .B(G2078), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(new_n662), .B2(new_n663), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n663), .B(KEYINPUT17), .Z(new_n668));
  INV_X1    g243(.A(new_n661), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n665), .B(new_n667), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT85), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n666), .A2(new_n663), .A3(new_n661), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT18), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n667), .A2(new_n661), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n674), .B1(new_n668), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2096), .B(G2100), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G227));
  XOR2_X1   g254(.A(G1971), .B(G1976), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  XOR2_X1   g256(.A(G1956), .B(G2474), .Z(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  AND2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT20), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n682), .A2(new_n683), .ZN(new_n687));
  NOR3_X1   g262(.A1(new_n681), .A2(new_n684), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(new_n681), .B2(new_n687), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n690), .B(new_n691), .Z(new_n692));
  XOR2_X1   g267(.A(G1991), .B(G1996), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT86), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n692), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(G229));
  NAND2_X1  g274(.A1(new_n487), .A2(G131), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n482), .A2(G119), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n477), .A2(G107), .ZN(new_n702));
  OAI21_X1  g277(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n700), .B(new_n701), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  MUX2_X1   g279(.A(G25), .B(new_n704), .S(G29), .Z(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT35), .B(G1991), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT87), .Z(new_n707));
  XOR2_X1   g282(.A(new_n705), .B(new_n707), .Z(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n709), .A2(G24), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G290), .B2(G16), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT88), .B(G1986), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n708), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n709), .A2(G23), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n589), .A2(new_n591), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n716), .B1(new_n717), .B2(new_n709), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n718), .A2(KEYINPUT89), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(KEYINPUT89), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT33), .B(G1976), .Z(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n719), .A2(new_n722), .A3(new_n720), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n709), .A2(G22), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G166), .B2(new_n709), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1971), .ZN(new_n728));
  NOR2_X1   g303(.A1(G6), .A2(G16), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n600), .B2(G16), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT32), .B(G1981), .Z(new_n731));
  XOR2_X1   g306(.A(new_n730), .B(new_n731), .Z(new_n732));
  NOR2_X1   g307(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n724), .A2(new_n725), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n715), .B1(new_n734), .B2(KEYINPUT34), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT34), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n724), .A2(new_n733), .A3(new_n736), .A4(new_n725), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(KEYINPUT36), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT36), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n735), .A2(new_n740), .A3(new_n737), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(G162), .A2(G29), .ZN(new_n743));
  OR2_X1    g318(.A1(G29), .A2(G35), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT29), .B(G2090), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G29), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G27), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G164), .B2(new_n748), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT96), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G2078), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n748), .A2(G32), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n487), .A2(G141), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n482), .A2(G129), .ZN(new_n755));
  NAND3_X1  g330(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT26), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  AOI22_X1  g334(.A1(G105), .A2(new_n474), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n754), .A2(new_n755), .A3(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n753), .B1(new_n762), .B2(new_n748), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT27), .B(G1996), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n747), .A2(new_n752), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(G5), .A2(G16), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT95), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G301), .B2(new_n709), .ZN(new_n769));
  INV_X1    g344(.A(G1961), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n709), .A2(G21), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G286), .B2(G16), .ZN(new_n773));
  INV_X1    g348(.A(G1966), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n751), .B2(G2078), .ZN(new_n776));
  NOR3_X1   g351(.A1(new_n766), .A2(new_n771), .A3(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(G4), .A2(G16), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n616), .B2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT90), .ZN(new_n780));
  INV_X1    g355(.A(G1348), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n709), .A2(G19), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n570), .B2(new_n709), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT91), .ZN(new_n785));
  INV_X1    g360(.A(G1341), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n748), .A2(G33), .ZN(new_n789));
  NAND2_X1  g364(.A1(G115), .A2(G2104), .ZN(new_n790));
  INV_X1    g365(.A(G127), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n469), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(G2105), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT93), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n477), .A2(G103), .A3(G2104), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT25), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n487), .B2(G139), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n789), .B1(new_n798), .B2(G29), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G2072), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n487), .A2(G140), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n482), .A2(G128), .ZN(new_n802));
  OR2_X1    g377(.A1(G104), .A2(G2105), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n803), .B(G2104), .C1(G116), .C2(new_n477), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT92), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n801), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(G29), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n748), .A2(G26), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT28), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(G2067), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(G34), .ZN(new_n813));
  AOI21_X1  g388(.A(G29), .B1(new_n813), .B2(KEYINPUT24), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(KEYINPUT24), .B2(new_n813), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n479), .B2(new_n748), .ZN(new_n816));
  INV_X1    g391(.A(G2084), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT30), .B(G28), .ZN(new_n820));
  OR2_X1    g395(.A1(KEYINPUT31), .A2(G11), .ZN(new_n821));
  NAND2_X1  g396(.A1(KEYINPUT31), .A2(G11), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n820), .A2(new_n748), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(new_n641), .B2(new_n748), .ZN(new_n824));
  NOR3_X1   g399(.A1(new_n818), .A2(new_n819), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n800), .A2(new_n812), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n788), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n777), .A2(new_n782), .A3(new_n787), .A4(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n773), .A2(new_n774), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT94), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n709), .A2(G20), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT23), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n623), .B2(new_n709), .ZN(new_n833));
  INV_X1    g408(.A(G1956), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n830), .B(new_n835), .C1(new_n770), .C2(new_n769), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n828), .A2(new_n836), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n742), .A2(new_n837), .ZN(G311));
  INV_X1    g413(.A(KEYINPUT97), .ZN(new_n839));
  INV_X1    g414(.A(new_n741), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n740), .B1(new_n735), .B2(new_n737), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n837), .B(new_n839), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n839), .B1(new_n742), .B2(new_n837), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(G150));
  AOI22_X1  g420(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n846), .A2(new_n511), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n556), .A2(G55), .A3(G543), .A4(new_n557), .ZN(new_n848));
  AND2_X1   g423(.A1(KEYINPUT98), .A2(G93), .ZN(new_n849));
  NOR2_X1   g424(.A1(KEYINPUT98), .A2(G93), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n532), .A2(new_n851), .ZN(new_n852));
  AND3_X1   g427(.A1(new_n848), .A2(KEYINPUT99), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(KEYINPUT99), .B1(new_n848), .B2(new_n852), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n847), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(G860), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT37), .Z(new_n857));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n626), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n855), .A2(KEYINPUT100), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n861), .B(new_n847), .C1(new_n853), .C2(new_n854), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n860), .A2(new_n570), .A3(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT38), .ZN(new_n864));
  INV_X1    g439(.A(new_n570), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n865), .A2(new_n855), .A3(KEYINPUT100), .ZN(new_n866));
  AND3_X1   g441(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n864), .B1(new_n863), .B2(new_n866), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n859), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n862), .A2(new_n570), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT99), .ZN(new_n871));
  INV_X1    g446(.A(G55), .ZN(new_n872));
  NOR3_X1   g447(.A1(new_n540), .A2(new_n542), .A3(new_n872), .ZN(new_n873));
  NOR3_X1   g448(.A1(new_n568), .A2(new_n850), .A3(new_n849), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n871), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n848), .A2(KEYINPUT99), .A3(new_n852), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n861), .B1(new_n877), .B2(new_n847), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n870), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n866), .ZN(new_n880));
  OAI21_X1  g455(.A(KEYINPUT38), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(new_n858), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n869), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT39), .ZN(new_n885));
  AOI21_X1  g460(.A(G860), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n869), .A2(KEYINPUT39), .A3(new_n883), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT101), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NOR3_X1   g463(.A1(new_n867), .A2(new_n868), .A3(new_n859), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n858), .B1(new_n881), .B2(new_n882), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n885), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(G860), .ZN(new_n892));
  AND4_X1   g467(.A1(KEYINPUT101), .A2(new_n891), .A3(new_n892), .A4(new_n887), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n857), .B1(new_n888), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(KEYINPUT102), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT102), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n896), .B(new_n857), .C1(new_n888), .C2(new_n893), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(G145));
  XNOR2_X1  g473(.A(new_n641), .B(new_n479), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n899), .B(G162), .Z(new_n900));
  XNOR2_X1  g475(.A(new_n806), .B(KEYINPUT104), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n798), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n482), .A2(G130), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n477), .A2(G118), .ZN(new_n904));
  OAI21_X1  g479(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n906), .B1(G142), .B2(new_n487), .ZN(new_n907));
  XOR2_X1   g482(.A(new_n907), .B(new_n704), .Z(new_n908));
  XNOR2_X1  g483(.A(new_n902), .B(new_n908), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n490), .A2(KEYINPUT103), .A3(new_n493), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT103), .B1(new_n490), .B2(new_n493), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n505), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(new_n762), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(new_n634), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n909), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n909), .A2(new_n914), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n900), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n917), .ZN(new_n919));
  INV_X1    g494(.A(new_n900), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(new_n920), .A3(new_n915), .ZN(new_n921));
  INV_X1    g496(.A(G37), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n918), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g499(.A(G290), .B(G305), .ZN(new_n925));
  XNOR2_X1  g500(.A(G288), .B(KEYINPUT106), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(G303), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n928));
  XNOR2_X1  g503(.A(G288), .B(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(G166), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n925), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n927), .A2(new_n930), .A3(new_n925), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XOR2_X1   g509(.A(KEYINPUT107), .B(KEYINPUT42), .Z(new_n935));
  OR2_X1    g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n933), .ZN(new_n937));
  OAI22_X1  g512(.A1(new_n937), .A2(new_n931), .B1(KEYINPUT107), .B2(KEYINPUT42), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n863), .A2(new_n866), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n939), .B(new_n628), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT105), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT9), .B1(new_n583), .B2(new_n584), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n543), .A2(new_n586), .A3(G53), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n944), .A2(new_n616), .A3(new_n582), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n608), .A2(new_n609), .B1(G651), .B2(new_n614), .ZN(new_n946));
  AOI22_X1  g521(.A1(new_n944), .A2(new_n582), .B1(new_n611), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n941), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(G299), .A2(new_n617), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n944), .A2(new_n616), .A3(new_n582), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(KEYINPUT105), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n940), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT41), .B1(new_n945), .B2(new_n947), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT41), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n949), .A2(new_n955), .A3(new_n950), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n940), .A2(new_n958), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n936), .B(new_n938), .C1(new_n953), .C2(new_n959), .ZN(new_n960));
  XOR2_X1   g535(.A(new_n939), .B(new_n628), .Z(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n957), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n938), .B1(new_n934), .B2(new_n935), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n940), .A2(new_n952), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n618), .B1(new_n960), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n855), .A2(new_n618), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT108), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n963), .B1(new_n962), .B2(new_n964), .ZN(new_n971));
  OAI21_X1  g546(.A(G868), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(new_n973), .A3(new_n967), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n969), .A2(new_n974), .ZN(G295));
  OAI21_X1  g550(.A(KEYINPUT109), .B1(new_n966), .B2(new_n968), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT109), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n972), .A2(new_n977), .A3(new_n967), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n978), .ZN(G331));
  INV_X1    g554(.A(KEYINPUT111), .ZN(new_n980));
  NAND2_X1  g555(.A1(G171), .A2(G168), .ZN(new_n981));
  NAND2_X1  g556(.A1(G301), .A2(G286), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n939), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n863), .A2(new_n866), .A3(new_n982), .A4(new_n981), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(new_n952), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n985), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT110), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n954), .A2(new_n988), .A3(new_n956), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n945), .A2(new_n947), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n990), .A2(KEYINPUT110), .A3(new_n955), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  AOI22_X1  g567(.A1(new_n980), .A2(new_n986), .B1(new_n987), .B2(new_n992), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n986), .A2(new_n980), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n934), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT43), .ZN(new_n996));
  INV_X1    g571(.A(new_n985), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n863), .A2(new_n866), .B1(new_n981), .B2(new_n982), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n957), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n984), .A2(new_n990), .A3(new_n985), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n999), .A2(new_n934), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n922), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n995), .A2(new_n996), .A3(new_n1002), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n1001), .A2(new_n922), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n999), .A2(new_n1000), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1005), .A2(new_n933), .A3(new_n932), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT43), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT44), .B1(new_n1003), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n995), .A2(KEYINPUT43), .A3(new_n1002), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n996), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1008), .A2(new_n1012), .ZN(G397));
  INV_X1    g588(.A(KEYINPUT103), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n494), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n492), .B1(new_n489), .B2(KEYINPUT4), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT103), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(G1384), .B1(new_n1018), .B2(new_n505), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT112), .B(KEYINPUT45), .Z(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n475), .A2(G40), .A3(new_n478), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT113), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n475), .A2(new_n1025), .A3(G40), .A4(new_n478), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1022), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT115), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT115), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1022), .A2(new_n1030), .A3(new_n1027), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n806), .B(G2067), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1029), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1033), .B(KEYINPUT116), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n704), .A2(new_n707), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n704), .A2(new_n707), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1035), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1029), .A2(new_n761), .A3(new_n1031), .ZN(new_n1039));
  INV_X1    g614(.A(G1996), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1022), .A2(new_n1040), .A3(new_n1027), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1042), .B1(G1996), .B2(new_n762), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1034), .A2(new_n1038), .A3(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(G290), .A2(G1986), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n1045), .B(KEYINPUT114), .ZN(new_n1046));
  NAND2_X1  g621(.A1(G290), .A2(G1986), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1028), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1044), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT122), .ZN(new_n1050));
  INV_X1    g625(.A(G1384), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT45), .B1(new_n912), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n503), .A2(new_n504), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1051), .B1(new_n1016), .B2(new_n1053), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1024), .B(new_n1026), .C1(new_n1054), .C2(new_n1020), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n774), .B1(new_n1052), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n1057));
  AOI21_X1  g632(.A(G1384), .B1(new_n494), .B2(new_n505), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT50), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1057), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1054), .A2(KEYINPUT117), .A3(KEYINPUT50), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n912), .A2(new_n1059), .A3(new_n1051), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1024), .A2(new_n1026), .A3(new_n817), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1056), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G8), .ZN(new_n1067));
  NOR2_X1   g642(.A1(G286), .A2(new_n1067), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n912), .A2(KEYINPUT45), .A3(new_n1051), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1054), .A2(new_n1020), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n1027), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G1971), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  XOR2_X1   g649(.A(KEYINPUT118), .B(G2090), .Z(new_n1075));
  NAND4_X1  g650(.A1(new_n1062), .A2(new_n1027), .A3(new_n1063), .A4(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1067), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(G303), .A2(G8), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT55), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1069), .B(KEYINPUT63), .C1(new_n1077), .C2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1067), .B1(new_n1019), .B2(new_n1027), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n717), .A2(G1976), .ZN(new_n1086));
  INV_X1    g661(.A(G1976), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT52), .B1(G288), .B2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .A4(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT49), .ZN(new_n1090));
  INV_X1    g665(.A(G1981), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n595), .A2(new_n596), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(G651), .ZN(new_n1093));
  INV_X1    g668(.A(new_n599), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1091), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n597), .A2(G1981), .A3(new_n599), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1090), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT121), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT121), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1099), .B(new_n1090), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  OR3_X1    g676(.A1(new_n1095), .A2(new_n1096), .A3(new_n1090), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1101), .A2(new_n1084), .A3(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n912), .A2(new_n1051), .A3(new_n1024), .A4(new_n1026), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1104), .A2(G8), .A3(new_n1086), .A4(new_n1088), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT120), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1104), .A2(G8), .A3(new_n1086), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT52), .ZN(new_n1108));
  AND4_X1   g683(.A1(new_n1089), .A2(new_n1103), .A3(new_n1106), .A4(new_n1108), .ZN(new_n1109));
  AND3_X1   g684(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT119), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1080), .A2(new_n1113), .A3(new_n1081), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1077), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1109), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1050), .B1(new_n1083), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1119));
  AOI211_X1 g694(.A(new_n1067), .B(new_n1119), .C1(new_n1074), .C2(new_n1076), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1089), .A2(new_n1103), .A3(new_n1106), .A4(new_n1108), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1069), .A2(KEYINPUT63), .ZN(new_n1123));
  OR2_X1    g698(.A1(new_n1077), .A2(new_n1082), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1122), .A2(new_n1123), .A3(KEYINPUT122), .A4(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1082), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1059), .B1(new_n912), .B2(new_n1051), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1024), .B(new_n1026), .C1(KEYINPUT50), .C2(new_n1054), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1129), .A2(new_n1075), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1126), .B1(new_n1130), .B2(new_n1067), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1109), .A2(new_n1131), .A3(new_n1116), .A4(new_n1069), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT63), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1118), .A2(new_n1125), .A3(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1056), .A2(new_n1065), .A3(G168), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(G8), .ZN(new_n1137));
  AOI21_X1  g712(.A(G168), .B1(new_n1056), .B2(new_n1065), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT51), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT51), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1136), .A2(new_n1140), .A3(G8), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT62), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1139), .A2(new_n1144), .A3(new_n1141), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1062), .A2(new_n1027), .A3(new_n1063), .ZN(new_n1146));
  INV_X1    g721(.A(G2078), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1070), .A2(new_n1147), .A3(new_n1027), .A4(new_n1071), .ZN(new_n1148));
  XOR2_X1   g723(.A(KEYINPUT125), .B(KEYINPUT53), .Z(new_n1149));
  AOI22_X1  g724(.A1(new_n770), .A2(new_n1146), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1147), .A2(KEYINPUT53), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(G301), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1154));
  AND4_X1   g729(.A1(new_n1154), .A2(new_n1109), .A3(new_n1131), .A4(new_n1116), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1143), .A2(new_n1145), .A3(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1103), .A2(new_n1087), .A3(new_n717), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(G1981), .B2(G305), .ZN(new_n1158));
  AOI22_X1  g733(.A1(new_n1158), .A2(new_n1084), .B1(new_n1109), .B2(new_n1120), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1135), .A2(new_n1156), .A3(new_n1159), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1109), .A2(new_n1131), .A3(new_n1116), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT54), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1146), .A2(new_n770), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1023), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1165), .A2(new_n1152), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1070), .B(new_n1166), .C1(new_n1019), .C2(new_n1021), .ZN(new_n1167));
  AND4_X1   g742(.A1(G301), .A2(new_n1163), .A3(new_n1164), .A4(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1162), .B1(new_n1154), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1163), .A2(new_n1164), .A3(new_n1167), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(G171), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1150), .A2(G301), .A3(new_n1153), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1171), .A2(new_n1172), .A3(KEYINPUT54), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1161), .A2(new_n1169), .A3(new_n1142), .A4(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n834), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT57), .ZN(new_n1176));
  AND3_X1   g751(.A1(new_n944), .A2(new_n1176), .A3(new_n582), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1176), .B1(new_n944), .B2(new_n582), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(KEYINPUT56), .B(G2072), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1070), .A2(new_n1027), .A3(new_n1071), .A4(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1175), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  AND2_X1   g757(.A1(new_n1175), .A2(new_n1181), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1178), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT123), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n944), .A2(new_n1176), .A3(new_n582), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(KEYINPUT123), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  OAI211_X1 g764(.A(KEYINPUT61), .B(new_n1182), .C1(new_n1183), .C2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1104), .A2(G2067), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1191), .B1(new_n1146), .B2(new_n781), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1192), .A2(KEYINPUT60), .A3(new_n617), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1070), .A2(new_n1040), .A3(new_n1027), .A4(new_n1071), .ZN(new_n1194));
  XOR2_X1   g769(.A(KEYINPUT58), .B(G1341), .Z(new_n1195));
  NAND2_X1  g770(.A1(new_n1104), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n865), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1197));
  OR2_X1    g772(.A1(new_n1197), .A2(KEYINPUT59), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1197), .A2(KEYINPUT59), .ZN(new_n1199));
  AND4_X1   g774(.A1(new_n1190), .A2(new_n1193), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT61), .ZN(new_n1201));
  AND3_X1   g776(.A1(new_n1175), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1179), .B1(new_n1175), .B2(new_n1181), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1201), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1204), .A2(KEYINPUT124), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT124), .ZN(new_n1206));
  OAI211_X1 g781(.A(new_n1206), .B(new_n1201), .C1(new_n1202), .C2(new_n1203), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n617), .B1(new_n1192), .B2(KEYINPUT60), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1209), .B1(KEYINPUT60), .B2(new_n1192), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1200), .A2(new_n1208), .A3(new_n1210), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1183), .A2(new_n1189), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n1192), .A2(new_n617), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1212), .B1(new_n1182), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1174), .B1(new_n1211), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1049), .B1(new_n1160), .B2(new_n1215), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n1046), .A2(new_n1028), .ZN(new_n1217));
  XOR2_X1   g792(.A(new_n1217), .B(KEYINPUT48), .Z(new_n1218));
  NAND4_X1  g793(.A1(new_n1034), .A2(new_n1043), .A3(new_n1218), .A4(new_n1038), .ZN(new_n1219));
  INV_X1    g794(.A(KEYINPUT47), .ZN(new_n1220));
  INV_X1    g795(.A(KEYINPUT126), .ZN(new_n1221));
  OAI211_X1 g796(.A(new_n1035), .B(new_n1221), .C1(new_n761), .C2(new_n1032), .ZN(new_n1222));
  NAND3_X1  g797(.A1(new_n1039), .A2(new_n1033), .A3(KEYINPUT126), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  XOR2_X1   g799(.A(new_n1041), .B(KEYINPUT46), .Z(new_n1225));
  INV_X1    g800(.A(new_n1225), .ZN(new_n1226));
  AOI21_X1  g801(.A(new_n1220), .B1(new_n1224), .B2(new_n1226), .ZN(new_n1227));
  AOI211_X1 g802(.A(KEYINPUT47), .B(new_n1225), .C1(new_n1222), .C2(new_n1223), .ZN(new_n1228));
  OAI21_X1  g803(.A(new_n1219), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g804(.A(new_n1035), .ZN(new_n1230));
  NAND3_X1  g805(.A1(new_n1034), .A2(new_n1037), .A3(new_n1043), .ZN(new_n1231));
  OR2_X1    g806(.A1(new_n806), .A2(G2067), .ZN(new_n1232));
  AOI21_X1  g807(.A(new_n1230), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  NOR2_X1   g808(.A1(new_n1229), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1216), .A2(new_n1234), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g810(.A1(G227), .A2(new_n462), .ZN(new_n1237));
  XNOR2_X1  g811(.A(new_n1237), .B(KEYINPUT127), .ZN(new_n1238));
  AND4_X1   g812(.A1(new_n659), .A2(new_n697), .A3(new_n698), .A4(new_n1238), .ZN(new_n1239));
  OAI211_X1 g813(.A(new_n923), .B(new_n1239), .C1(new_n1010), .C2(new_n1011), .ZN(G225));
  INV_X1    g814(.A(G225), .ZN(G308));
endmodule


