//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0 0 1 1 1 0 1 1 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 0 1 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1007, new_n1008, new_n1009, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047;
  INV_X1    g000(.A(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G217), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT71), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XOR2_X1   g004(.A(KEYINPUT24), .B(G110), .Z(new_n191));
  INV_X1    g005(.A(KEYINPUT73), .ZN(new_n192));
  XNOR2_X1  g006(.A(G119), .B(G128), .ZN(new_n193));
  OR3_X1    g007(.A1(new_n191), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n192), .B1(new_n191), .B2(new_n193), .ZN(new_n195));
  INV_X1    g009(.A(G119), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G128), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT23), .B1(new_n197), .B2(KEYINPUT72), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT72), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n199), .B(new_n200), .C1(new_n196), .C2(G128), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n198), .B(new_n201), .C1(G119), .C2(new_n202), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n194), .B(new_n195), .C1(G110), .C2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G140), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G125), .ZN(new_n206));
  INV_X1    g020(.A(G125), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G140), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(new_n208), .A3(KEYINPUT16), .ZN(new_n209));
  OR3_X1    g023(.A1(new_n207), .A2(KEYINPUT16), .A3(G140), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G146), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT74), .ZN(new_n212));
  XNOR2_X1  g026(.A(new_n211), .B(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n206), .A2(new_n208), .A3(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n204), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  AOI22_X1  g030(.A1(new_n203), .A2(G110), .B1(new_n193), .B2(new_n191), .ZN(new_n217));
  AOI21_X1  g031(.A(G146), .B1(new_n209), .B2(new_n210), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n209), .A2(G146), .A3(new_n210), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n216), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G953), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(G221), .A3(G234), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n223), .B(KEYINPUT22), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n224), .B(G137), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n221), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G902), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n216), .A2(new_n220), .A3(new_n225), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n190), .B1(new_n230), .B2(KEYINPUT25), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n231), .B1(KEYINPUT25), .B2(new_n230), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n189), .A2(G902), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n227), .A2(new_n229), .A3(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n234), .B(KEYINPUT75), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT11), .ZN(new_n239));
  INV_X1    g053(.A(G134), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n239), .B1(new_n240), .B2(G137), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(G137), .ZN(new_n242));
  INV_X1    g056(.A(G137), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(KEYINPUT11), .A3(G134), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n241), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G131), .ZN(new_n246));
  INV_X1    g060(.A(G131), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n241), .A2(new_n244), .A3(new_n247), .A4(new_n242), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n214), .A2(G143), .ZN(new_n252));
  INV_X1    g066(.A(G143), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G146), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(KEYINPUT0), .A2(G128), .ZN(new_n256));
  OR2_X1    g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(G143), .B(G146), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(KEYINPUT0), .A3(G128), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n246), .A2(KEYINPUT68), .A3(new_n248), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n251), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(KEYINPUT2), .A2(G113), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT65), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n266), .A2(KEYINPUT2), .A3(G113), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT2), .ZN(new_n268));
  INV_X1    g082(.A(G113), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT65), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n265), .B1(new_n267), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n196), .A2(G116), .ZN(new_n272));
  INV_X1    g086(.A(G116), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n273), .A2(KEYINPUT66), .A3(G119), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT66), .B1(new_n273), .B2(G119), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n272), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n271), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT67), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n268), .A2(new_n269), .A3(KEYINPUT65), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n266), .B1(KEYINPUT2), .B2(G113), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n279), .A2(new_n280), .B1(KEYINPUT2), .B2(G113), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n273), .A2(G119), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT66), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n283), .B1(new_n196), .B2(G116), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n273), .A2(KEYINPUT66), .A3(G119), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n282), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n277), .A2(new_n278), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n287), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n281), .A2(new_n286), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT67), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n242), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n240), .A2(G137), .ZN(new_n293));
  OAI21_X1  g107(.A(G131), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT1), .B1(new_n253), .B2(G146), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT64), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n202), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n252), .A2(KEYINPUT64), .A3(KEYINPUT1), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n259), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n300), .A2(new_n252), .A3(new_n254), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n248), .B(new_n294), .C1(new_n299), .C2(new_n302), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n264), .A2(new_n288), .A3(new_n291), .A4(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT28), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n291), .A2(new_n288), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n262), .A2(new_n249), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  AND3_X1   g124(.A1(new_n277), .A2(new_n278), .A3(new_n287), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n278), .B1(new_n277), .B2(new_n287), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n313), .A2(KEYINPUT28), .A3(new_n303), .A4(new_n264), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n306), .A2(new_n310), .A3(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n316));
  NOR2_X1   g130(.A1(G237), .A2(G953), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G210), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n316), .B(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT26), .B(G101), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n319), .B(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n315), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n321), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n304), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT30), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n309), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n264), .A2(KEYINPUT30), .A3(new_n303), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(new_n307), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT29), .B1(new_n322), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n264), .A2(new_n303), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n307), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n306), .A2(new_n314), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n321), .A2(KEYINPUT29), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n228), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n238), .B(G472), .C1(new_n330), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n328), .A2(new_n304), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT31), .B1(new_n337), .B2(new_n323), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n315), .A2(new_n323), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT31), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n328), .A2(new_n340), .A3(new_n304), .A4(new_n321), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n338), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(G472), .A2(G902), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(KEYINPUT32), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n336), .A2(new_n344), .ZN(new_n345));
  OR2_X1    g159(.A1(new_n333), .A2(new_n334), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n315), .A2(new_n321), .B1(new_n328), .B2(new_n324), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n346), .B(new_n228), .C1(new_n347), .C2(KEYINPUT29), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n238), .B1(new_n348), .B2(G472), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT32), .B1(new_n342), .B2(new_n343), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n237), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT9), .B(G234), .ZN(new_n354));
  OAI21_X1  g168(.A(G221), .B1(new_n354), .B2(G902), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT79), .ZN(new_n357));
  INV_X1    g171(.A(G104), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT3), .B1(new_n358), .B2(G107), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT3), .ZN(new_n360));
  INV_X1    g174(.A(G107), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n361), .A3(G104), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n358), .A2(G107), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n359), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G101), .ZN(new_n365));
  INV_X1    g179(.A(G101), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n359), .A2(new_n362), .A3(new_n366), .A4(new_n363), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n365), .A2(KEYINPUT4), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT4), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n364), .A2(new_n369), .A3(G101), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n262), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n295), .A2(new_n296), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(G128), .A3(new_n298), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n255), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n301), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n361), .A2(G104), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n363), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G101), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT76), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n366), .B1(new_n376), .B2(new_n363), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT76), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n359), .A2(new_n362), .A3(new_n363), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n380), .A2(new_n382), .B1(new_n366), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n375), .A2(new_n384), .A3(KEYINPUT10), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n202), .B1(new_n252), .B2(KEYINPUT1), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n301), .B1(new_n386), .B2(new_n259), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n381), .A2(KEYINPUT76), .ZN(new_n388));
  AOI211_X1 g202(.A(new_n379), .B(new_n366), .C1(new_n376), .C2(new_n363), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n387), .B(new_n367), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT77), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT10), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n391), .B1(new_n390), .B2(new_n392), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n371), .B(new_n385), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n251), .A2(new_n263), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n390), .B1(new_n375), .B2(new_n384), .ZN(new_n397));
  AOI21_X1  g211(.A(KEYINPUT12), .B1(new_n397), .B2(new_n396), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n249), .A2(KEYINPUT12), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n299), .A2(new_n302), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n367), .B1(new_n388), .B2(new_n389), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n399), .B1(new_n402), .B2(new_n390), .ZN(new_n403));
  OAI22_X1  g217(.A1(new_n395), .A2(new_n396), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(G110), .B(G140), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n222), .A2(G227), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n405), .B(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n251), .A2(new_n263), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT78), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n395), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n390), .A2(new_n392), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT77), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n368), .A2(new_n370), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  OAI211_X1 g231(.A(KEYINPUT10), .B(new_n367), .C1(new_n388), .C2(new_n389), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n417), .A2(new_n262), .B1(new_n419), .B2(new_n375), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n415), .A2(new_n420), .A3(KEYINPUT78), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n409), .B1(new_n411), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n415), .A2(new_n420), .A3(new_n409), .ZN(new_n423));
  INV_X1    g237(.A(new_n407), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n408), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n228), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n357), .B1(new_n427), .B2(G469), .ZN(new_n428));
  INV_X1    g242(.A(G469), .ZN(new_n429));
  AOI211_X1 g243(.A(KEYINPUT79), .B(new_n429), .C1(new_n426), .C2(new_n228), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  OR2_X1    g245(.A1(new_n398), .A2(new_n403), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n432), .A2(new_n423), .A3(new_n424), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n393), .A2(new_n394), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n385), .A2(new_n371), .ZN(new_n436));
  NOR3_X1   g250(.A1(new_n435), .A2(new_n410), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT78), .B1(new_n415), .B2(new_n420), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n396), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n424), .B1(new_n439), .B2(new_n423), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT80), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n434), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n395), .A2(new_n396), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n441), .B(new_n407), .C1(new_n422), .C2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n429), .B(new_n228), .C1(new_n442), .C2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n356), .B1(new_n431), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G237), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(new_n222), .A3(G214), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT88), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n450), .A2(G143), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n253), .A2(KEYINPUT88), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(G214), .A3(new_n317), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(KEYINPUT18), .A2(G131), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(KEYINPUT89), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT89), .ZN(new_n459));
  AOI211_X1 g273(.A(new_n459), .B(new_n456), .C1(new_n452), .C2(new_n454), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT90), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n206), .A2(new_n208), .A3(new_n214), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n214), .B1(new_n206), .B2(new_n208), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n207), .A2(G140), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n205), .A2(G125), .ZN(new_n467));
  OAI21_X1  g281(.A(G146), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n468), .A2(KEYINPUT90), .A3(new_n215), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n452), .A2(new_n454), .A3(new_n456), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n465), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT91), .B1(new_n461), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n455), .A2(new_n457), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n459), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n455), .A2(KEYINPUT89), .A3(new_n457), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n465), .A2(new_n469), .A3(new_n470), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT91), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n472), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT92), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n481), .B1(new_n455), .B2(G131), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n455), .A2(G131), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n452), .A2(new_n454), .A3(KEYINPUT92), .A4(new_n247), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n206), .A2(new_n208), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(KEYINPUT19), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n213), .B(new_n485), .C1(G146), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n480), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(G113), .B(G122), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(new_n358), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT93), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n494), .B1(new_n219), .B2(new_n218), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n209), .A2(new_n210), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n214), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(KEYINPUT93), .A3(new_n211), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n455), .A2(KEYINPUT17), .A3(G131), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n495), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT94), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n495), .A2(new_n498), .A3(KEYINPUT94), .A4(new_n499), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT17), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n502), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(new_n491), .A3(new_n480), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n493), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT20), .ZN(new_n510));
  NOR2_X1   g324(.A1(G475), .A2(G902), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  XOR2_X1   g326(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n513));
  INV_X1    g327(.A(new_n511), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n514), .B1(new_n493), .B2(new_n508), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n512), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n222), .A2(G952), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n517), .B1(new_n187), .B2(new_n448), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  AOI211_X1 g333(.A(new_n228), .B(new_n222), .C1(G234), .C2(G237), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT21), .B(G898), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n508), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n491), .B1(new_n507), .B2(new_n480), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n228), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G475), .ZN(new_n527));
  INV_X1    g341(.A(G217), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n354), .A2(new_n528), .A3(G953), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n253), .A2(G128), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n202), .A2(G143), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n532), .A3(new_n240), .ZN(new_n533));
  INV_X1    g347(.A(G122), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(G116), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n273), .A2(G122), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n535), .A2(new_n536), .A3(new_n361), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n361), .B1(new_n535), .B2(new_n536), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n533), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT13), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT95), .B1(new_n531), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT95), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n542), .A2(new_n253), .A3(KEYINPUT13), .A4(G128), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n531), .A2(new_n540), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n541), .A2(new_n543), .A3(new_n532), .A4(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n539), .B1(G134), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n531), .A2(new_n532), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(G134), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n533), .ZN(new_n549));
  INV_X1    g363(.A(new_n537), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n273), .A2(KEYINPUT14), .A3(G122), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n535), .A2(new_n536), .ZN(new_n552));
  OAI211_X1 g366(.A(G107), .B(new_n551), .C1(new_n552), .C2(KEYINPUT14), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n549), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n530), .B1(new_n546), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n545), .A2(G134), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n537), .A2(new_n538), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n533), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n549), .A2(new_n550), .A3(new_n553), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n559), .A3(new_n529), .ZN(new_n560));
  AOI21_X1  g374(.A(G902), .B1(new_n555), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT96), .ZN(new_n562));
  INV_X1    g376(.A(G478), .ZN(new_n563));
  OAI22_X1  g377(.A1(new_n561), .A2(new_n562), .B1(KEYINPUT15), .B2(new_n563), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n546), .A2(new_n554), .A3(new_n530), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n529), .B1(new_n558), .B2(new_n559), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n228), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n563), .A2(KEYINPUT15), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(KEYINPUT96), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n561), .A2(new_n562), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n564), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n516), .A2(new_n523), .A3(new_n527), .A4(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(G214), .B1(G237), .B2(G902), .ZN(new_n573));
  XNOR2_X1  g387(.A(G110), .B(G122), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(KEYINPUT81), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n416), .B1(new_n291), .B2(new_n288), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT5), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n269), .B1(new_n282), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n276), .B2(new_n577), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n287), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(new_n401), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n575), .B1(new_n576), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT81), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n574), .B(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n384), .A2(new_n287), .A3(new_n579), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n584), .B(new_n585), .C1(new_n313), .C2(new_n416), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n582), .A2(new_n586), .A3(KEYINPUT6), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n400), .A2(new_n207), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n207), .B1(new_n258), .B2(new_n260), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n222), .A2(G224), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(KEYINPUT82), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n591), .B(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT6), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n595), .B(new_n575), .C1(new_n576), .C2(new_n581), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n587), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(G210), .B1(G237), .B2(G902), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT8), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n584), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n575), .A2(KEYINPUT8), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n580), .A2(new_n401), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n602), .B1(new_n585), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT7), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n592), .B1(KEYINPUT83), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n606), .B1(KEYINPUT83), .B2(new_n605), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n607), .B1(new_n588), .B2(new_n590), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT84), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n605), .B1(new_n592), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n610), .B1(new_n609), .B2(new_n592), .ZN(new_n611));
  AOI211_X1 g425(.A(new_n611), .B(new_n589), .C1(new_n400), .C2(new_n207), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n604), .A2(new_n608), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(G902), .B1(new_n613), .B2(new_n586), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n597), .A2(new_n598), .A3(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(new_n598), .B(KEYINPUT85), .Z(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n597), .B2(new_n614), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n573), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT86), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT86), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n621), .B(new_n573), .C1(new_n615), .C2(new_n618), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n572), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n353), .A2(new_n447), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G101), .ZN(G3));
  NAND2_X1  g439(.A1(new_n342), .A2(new_n228), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(G472), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n342), .A2(new_n343), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n627), .A2(new_n236), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n407), .B1(new_n422), .B2(new_n443), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n433), .B1(new_n630), .B2(KEYINPUT80), .ZN(new_n631));
  AOI211_X1 g445(.A(G469), .B(G902), .C1(new_n631), .C2(new_n444), .ZN(new_n632));
  INV_X1    g446(.A(new_n425), .ZN(new_n633));
  AOI22_X1  g447(.A1(new_n439), .A2(new_n633), .B1(new_n407), .B2(new_n404), .ZN(new_n634));
  OAI21_X1  g448(.A(G469), .B1(new_n634), .B2(G902), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(KEYINPUT79), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n429), .B1(new_n426), .B2(new_n228), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n357), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n629), .B(new_n355), .C1(new_n632), .C2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n598), .B1(new_n597), .B2(new_n614), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n573), .B1(new_n615), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n523), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n567), .A2(new_n563), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT97), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n555), .A2(new_n560), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT33), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n649), .A2(G478), .A3(new_n228), .ZN(new_n650));
  AOI22_X1  g464(.A1(new_n516), .A2(new_n527), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n645), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n641), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT34), .B(G104), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G6));
  INV_X1    g470(.A(new_n513), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n491), .B1(new_n480), .B2(new_n488), .ZN(new_n658));
  AOI22_X1  g472(.A1(new_n500), .A2(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n659));
  AOI22_X1  g473(.A1(new_n659), .A2(new_n503), .B1(new_n479), .B2(new_n472), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n658), .B1(new_n660), .B2(new_n491), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n657), .B1(new_n661), .B2(new_n514), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n515), .A2(new_n513), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n662), .A2(KEYINPUT98), .A3(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT98), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n515), .A2(new_n665), .A3(new_n513), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n571), .B1(new_n526), .B2(G475), .ZN(new_n668));
  AND4_X1   g482(.A1(new_n523), .A2(new_n667), .A3(new_n644), .A4(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n641), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT35), .B(G107), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G9));
  NAND3_X1  g486(.A1(new_n446), .A2(new_n636), .A3(new_n638), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n221), .A2(KEYINPUT99), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n221), .A2(KEYINPUT99), .ZN(new_n676));
  OAI22_X1  g490(.A1(new_n675), .A2(new_n676), .B1(KEYINPUT36), .B2(new_n226), .ZN(new_n677));
  INV_X1    g491(.A(new_n676), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n226), .A2(KEYINPUT36), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n679), .A3(new_n674), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n233), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n232), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n627), .A2(new_n628), .A3(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n673), .A2(new_n623), .A3(new_n355), .A4(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT37), .B(G110), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G12));
  INV_X1    g501(.A(G900), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n519), .B1(new_n520), .B2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n664), .A2(new_n666), .A3(new_n668), .A4(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT100), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n683), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n694), .B1(new_n350), .B2(new_n352), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n693), .A2(new_n695), .A3(new_n447), .A4(new_n644), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G128), .ZN(G30));
  XOR2_X1   g511(.A(new_n689), .B(KEYINPUT39), .Z(new_n698));
  NAND2_X1  g512(.A1(new_n447), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(new_n699), .B(KEYINPUT40), .Z(new_n700));
  NAND2_X1  g514(.A1(new_n337), .A2(new_n321), .ZN(new_n701));
  AOI21_X1  g515(.A(G902), .B1(new_n324), .B2(new_n332), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(G472), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n352), .A2(new_n344), .A3(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(new_n705), .B(KEYINPUT101), .Z(new_n706));
  INV_X1    g520(.A(new_n618), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n597), .A2(new_n614), .A3(new_n598), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(new_n709), .B(KEYINPUT38), .Z(new_n710));
  NAND2_X1  g524(.A1(new_n516), .A2(new_n527), .ZN(new_n711));
  INV_X1    g525(.A(new_n571), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n694), .A2(new_n573), .ZN(new_n714));
  NOR4_X1   g528(.A1(new_n706), .A2(new_n710), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n700), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G143), .ZN(G45));
  NAND2_X1  g531(.A1(new_n647), .A2(new_n650), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n711), .A2(new_n718), .A3(new_n690), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n695), .A2(new_n447), .A3(new_n644), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G146), .ZN(G48));
  NAND2_X1  g536(.A1(new_n630), .A2(KEYINPUT80), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n444), .A3(new_n434), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n429), .B1(new_n724), .B2(new_n228), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n632), .A2(new_n725), .A3(new_n356), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(new_n353), .A3(new_n653), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(KEYINPUT102), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT102), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n726), .A2(new_n353), .A3(new_n729), .A4(new_n653), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(KEYINPUT41), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G113), .ZN(G15));
  NAND3_X1  g547(.A1(new_n726), .A2(new_n353), .A3(new_n669), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G116), .ZN(G18));
  OAI21_X1  g549(.A(G472), .B1(new_n330), .B2(new_n335), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(KEYINPUT70), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n737), .A2(new_n352), .A3(new_n336), .A4(new_n344), .ZN(new_n738));
  INV_X1    g552(.A(new_n572), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n738), .A2(new_n739), .A3(new_n683), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n726), .A3(new_n644), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G119), .ZN(G21));
  NAND2_X1  g556(.A1(new_n333), .A2(new_n323), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n338), .A2(new_n341), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n343), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n627), .A2(new_n236), .A3(new_n745), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n645), .A2(new_n746), .A3(new_n713), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n726), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G122), .ZN(G24));
  NOR2_X1   g563(.A1(new_n632), .A2(new_n725), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n627), .A2(new_n683), .A3(new_n745), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n719), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n750), .A2(new_n355), .A3(new_n752), .A4(new_n644), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G125), .ZN(G27));
  INV_X1    g568(.A(KEYINPUT42), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n719), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n351), .B(KEYINPUT105), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n737), .A2(new_n336), .A3(new_n344), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n756), .B(new_n236), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n446), .A2(new_n635), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT103), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n707), .A2(new_n355), .A3(new_n573), .A4(new_n708), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n760), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(G902), .B1(new_n631), .B2(new_n444), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n637), .B1(new_n765), .B2(new_n429), .ZN(new_n766));
  OAI21_X1  g580(.A(KEYINPUT103), .B1(new_n766), .B2(new_n762), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n759), .B1(new_n764), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n761), .B1(new_n760), .B2(new_n763), .ZN(new_n769));
  AOI211_X1 g583(.A(KEYINPUT103), .B(new_n762), .C1(new_n446), .C2(new_n635), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n353), .B(new_n720), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  XOR2_X1   g585(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n768), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(new_n247), .ZN(G33));
  NAND2_X1  g589(.A1(new_n738), .A2(new_n236), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n776), .B1(new_n767), .B2(new_n764), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n693), .ZN(new_n778));
  XOR2_X1   g592(.A(KEYINPUT106), .B(G134), .Z(new_n779));
  XNOR2_X1  g593(.A(new_n778), .B(new_n779), .ZN(G36));
  NAND3_X1  g594(.A1(new_n516), .A2(new_n718), .A3(new_n527), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT43), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n627), .A2(new_n628), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(new_n784), .A3(new_n683), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT44), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n573), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n709), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n785), .A2(new_n786), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n787), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n634), .A2(KEYINPUT45), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(G469), .B1(new_n634), .B2(KEYINPUT45), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(G469), .B2(G902), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT46), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(KEYINPUT107), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n797), .A2(KEYINPUT46), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n800), .A2(new_n632), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n356), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(KEYINPUT108), .A3(new_n698), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT108), .B1(new_n802), .B2(new_n698), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n792), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G137), .ZN(G39));
  XOR2_X1   g621(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n808));
  OR2_X1    g622(.A1(new_n802), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n802), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n789), .ZN(new_n812));
  NOR4_X1   g626(.A1(new_n738), .A2(new_n812), .A3(new_n719), .A4(new_n236), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n809), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT110), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G140), .ZN(G42));
  INV_X1    g630(.A(new_n726), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(new_n812), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n782), .A2(new_n518), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n236), .B1(new_n757), .B2(new_n758), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(KEYINPUT48), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n726), .A2(new_n644), .ZN(new_n824));
  INV_X1    g638(.A(new_n746), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n819), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n818), .A2(new_n706), .A3(new_n236), .A4(new_n519), .ZN(new_n827));
  OAI221_X1 g641(.A(new_n517), .B1(new_n824), .B2(new_n826), .C1(new_n827), .C2(new_n652), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT51), .ZN(new_n830));
  INV_X1    g644(.A(new_n710), .ZN(new_n831));
  NOR4_X1   g645(.A1(new_n826), .A2(new_n817), .A3(new_n573), .A4(new_n831), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n832), .A2(KEYINPUT50), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(KEYINPUT50), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n830), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n809), .A2(new_n811), .B1(new_n356), .B2(new_n750), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n826), .A2(new_n812), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n835), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n711), .A2(new_n718), .ZN(new_n840));
  OAI22_X1  g654(.A1(new_n827), .A2(new_n840), .B1(new_n820), .B2(new_n751), .ZN(new_n841));
  XOR2_X1   g655(.A(new_n841), .B(KEYINPUT118), .Z(new_n842));
  OAI21_X1  g656(.A(new_n829), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n841), .B1(new_n833), .B2(new_n834), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n836), .A2(KEYINPUT117), .A3(new_n838), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n750), .A2(new_n356), .ZN(new_n847));
  INV_X1    g661(.A(new_n811), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n802), .A2(new_n808), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n846), .B1(new_n850), .B2(new_n837), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n844), .B1(new_n845), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n843), .B1(new_n852), .B2(new_n830), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n741), .A2(new_n734), .A3(new_n748), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n855), .B1(new_n730), .B2(new_n728), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n651), .A2(new_n627), .A3(new_n745), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n858), .B1(new_n769), .B2(new_n770), .ZN(new_n859));
  INV_X1    g673(.A(new_n738), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n789), .A2(new_n667), .A3(new_n527), .A4(new_n571), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n447), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n694), .A2(new_n689), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n864), .A2(new_n865), .B1(new_n693), .B2(new_n777), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT113), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n673), .A2(new_n623), .A3(new_n355), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n685), .B1(new_n868), .B2(new_n776), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n516), .A2(new_n527), .A3(new_n571), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT112), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n718), .B1(new_n516), .B2(new_n527), .ZN(new_n872));
  OAI22_X1  g686(.A1(new_n871), .A2(new_n872), .B1(new_n651), .B2(KEYINPUT112), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n522), .B1(new_n620), .B2(new_n622), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n640), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n867), .B1(new_n869), .B2(new_n876), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n447), .B(new_n623), .C1(new_n353), .C2(new_n684), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n447), .A2(new_n873), .A3(new_n629), .A4(new_n874), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n878), .A2(KEYINPUT113), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n768), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n771), .A2(new_n773), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n856), .A2(new_n866), .A3(new_n881), .A4(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n713), .A2(new_n643), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n683), .A2(new_n356), .A3(new_n689), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n760), .A2(new_n886), .A3(new_n705), .A4(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n696), .A2(new_n721), .A3(new_n753), .A4(new_n888), .ZN(new_n889));
  XOR2_X1   g703(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n890));
  AND2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT52), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n854), .B1(new_n885), .B2(new_n894), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n741), .A2(new_n734), .A3(new_n748), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n878), .A2(KEYINPUT113), .A3(new_n879), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT113), .B1(new_n878), .B2(new_n879), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n731), .B(new_n896), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n857), .B1(new_n767), .B2(new_n764), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n673), .A2(new_n355), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n902), .A2(new_n860), .A3(new_n861), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n865), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n778), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(new_n774), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n889), .B(new_n892), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n900), .A2(new_n906), .A3(new_n907), .A4(KEYINPUT53), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n895), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT115), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT115), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n889), .B(KEYINPUT52), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n854), .B1(new_n885), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT54), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n889), .A2(new_n890), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n917), .B1(new_n892), .B2(new_n889), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n900), .A2(new_n906), .A3(KEYINPUT53), .A4(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n915), .A2(new_n916), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(KEYINPUT116), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT116), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n915), .A2(new_n919), .A3(new_n922), .A4(new_n916), .ZN(new_n923));
  AOI22_X1  g737(.A1(new_n913), .A2(KEYINPUT54), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n853), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(G952), .B2(G953), .ZN(new_n926));
  NOR4_X1   g740(.A1(new_n237), .A2(new_n781), .A3(new_n356), .A4(new_n788), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT49), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n927), .B1(new_n750), .B2(new_n928), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT111), .Z(new_n930));
  AOI21_X1  g744(.A(new_n831), .B1(new_n750), .B2(new_n928), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n930), .A2(new_n706), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n926), .A2(new_n932), .ZN(G75));
  NOR2_X1   g747(.A1(new_n222), .A2(G952), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT119), .Z(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n587), .A2(new_n596), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(new_n594), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT55), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n228), .B1(new_n915), .B2(new_n919), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(G210), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT56), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n940), .A2(new_n616), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n939), .A2(new_n942), .ZN(new_n945));
  AOI211_X1 g759(.A(new_n936), .B(new_n943), .C1(new_n944), .C2(new_n945), .ZN(G51));
  NAND2_X1  g760(.A1(new_n940), .A2(new_n796), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT121), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n915), .A2(new_n916), .A3(new_n919), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n916), .B1(new_n915), .B2(new_n919), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(G469), .A2(G902), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT57), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n724), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT120), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n949), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n955), .A2(new_n956), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n934), .B1(new_n957), .B2(new_n958), .ZN(G54));
  AND3_X1   g773(.A1(new_n940), .A2(KEYINPUT58), .A3(G475), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n960), .A2(new_n509), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n960), .A2(new_n509), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n961), .A2(new_n962), .A3(new_n934), .ZN(G60));
  AOI21_X1  g777(.A(new_n772), .B1(new_n777), .B2(new_n720), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n904), .B(new_n778), .C1(new_n964), .C2(new_n768), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n899), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(KEYINPUT53), .B1(new_n966), .B2(new_n907), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n885), .A2(new_n894), .A3(new_n854), .ZN(new_n968));
  OAI21_X1  g782(.A(KEYINPUT54), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n920), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n649), .B(KEYINPUT122), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(G478), .A2(G902), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT59), .Z(new_n974));
  NOR2_X1   g788(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(KEYINPUT123), .B1(new_n970), .B2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT123), .ZN(new_n977));
  INV_X1    g791(.A(new_n975), .ZN(new_n978));
  AOI211_X1 g792(.A(new_n977), .B(new_n978), .C1(new_n969), .C2(new_n920), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n935), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n921), .A2(new_n923), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n911), .B1(new_n895), .B2(new_n908), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n908), .A2(new_n911), .ZN(new_n983));
  OAI21_X1  g797(.A(KEYINPUT54), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n974), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n971), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(KEYINPUT124), .B1(new_n980), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n972), .B1(new_n924), .B2(new_n974), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n975), .B1(new_n950), .B2(new_n951), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n977), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n970), .A2(KEYINPUT123), .A3(new_n975), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n936), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT124), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n989), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n988), .A2(new_n995), .ZN(G63));
  NAND2_X1  g810(.A1(new_n915), .A2(new_n919), .ZN(new_n997));
  NAND2_X1  g811(.A1(G217), .A2(G902), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT60), .Z(new_n999));
  AND2_X1   g813(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n681), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n227), .A2(new_n229), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n1001), .B(new_n935), .C1(new_n1002), .C2(new_n1000), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT125), .ZN(new_n1004));
  AOI21_X1  g818(.A(KEYINPUT61), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1003), .B(new_n1005), .ZN(G66));
  NAND2_X1  g820(.A1(G224), .A2(G953), .ZN(new_n1007));
  OAI22_X1  g821(.A1(new_n899), .A2(G953), .B1(new_n521), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n937), .B1(G898), .B2(new_n222), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1008), .B(new_n1009), .Z(G69));
  NAND2_X1  g824(.A1(new_n326), .A2(new_n327), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1011), .B(new_n487), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1012), .B1(new_n688), .B2(new_n222), .ZN(new_n1013));
  NOR3_X1   g827(.A1(new_n821), .A2(new_n643), .A3(new_n713), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1014), .B1(new_n804), .B2(new_n805), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n1015), .A2(new_n884), .A3(new_n778), .A4(new_n814), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n696), .A2(new_n721), .A3(new_n753), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n806), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT126), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n806), .A2(KEYINPUT126), .A3(new_n1018), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1016), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1013), .B1(new_n1023), .B2(new_n222), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n222), .B1(G227), .B2(G900), .ZN(new_n1025));
  INV_X1    g839(.A(new_n699), .ZN(new_n1026));
  NAND4_X1  g840(.A1(new_n1026), .A2(new_n353), .A3(new_n789), .A4(new_n873), .ZN(new_n1027));
  AND2_X1   g841(.A1(new_n814), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1017), .B1(new_n700), .B2(new_n715), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT62), .ZN(new_n1030));
  OR2_X1    g844(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1032));
  NAND4_X1  g846(.A1(new_n1028), .A2(new_n806), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1012), .B1(new_n1033), .B2(new_n222), .ZN(new_n1034));
  OR3_X1    g848(.A1(new_n1024), .A2(new_n1025), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n1025), .B1(new_n1024), .B2(new_n1034), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1035), .A2(new_n1036), .ZN(G72));
  NAND2_X1  g851(.A1(G472), .A2(G902), .ZN(new_n1038));
  XOR2_X1   g852(.A(new_n1038), .B(KEYINPUT63), .Z(new_n1039));
  XOR2_X1   g853(.A(new_n1039), .B(KEYINPUT127), .Z(new_n1040));
  OAI21_X1  g854(.A(new_n1040), .B1(new_n1033), .B2(new_n899), .ZN(new_n1041));
  INV_X1    g855(.A(new_n701), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n934), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g857(.A(new_n1040), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1044), .B1(new_n1023), .B2(new_n900), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n1043), .B1(new_n1045), .B2(new_n329), .ZN(new_n1046));
  AND4_X1   g860(.A1(new_n329), .A2(new_n913), .A3(new_n701), .A4(new_n1039), .ZN(new_n1047));
  NOR2_X1   g861(.A1(new_n1046), .A2(new_n1047), .ZN(G57));
endmodule


