

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U551 ( .A1(n642), .A2(n523), .ZN(n645) );
  NAND2_X2 U552 ( .A1(n705), .A2(n704), .ZN(n752) );
  XNOR2_X2 U553 ( .A(n692), .B(KEYINPUT91), .ZN(n704) );
  AND2_X2 U554 ( .A1(n557), .A2(G2104), .ZN(n886) );
  OR2_X1 U555 ( .A1(n788), .A2(n787), .ZN(n516) );
  XOR2_X1 U556 ( .A(KEYINPUT29), .B(n741), .Z(n517) );
  INV_X1 U557 ( .A(KEYINPUT28), .ZN(n713) );
  NOR2_X1 U558 ( .A1(n788), .A2(n770), .ZN(n771) );
  NAND2_X1 U559 ( .A1(G160), .A2(G40), .ZN(n692) );
  NAND2_X1 U560 ( .A1(n789), .A2(n516), .ZN(n790) );
  NOR2_X1 U561 ( .A1(G2105), .A2(G2104), .ZN(n554) );
  NOR2_X1 U562 ( .A1(n811), .A2(n810), .ZN(n813) );
  NOR2_X1 U563 ( .A1(G651), .A2(G543), .ZN(n654) );
  NOR2_X1 U564 ( .A1(G651), .A2(n642), .ZN(n647) );
  NAND2_X1 U565 ( .A1(n654), .A2(G89), .ZN(n518) );
  XNOR2_X1 U566 ( .A(KEYINPUT4), .B(n518), .ZN(n521) );
  XOR2_X1 U567 ( .A(G543), .B(KEYINPUT0), .Z(n642) );
  INV_X1 U568 ( .A(G651), .ZN(n523) );
  NAND2_X1 U569 ( .A1(n645), .A2(G76), .ZN(n519) );
  XOR2_X1 U570 ( .A(KEYINPUT75), .B(n519), .Z(n520) );
  NAND2_X1 U571 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U572 ( .A(n522), .B(KEYINPUT5), .ZN(n530) );
  NOR2_X1 U573 ( .A1(G543), .A2(n523), .ZN(n525) );
  XNOR2_X1 U574 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n524) );
  XNOR2_X1 U575 ( .A(n525), .B(n524), .ZN(n648) );
  NAND2_X1 U576 ( .A1(G63), .A2(n648), .ZN(n527) );
  NAND2_X1 U577 ( .A1(G51), .A2(n647), .ZN(n526) );
  NAND2_X1 U578 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U579 ( .A(KEYINPUT6), .B(n528), .Z(n529) );
  NAND2_X1 U580 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U581 ( .A(n531), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U582 ( .A(G168), .B(KEYINPUT8), .Z(n532) );
  XNOR2_X1 U583 ( .A(KEYINPUT76), .B(n532), .ZN(G286) );
  XOR2_X1 U584 ( .A(G2446), .B(G2451), .Z(n534) );
  XNOR2_X1 U585 ( .A(G2454), .B(KEYINPUT105), .ZN(n533) );
  XNOR2_X1 U586 ( .A(n534), .B(n533), .ZN(n541) );
  XOR2_X1 U587 ( .A(G2438), .B(G2430), .Z(n536) );
  XNOR2_X1 U588 ( .A(G2435), .B(G2443), .ZN(n535) );
  XNOR2_X1 U589 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U590 ( .A(n537), .B(G2427), .Z(n539) );
  XNOR2_X1 U591 ( .A(G1348), .B(G1341), .ZN(n538) );
  XNOR2_X1 U592 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U593 ( .A(n541), .B(n540), .ZN(n542) );
  AND2_X1 U594 ( .A1(n542), .A2(G14), .ZN(G401) );
  NAND2_X1 U595 ( .A1(G77), .A2(n645), .ZN(n544) );
  NAND2_X1 U596 ( .A1(G90), .A2(n654), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n544), .A2(n543), .ZN(n546) );
  XOR2_X1 U598 ( .A(KEYINPUT9), .B(KEYINPUT70), .Z(n545) );
  XNOR2_X1 U599 ( .A(n546), .B(n545), .ZN(n551) );
  NAND2_X1 U600 ( .A1(G64), .A2(n648), .ZN(n548) );
  NAND2_X1 U601 ( .A1(G52), .A2(n647), .ZN(n547) );
  NAND2_X1 U602 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U603 ( .A(KEYINPUT69), .B(n549), .Z(n550) );
  NOR2_X1 U604 ( .A1(n551), .A2(n550), .ZN(G171) );
  AND2_X1 U605 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U606 ( .A(G2105), .ZN(n557) );
  NAND2_X1 U607 ( .A1(G101), .A2(n886), .ZN(n552) );
  XNOR2_X1 U608 ( .A(n552), .B(KEYINPUT23), .ZN(n553) );
  XNOR2_X1 U609 ( .A(n553), .B(KEYINPUT65), .ZN(n556) );
  XOR2_X1 U610 ( .A(KEYINPUT17), .B(n554), .Z(n887) );
  NAND2_X1 U611 ( .A1(G137), .A2(n887), .ZN(n555) );
  NAND2_X1 U612 ( .A1(n556), .A2(n555), .ZN(n561) );
  NOR2_X1 U613 ( .A1(G2104), .A2(n557), .ZN(n882) );
  NAND2_X1 U614 ( .A1(G125), .A2(n882), .ZN(n559) );
  AND2_X1 U615 ( .A1(G2105), .A2(G2104), .ZN(n883) );
  NAND2_X1 U616 ( .A1(G113), .A2(n883), .ZN(n558) );
  NAND2_X1 U617 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U618 ( .A1(n561), .A2(n560), .ZN(G160) );
  INV_X1 U619 ( .A(G132), .ZN(G219) );
  INV_X1 U620 ( .A(G82), .ZN(G220) );
  INV_X1 U621 ( .A(G120), .ZN(G236) );
  INV_X1 U622 ( .A(G69), .ZN(G235) );
  INV_X1 U623 ( .A(G57), .ZN(G237) );
  NAND2_X1 U624 ( .A1(G7), .A2(G661), .ZN(n562) );
  XNOR2_X1 U625 ( .A(n562), .B(KEYINPUT10), .ZN(n563) );
  XNOR2_X1 U626 ( .A(KEYINPUT72), .B(n563), .ZN(G223) );
  INV_X1 U627 ( .A(G223), .ZN(n831) );
  NAND2_X1 U628 ( .A1(n831), .A2(G567), .ZN(n564) );
  XOR2_X1 U629 ( .A(KEYINPUT11), .B(n564), .Z(G234) );
  NAND2_X1 U630 ( .A1(n654), .A2(G81), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(KEYINPUT12), .ZN(n567) );
  NAND2_X1 U632 ( .A1(G68), .A2(n645), .ZN(n566) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(KEYINPUT13), .ZN(n570) );
  NAND2_X1 U635 ( .A1(G43), .A2(n647), .ZN(n569) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n573) );
  NAND2_X1 U637 ( .A1(n648), .A2(G56), .ZN(n571) );
  XOR2_X1 U638 ( .A(KEYINPUT14), .B(n571), .Z(n572) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n980) );
  NAND2_X1 U640 ( .A1(n980), .A2(G860), .ZN(G153) );
  INV_X1 U641 ( .A(G171), .ZN(G301) );
  INV_X1 U642 ( .A(G868), .ZN(n666) );
  NOR2_X1 U643 ( .A1(G301), .A2(n666), .ZN(n583) );
  NAND2_X1 U644 ( .A1(n647), .A2(G54), .ZN(n580) );
  NAND2_X1 U645 ( .A1(G66), .A2(n648), .ZN(n575) );
  NAND2_X1 U646 ( .A1(G92), .A2(n654), .ZN(n574) );
  NAND2_X1 U647 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U648 ( .A1(G79), .A2(n645), .ZN(n576) );
  XNOR2_X1 U649 ( .A(KEYINPUT73), .B(n576), .ZN(n577) );
  NOR2_X1 U650 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U651 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X2 U652 ( .A(KEYINPUT15), .B(n581), .Z(n968) );
  NOR2_X1 U653 ( .A1(G868), .A2(n968), .ZN(n582) );
  NOR2_X1 U654 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U655 ( .A(KEYINPUT74), .B(n584), .ZN(G284) );
  NAND2_X1 U656 ( .A1(G65), .A2(n648), .ZN(n586) );
  NAND2_X1 U657 ( .A1(G91), .A2(n654), .ZN(n585) );
  NAND2_X1 U658 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U659 ( .A1(G78), .A2(n645), .ZN(n587) );
  XNOR2_X1 U660 ( .A(KEYINPUT71), .B(n587), .ZN(n588) );
  NOR2_X1 U661 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U662 ( .A1(n647), .A2(G53), .ZN(n590) );
  NAND2_X1 U663 ( .A1(n591), .A2(n590), .ZN(G299) );
  XNOR2_X1 U664 ( .A(KEYINPUT77), .B(G868), .ZN(n592) );
  NOR2_X1 U665 ( .A1(G286), .A2(n592), .ZN(n593) );
  XNOR2_X1 U666 ( .A(n593), .B(KEYINPUT78), .ZN(n595) );
  NOR2_X1 U667 ( .A1(G299), .A2(G868), .ZN(n594) );
  NOR2_X1 U668 ( .A1(n595), .A2(n594), .ZN(G297) );
  INV_X1 U669 ( .A(G860), .ZN(n615) );
  NAND2_X1 U670 ( .A1(n615), .A2(G559), .ZN(n596) );
  INV_X1 U671 ( .A(n968), .ZN(n613) );
  NAND2_X1 U672 ( .A1(n596), .A2(n613), .ZN(n597) );
  XNOR2_X1 U673 ( .A(n597), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U674 ( .A1(n968), .A2(n666), .ZN(n598) );
  XNOR2_X1 U675 ( .A(n598), .B(KEYINPUT79), .ZN(n599) );
  NOR2_X1 U676 ( .A1(G559), .A2(n599), .ZN(n600) );
  XNOR2_X1 U677 ( .A(n600), .B(KEYINPUT80), .ZN(n602) );
  AND2_X1 U678 ( .A1(n980), .A2(n666), .ZN(n601) );
  NOR2_X1 U679 ( .A1(n602), .A2(n601), .ZN(G282) );
  NAND2_X1 U680 ( .A1(G123), .A2(n882), .ZN(n603) );
  XOR2_X1 U681 ( .A(KEYINPUT18), .B(n603), .Z(n604) );
  XNOR2_X1 U682 ( .A(n604), .B(KEYINPUT81), .ZN(n606) );
  NAND2_X1 U683 ( .A1(G99), .A2(n886), .ZN(n605) );
  NAND2_X1 U684 ( .A1(n606), .A2(n605), .ZN(n610) );
  NAND2_X1 U685 ( .A1(G135), .A2(n887), .ZN(n608) );
  NAND2_X1 U686 ( .A1(G111), .A2(n883), .ZN(n607) );
  NAND2_X1 U687 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U688 ( .A1(n610), .A2(n609), .ZN(n926) );
  XNOR2_X1 U689 ( .A(G2096), .B(n926), .ZN(n612) );
  INV_X1 U690 ( .A(G2100), .ZN(n611) );
  NAND2_X1 U691 ( .A1(n612), .A2(n611), .ZN(G156) );
  NAND2_X1 U692 ( .A1(G559), .A2(n613), .ZN(n614) );
  XNOR2_X1 U693 ( .A(n614), .B(n980), .ZN(n663) );
  NAND2_X1 U694 ( .A1(n615), .A2(n663), .ZN(n624) );
  NAND2_X1 U695 ( .A1(G80), .A2(n645), .ZN(n616) );
  XNOR2_X1 U696 ( .A(n616), .B(KEYINPUT82), .ZN(n623) );
  NAND2_X1 U697 ( .A1(G55), .A2(n647), .ZN(n618) );
  NAND2_X1 U698 ( .A1(G93), .A2(n654), .ZN(n617) );
  NAND2_X1 U699 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U700 ( .A1(G67), .A2(n648), .ZN(n619) );
  XNOR2_X1 U701 ( .A(KEYINPUT83), .B(n619), .ZN(n620) );
  NOR2_X1 U702 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U703 ( .A1(n623), .A2(n622), .ZN(n667) );
  XNOR2_X1 U704 ( .A(n624), .B(n667), .ZN(G145) );
  NAND2_X1 U705 ( .A1(G75), .A2(n645), .ZN(n626) );
  NAND2_X1 U706 ( .A1(G88), .A2(n654), .ZN(n625) );
  NAND2_X1 U707 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U708 ( .A1(G62), .A2(n648), .ZN(n628) );
  NAND2_X1 U709 ( .A1(G50), .A2(n647), .ZN(n627) );
  NAND2_X1 U710 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U711 ( .A1(n630), .A2(n629), .ZN(G166) );
  NAND2_X1 U712 ( .A1(G61), .A2(n648), .ZN(n632) );
  NAND2_X1 U713 ( .A1(G86), .A2(n654), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n645), .A2(G73), .ZN(n633) );
  XOR2_X1 U716 ( .A(KEYINPUT2), .B(n633), .Z(n634) );
  NOR2_X1 U717 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U718 ( .A(n636), .B(KEYINPUT84), .ZN(n638) );
  NAND2_X1 U719 ( .A1(G48), .A2(n647), .ZN(n637) );
  NAND2_X1 U720 ( .A1(n638), .A2(n637), .ZN(G305) );
  NAND2_X1 U721 ( .A1(G49), .A2(n647), .ZN(n640) );
  NAND2_X1 U722 ( .A1(G74), .A2(G651), .ZN(n639) );
  NAND2_X1 U723 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U724 ( .A1(n648), .A2(n641), .ZN(n644) );
  NAND2_X1 U725 ( .A1(n642), .A2(G87), .ZN(n643) );
  NAND2_X1 U726 ( .A1(n644), .A2(n643), .ZN(G288) );
  NAND2_X1 U727 ( .A1(n645), .A2(G72), .ZN(n646) );
  XOR2_X1 U728 ( .A(KEYINPUT66), .B(n646), .Z(n653) );
  NAND2_X1 U729 ( .A1(n647), .A2(G47), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n648), .A2(G60), .ZN(n649) );
  NAND2_X1 U731 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U732 ( .A(KEYINPUT68), .B(n651), .ZN(n652) );
  NOR2_X1 U733 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U734 ( .A1(n654), .A2(G85), .ZN(n655) );
  NAND2_X1 U735 ( .A1(n656), .A2(n655), .ZN(G290) );
  XOR2_X1 U736 ( .A(KEYINPUT19), .B(KEYINPUT85), .Z(n657) );
  XNOR2_X1 U737 ( .A(n667), .B(n657), .ZN(n658) );
  XNOR2_X1 U738 ( .A(n658), .B(G305), .ZN(n659) );
  XNOR2_X1 U739 ( .A(n659), .B(G288), .ZN(n660) );
  XNOR2_X1 U740 ( .A(G166), .B(n660), .ZN(n662) );
  INV_X1 U741 ( .A(G299), .ZN(n735) );
  XNOR2_X1 U742 ( .A(G290), .B(n735), .ZN(n661) );
  XNOR2_X1 U743 ( .A(n662), .B(n661), .ZN(n903) );
  XNOR2_X1 U744 ( .A(n663), .B(n903), .ZN(n664) );
  XNOR2_X1 U745 ( .A(KEYINPUT86), .B(n664), .ZN(n665) );
  NOR2_X1 U746 ( .A1(n666), .A2(n665), .ZN(n669) );
  NOR2_X1 U747 ( .A1(G868), .A2(n667), .ZN(n668) );
  NOR2_X1 U748 ( .A1(n669), .A2(n668), .ZN(G295) );
  NAND2_X1 U749 ( .A1(G2084), .A2(G2078), .ZN(n670) );
  XOR2_X1 U750 ( .A(KEYINPUT20), .B(n670), .Z(n671) );
  NAND2_X1 U751 ( .A1(G2090), .A2(n671), .ZN(n672) );
  XNOR2_X1 U752 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U753 ( .A1(n673), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U755 ( .A1(G235), .A2(G236), .ZN(n674) );
  XNOR2_X1 U756 ( .A(n674), .B(KEYINPUT87), .ZN(n675) );
  NOR2_X1 U757 ( .A1(G237), .A2(n675), .ZN(n676) );
  XNOR2_X1 U758 ( .A(KEYINPUT88), .B(n676), .ZN(n677) );
  NAND2_X1 U759 ( .A1(n677), .A2(G108), .ZN(n835) );
  NAND2_X1 U760 ( .A1(G567), .A2(n835), .ZN(n682) );
  NOR2_X1 U761 ( .A1(G220), .A2(G219), .ZN(n678) );
  XOR2_X1 U762 ( .A(KEYINPUT22), .B(n678), .Z(n679) );
  NOR2_X1 U763 ( .A1(G218), .A2(n679), .ZN(n680) );
  NAND2_X1 U764 ( .A1(G96), .A2(n680), .ZN(n836) );
  NAND2_X1 U765 ( .A1(G2106), .A2(n836), .ZN(n681) );
  NAND2_X1 U766 ( .A1(n682), .A2(n681), .ZN(n857) );
  NAND2_X1 U767 ( .A1(G661), .A2(G483), .ZN(n683) );
  NOR2_X1 U768 ( .A1(n857), .A2(n683), .ZN(n834) );
  NAND2_X1 U769 ( .A1(n834), .A2(G36), .ZN(G176) );
  NAND2_X1 U770 ( .A1(n887), .A2(G138), .ZN(n686) );
  NAND2_X1 U771 ( .A1(G102), .A2(n886), .ZN(n684) );
  XOR2_X1 U772 ( .A(KEYINPUT89), .B(n684), .Z(n685) );
  NAND2_X1 U773 ( .A1(n686), .A2(n685), .ZN(n690) );
  NAND2_X1 U774 ( .A1(G126), .A2(n882), .ZN(n688) );
  NAND2_X1 U775 ( .A1(G114), .A2(n883), .ZN(n687) );
  NAND2_X1 U776 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U777 ( .A1(n690), .A2(n689), .ZN(G164) );
  XOR2_X1 U778 ( .A(KEYINPUT90), .B(G166), .Z(G303) );
  NOR2_X1 U779 ( .A1(G164), .A2(G1384), .ZN(n705) );
  INV_X1 U780 ( .A(n704), .ZN(n693) );
  NOR2_X1 U781 ( .A1(n705), .A2(n693), .ZN(n826) );
  XNOR2_X1 U782 ( .A(KEYINPUT37), .B(G2067), .ZN(n824) );
  NAND2_X1 U783 ( .A1(G128), .A2(n882), .ZN(n695) );
  NAND2_X1 U784 ( .A1(G116), .A2(n883), .ZN(n694) );
  NAND2_X1 U785 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U786 ( .A(n696), .B(KEYINPUT35), .ZN(n701) );
  NAND2_X1 U787 ( .A1(G104), .A2(n886), .ZN(n698) );
  NAND2_X1 U788 ( .A1(G140), .A2(n887), .ZN(n697) );
  NAND2_X1 U789 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U790 ( .A(KEYINPUT34), .B(n699), .Z(n700) );
  NAND2_X1 U791 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U792 ( .A(n702), .B(KEYINPUT36), .Z(n900) );
  OR2_X1 U793 ( .A1(n824), .A2(n900), .ZN(n703) );
  XOR2_X1 U794 ( .A(KEYINPUT92), .B(n703), .Z(n933) );
  NAND2_X1 U795 ( .A1(n826), .A2(n933), .ZN(n821) );
  INV_X1 U796 ( .A(n821), .ZN(n811) );
  XNOR2_X1 U797 ( .A(G1981), .B(G305), .ZN(n985) );
  NAND2_X1 U798 ( .A1(G8), .A2(n752), .ZN(n788) );
  INV_X2 U799 ( .A(n752), .ZN(n729) );
  OR2_X1 U800 ( .A1(n729), .A2(G1961), .ZN(n708) );
  XOR2_X1 U801 ( .A(G2078), .B(KEYINPUT25), .Z(n706) );
  XNOR2_X1 U802 ( .A(KEYINPUT95), .B(n706), .ZN(n946) );
  NAND2_X1 U803 ( .A1(n729), .A2(n946), .ZN(n707) );
  NAND2_X1 U804 ( .A1(n708), .A2(n707), .ZN(n746) );
  AND2_X1 U805 ( .A1(n746), .A2(G171), .ZN(n709) );
  XOR2_X1 U806 ( .A(KEYINPUT96), .B(n709), .Z(n742) );
  NAND2_X1 U807 ( .A1(n729), .A2(G2072), .ZN(n710) );
  XNOR2_X1 U808 ( .A(n710), .B(KEYINPUT27), .ZN(n712) );
  XNOR2_X1 U809 ( .A(G1956), .B(KEYINPUT97), .ZN(n992) );
  NOR2_X1 U810 ( .A1(n992), .A2(n729), .ZN(n711) );
  NOR2_X1 U811 ( .A1(n712), .A2(n711), .ZN(n736) );
  NOR2_X1 U812 ( .A1(n736), .A2(n735), .ZN(n714) );
  XNOR2_X1 U813 ( .A(n714), .B(n713), .ZN(n740) );
  NAND2_X1 U814 ( .A1(G1348), .A2(n752), .ZN(n716) );
  NAND2_X1 U815 ( .A1(G2067), .A2(n729), .ZN(n715) );
  NAND2_X1 U816 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U817 ( .A1(n968), .A2(n717), .ZN(n734) );
  NAND2_X1 U818 ( .A1(G1348), .A2(n968), .ZN(n967) );
  INV_X1 U819 ( .A(G1341), .ZN(n718) );
  NAND2_X1 U820 ( .A1(n967), .A2(n718), .ZN(n719) );
  NAND2_X1 U821 ( .A1(n719), .A2(n752), .ZN(n723) );
  NAND2_X1 U822 ( .A1(n729), .A2(G1996), .ZN(n721) );
  XOR2_X1 U823 ( .A(KEYINPUT26), .B(KEYINPUT98), .Z(n720) );
  XNOR2_X1 U824 ( .A(KEYINPUT64), .B(n720), .ZN(n724) );
  NAND2_X1 U825 ( .A1(n721), .A2(n724), .ZN(n722) );
  NAND2_X1 U826 ( .A1(n723), .A2(n722), .ZN(n732) );
  INV_X1 U827 ( .A(n724), .ZN(n725) );
  NAND2_X1 U828 ( .A1(G1996), .A2(n725), .ZN(n727) );
  NAND2_X1 U829 ( .A1(G2067), .A2(n968), .ZN(n726) );
  NAND2_X1 U830 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U831 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U832 ( .A1(n980), .A2(n730), .ZN(n731) );
  NOR2_X1 U833 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U834 ( .A1(n734), .A2(n733), .ZN(n738) );
  NAND2_X1 U835 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U836 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U837 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U838 ( .A1(n742), .A2(n517), .ZN(n751) );
  NOR2_X1 U839 ( .A1(G1966), .A2(n788), .ZN(n763) );
  NOR2_X1 U840 ( .A1(G2084), .A2(n752), .ZN(n760) );
  NOR2_X1 U841 ( .A1(n763), .A2(n760), .ZN(n743) );
  NAND2_X1 U842 ( .A1(G8), .A2(n743), .ZN(n744) );
  XNOR2_X1 U843 ( .A(KEYINPUT30), .B(n744), .ZN(n745) );
  NOR2_X1 U844 ( .A1(G168), .A2(n745), .ZN(n748) );
  NOR2_X1 U845 ( .A1(G171), .A2(n746), .ZN(n747) );
  NOR2_X1 U846 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U847 ( .A(KEYINPUT31), .B(n749), .Z(n750) );
  NAND2_X1 U848 ( .A1(n751), .A2(n750), .ZN(n761) );
  NAND2_X1 U849 ( .A1(n761), .A2(G286), .ZN(n757) );
  NOR2_X1 U850 ( .A1(G1971), .A2(n788), .ZN(n754) );
  NOR2_X1 U851 ( .A1(G2090), .A2(n752), .ZN(n753) );
  NOR2_X1 U852 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U853 ( .A1(n755), .A2(G303), .ZN(n756) );
  NAND2_X1 U854 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U855 ( .A1(G8), .A2(n758), .ZN(n759) );
  XNOR2_X1 U856 ( .A(n759), .B(KEYINPUT32), .ZN(n767) );
  NAND2_X1 U857 ( .A1(G8), .A2(n760), .ZN(n765) );
  XNOR2_X1 U858 ( .A(KEYINPUT99), .B(n761), .ZN(n762) );
  NOR2_X1 U859 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U860 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U861 ( .A1(n767), .A2(n766), .ZN(n783) );
  INV_X1 U862 ( .A(n783), .ZN(n769) );
  NOR2_X1 U863 ( .A1(G303), .A2(G1971), .ZN(n768) );
  NOR2_X1 U864 ( .A1(G1976), .A2(G288), .ZN(n773) );
  OR2_X1 U865 ( .A1(n768), .A2(n773), .ZN(n965) );
  NOR2_X1 U866 ( .A1(n769), .A2(n965), .ZN(n770) );
  NAND2_X1 U867 ( .A1(G1976), .A2(G288), .ZN(n971) );
  NAND2_X1 U868 ( .A1(n771), .A2(n971), .ZN(n772) );
  INV_X1 U869 ( .A(KEYINPUT33), .ZN(n776) );
  NAND2_X1 U870 ( .A1(n772), .A2(n776), .ZN(n779) );
  INV_X1 U871 ( .A(n788), .ZN(n774) );
  NAND2_X1 U872 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U873 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U874 ( .A(n777), .B(KEYINPUT100), .Z(n778) );
  NAND2_X1 U875 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U876 ( .A1(n985), .A2(n780), .ZN(n791) );
  NOR2_X1 U877 ( .A1(G2090), .A2(G303), .ZN(n781) );
  NAND2_X1 U878 ( .A1(G8), .A2(n781), .ZN(n782) );
  NAND2_X1 U879 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U880 ( .A(KEYINPUT101), .B(n784), .Z(n785) );
  NAND2_X1 U881 ( .A1(n788), .A2(n785), .ZN(n789) );
  NOR2_X1 U882 ( .A1(G1981), .A2(G305), .ZN(n786) );
  XOR2_X1 U883 ( .A(n786), .B(KEYINPUT24), .Z(n787) );
  OR2_X1 U884 ( .A1(n791), .A2(n790), .ZN(n809) );
  NAND2_X1 U885 ( .A1(G105), .A2(n886), .ZN(n792) );
  XNOR2_X1 U886 ( .A(n792), .B(KEYINPUT38), .ZN(n799) );
  NAND2_X1 U887 ( .A1(G129), .A2(n882), .ZN(n794) );
  NAND2_X1 U888 ( .A1(G141), .A2(n887), .ZN(n793) );
  NAND2_X1 U889 ( .A1(n794), .A2(n793), .ZN(n797) );
  NAND2_X1 U890 ( .A1(G117), .A2(n883), .ZN(n795) );
  XNOR2_X1 U891 ( .A(KEYINPUT93), .B(n795), .ZN(n796) );
  NOR2_X1 U892 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U893 ( .A1(n799), .A2(n798), .ZN(n896) );
  NAND2_X1 U894 ( .A1(n896), .A2(G1996), .ZN(n807) );
  NAND2_X1 U895 ( .A1(G119), .A2(n882), .ZN(n801) );
  NAND2_X1 U896 ( .A1(G131), .A2(n887), .ZN(n800) );
  NAND2_X1 U897 ( .A1(n801), .A2(n800), .ZN(n805) );
  NAND2_X1 U898 ( .A1(G95), .A2(n886), .ZN(n803) );
  NAND2_X1 U899 ( .A1(G107), .A2(n883), .ZN(n802) );
  NAND2_X1 U900 ( .A1(n803), .A2(n802), .ZN(n804) );
  OR2_X1 U901 ( .A1(n805), .A2(n804), .ZN(n868) );
  NAND2_X1 U902 ( .A1(G1991), .A2(n868), .ZN(n806) );
  NAND2_X1 U903 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U904 ( .A(n808), .B(KEYINPUT94), .ZN(n929) );
  NAND2_X1 U905 ( .A1(n826), .A2(n929), .ZN(n816) );
  NAND2_X1 U906 ( .A1(n809), .A2(n816), .ZN(n810) );
  XNOR2_X1 U907 ( .A(G1986), .B(G290), .ZN(n978) );
  NAND2_X1 U908 ( .A1(n978), .A2(n826), .ZN(n812) );
  NAND2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n829) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n896), .ZN(n916) );
  NOR2_X1 U911 ( .A1(G1991), .A2(n868), .ZN(n927) );
  NOR2_X1 U912 ( .A1(G1986), .A2(G290), .ZN(n814) );
  NOR2_X1 U913 ( .A1(n927), .A2(n814), .ZN(n815) );
  XOR2_X1 U914 ( .A(KEYINPUT102), .B(n815), .Z(n817) );
  NAND2_X1 U915 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U916 ( .A(KEYINPUT103), .B(n818), .ZN(n819) );
  NOR2_X1 U917 ( .A1(n916), .A2(n819), .ZN(n820) );
  XNOR2_X1 U918 ( .A(n820), .B(KEYINPUT39), .ZN(n822) );
  NAND2_X1 U919 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U920 ( .A(n823), .B(KEYINPUT104), .ZN(n825) );
  NAND2_X1 U921 ( .A1(n900), .A2(n824), .ZN(n936) );
  NAND2_X1 U922 ( .A1(n825), .A2(n936), .ZN(n827) );
  NAND2_X1 U923 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U924 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U925 ( .A(KEYINPUT40), .B(n830), .ZN(G329) );
  NAND2_X1 U926 ( .A1(G2106), .A2(n831), .ZN(G217) );
  AND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n832) );
  NAND2_X1 U928 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U930 ( .A1(n834), .A2(n833), .ZN(G188) );
  INV_X1 U932 ( .A(G108), .ZN(G238) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  NOR2_X1 U934 ( .A1(n836), .A2(n835), .ZN(G325) );
  INV_X1 U935 ( .A(G325), .ZN(G261) );
  XOR2_X1 U936 ( .A(G2096), .B(G2100), .Z(n838) );
  XNOR2_X1 U937 ( .A(KEYINPUT42), .B(G2678), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U939 ( .A(KEYINPUT43), .B(G2090), .Z(n840) );
  XNOR2_X1 U940 ( .A(G2067), .B(G2072), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U942 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U943 ( .A(G2084), .B(G2078), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(G227) );
  XOR2_X1 U945 ( .A(G1976), .B(G1971), .Z(n846) );
  XNOR2_X1 U946 ( .A(G1996), .B(G1991), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(n856) );
  XOR2_X1 U948 ( .A(KEYINPUT107), .B(KEYINPUT41), .Z(n848) );
  XNOR2_X1 U949 ( .A(G1981), .B(KEYINPUT109), .ZN(n847) );
  XNOR2_X1 U950 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U951 ( .A(G1961), .B(G1956), .Z(n850) );
  XNOR2_X1 U952 ( .A(G1986), .B(G1966), .ZN(n849) );
  XNOR2_X1 U953 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U954 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U955 ( .A(KEYINPUT108), .B(G2474), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U957 ( .A(n856), .B(n855), .Z(G229) );
  XOR2_X1 U958 ( .A(KEYINPUT106), .B(n857), .Z(G319) );
  NAND2_X1 U959 ( .A1(G124), .A2(n882), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n858), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U961 ( .A1(n886), .A2(G100), .ZN(n859) );
  NAND2_X1 U962 ( .A1(n860), .A2(n859), .ZN(n864) );
  NAND2_X1 U963 ( .A1(G136), .A2(n887), .ZN(n862) );
  NAND2_X1 U964 ( .A1(G112), .A2(n883), .ZN(n861) );
  NAND2_X1 U965 ( .A1(n862), .A2(n861), .ZN(n863) );
  NOR2_X1 U966 ( .A1(n864), .A2(n863), .ZN(G162) );
  XNOR2_X1 U967 ( .A(G164), .B(G160), .ZN(n865) );
  XNOR2_X1 U968 ( .A(n865), .B(n926), .ZN(n871) );
  XOR2_X1 U969 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n867) );
  XNOR2_X1 U970 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n866) );
  XNOR2_X1 U971 ( .A(n867), .B(n866), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U973 ( .A(n871), .B(n870), .Z(n899) );
  NAND2_X1 U974 ( .A1(G127), .A2(n882), .ZN(n873) );
  NAND2_X1 U975 ( .A1(G115), .A2(n883), .ZN(n872) );
  NAND2_X1 U976 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U977 ( .A(n874), .B(KEYINPUT47), .ZN(n880) );
  NAND2_X1 U978 ( .A1(n887), .A2(G139), .ZN(n875) );
  XOR2_X1 U979 ( .A(KEYINPUT111), .B(n875), .Z(n877) );
  NAND2_X1 U980 ( .A1(n886), .A2(G103), .ZN(n876) );
  NAND2_X1 U981 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U982 ( .A(KEYINPUT112), .B(n878), .Z(n879) );
  NAND2_X1 U983 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U984 ( .A(n881), .B(KEYINPUT113), .ZN(n919) );
  NAND2_X1 U985 ( .A1(G130), .A2(n882), .ZN(n885) );
  NAND2_X1 U986 ( .A1(G118), .A2(n883), .ZN(n884) );
  NAND2_X1 U987 ( .A1(n885), .A2(n884), .ZN(n893) );
  NAND2_X1 U988 ( .A1(G106), .A2(n886), .ZN(n889) );
  NAND2_X1 U989 ( .A1(G142), .A2(n887), .ZN(n888) );
  NAND2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U991 ( .A(KEYINPUT110), .B(n890), .Z(n891) );
  XNOR2_X1 U992 ( .A(KEYINPUT45), .B(n891), .ZN(n892) );
  NOR2_X1 U993 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U994 ( .A(G162), .B(n894), .Z(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n919), .B(n897), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U999 ( .A1(G37), .A2(n902), .ZN(G395) );
  XNOR2_X1 U1000 ( .A(G286), .B(n903), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(n980), .B(G171), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(n906), .B(n968), .ZN(n907) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n907), .ZN(G397) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(n908), .ZN(n909) );
  NOR2_X1 U1007 ( .A1(G401), .A2(n909), .ZN(n910) );
  NAND2_X1 U1008 ( .A1(n910), .A2(G319), .ZN(n913) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n911) );
  XOR2_X1 U1010 ( .A(KEYINPUT116), .B(n911), .Z(n912) );
  NOR2_X1 U1011 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(KEYINPUT117), .B(n914), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1014 ( .A(G2090), .B(G162), .Z(n915) );
  NOR2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(n917) );
  XOR2_X1 U1016 ( .A(KEYINPUT119), .B(n917), .Z(n918) );
  XOR2_X1 U1017 ( .A(KEYINPUT51), .B(n918), .Z(n925) );
  XOR2_X1 U1018 ( .A(G2072), .B(n919), .Z(n920) );
  XNOR2_X1 U1019 ( .A(KEYINPUT120), .B(n920), .ZN(n922) );
  XOR2_X1 U1020 ( .A(G164), .B(G2078), .Z(n921) );
  NOR2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1022 ( .A(KEYINPUT50), .B(n923), .ZN(n924) );
  NAND2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n938) );
  NOR2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n931) );
  XOR2_X1 U1025 ( .A(G160), .B(G2084), .Z(n928) );
  NOR2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1029 ( .A(n934), .B(KEYINPUT118), .ZN(n935) );
  NAND2_X1 U1030 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1031 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1032 ( .A(KEYINPUT52), .B(n939), .ZN(n941) );
  INV_X1 U1033 ( .A(KEYINPUT55), .ZN(n940) );
  NAND2_X1 U1034 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1035 ( .A1(n942), .A2(G29), .ZN(n1022) );
  XNOR2_X1 U1036 ( .A(G1996), .B(G32), .ZN(n944) );
  XNOR2_X1 U1037 ( .A(G33), .B(G2072), .ZN(n943) );
  NOR2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n951) );
  XOR2_X1 U1039 ( .A(G2067), .B(G26), .Z(n945) );
  NAND2_X1 U1040 ( .A1(n945), .A2(G28), .ZN(n949) );
  XNOR2_X1 U1041 ( .A(G27), .B(n946), .ZN(n947) );
  XNOR2_X1 U1042 ( .A(KEYINPUT121), .B(n947), .ZN(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1044 ( .A1(n951), .A2(n950), .ZN(n953) );
  XNOR2_X1 U1045 ( .A(G25), .B(G1991), .ZN(n952) );
  NOR2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1047 ( .A(KEYINPUT53), .B(n954), .Z(n957) );
  XOR2_X1 U1048 ( .A(G34), .B(KEYINPUT54), .Z(n955) );
  XNOR2_X1 U1049 ( .A(G2084), .B(n955), .ZN(n956) );
  NAND2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n959) );
  XNOR2_X1 U1051 ( .A(G35), .B(G2090), .ZN(n958) );
  NOR2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1053 ( .A(KEYINPUT55), .B(n960), .Z(n961) );
  NOR2_X1 U1054 ( .A1(G29), .A2(n961), .ZN(n962) );
  XOR2_X1 U1055 ( .A(KEYINPUT122), .B(n962), .Z(n963) );
  NAND2_X1 U1056 ( .A1(G11), .A2(n963), .ZN(n1020) );
  XNOR2_X1 U1057 ( .A(G16), .B(KEYINPUT56), .ZN(n990) );
  XNOR2_X1 U1058 ( .A(G1961), .B(G301), .ZN(n964) );
  NOR2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n976) );
  NAND2_X1 U1060 ( .A1(G303), .A2(G1971), .ZN(n966) );
  NAND2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n974) );
  XNOR2_X1 U1062 ( .A(G299), .B(G1956), .ZN(n970) );
  NOR2_X1 U1063 ( .A1(n968), .A2(G1348), .ZN(n969) );
  NOR2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n972) );
  NAND2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1067 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1069 ( .A(KEYINPUT124), .B(n979), .Z(n982) );
  XOR2_X1 U1070 ( .A(n980), .B(G1341), .Z(n981) );
  NOR2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n988) );
  XNOR2_X1 U1072 ( .A(G1966), .B(G168), .ZN(n983) );
  XNOR2_X1 U1073 ( .A(n983), .B(KEYINPUT123), .ZN(n984) );
  NOR2_X1 U1074 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1075 ( .A(KEYINPUT57), .B(n986), .Z(n987) );
  NAND2_X1 U1076 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1077 ( .A1(n990), .A2(n989), .ZN(n1018) );
  INV_X1 U1078 ( .A(G16), .ZN(n1016) );
  XNOR2_X1 U1079 ( .A(G1348), .B(KEYINPUT59), .ZN(n991) );
  XNOR2_X1 U1080 ( .A(n991), .B(G4), .ZN(n996) );
  XOR2_X1 U1081 ( .A(n992), .B(G20), .Z(n994) );
  XNOR2_X1 U1082 ( .A(G19), .B(G1341), .ZN(n993) );
  NOR2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n999) );
  XOR2_X1 U1085 ( .A(KEYINPUT125), .B(G1981), .Z(n997) );
  XNOR2_X1 U1086 ( .A(G6), .B(n997), .ZN(n998) );
  NOR2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(KEYINPUT60), .B(n1000), .ZN(n1001) );
  XNOR2_X1 U1089 ( .A(n1001), .B(KEYINPUT126), .ZN(n1011) );
  XOR2_X1 U1090 ( .A(G1966), .B(KEYINPUT127), .Z(n1002) );
  XNOR2_X1 U1091 ( .A(G21), .B(n1002), .ZN(n1009) );
  XNOR2_X1 U1092 ( .A(G1971), .B(G22), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(G23), .B(G1976), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  XOR2_X1 U1095 ( .A(G1986), .B(G24), .Z(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(KEYINPUT58), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(G5), .B(G1961), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(KEYINPUT61), .B(n1014), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1023), .Z(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

