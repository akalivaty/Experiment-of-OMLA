//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0 1 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n863,
    new_n864, new_n865, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943;
  NAND2_X1  g000(.A1(KEYINPUT0), .A2(G128), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(G143), .B(G146), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n190), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n187), .A3(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n191), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT11), .ZN(new_n201));
  INV_X1    g015(.A(G134), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G137), .ZN(new_n203));
  INV_X1    g017(.A(G137), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT11), .A3(G134), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(G137), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G131), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT65), .B(G131), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n209), .A2(new_n203), .A3(new_n205), .A4(new_n206), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n200), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n193), .A2(KEYINPUT1), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n196), .A2(new_n213), .A3(G128), .ZN(new_n214));
  INV_X1    g028(.A(G128), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n193), .B(new_n195), .C1(KEYINPUT1), .C2(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n202), .A2(G137), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n204), .A2(G134), .ZN(new_n218));
  OAI21_X1  g032(.A(G131), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n210), .A2(new_n214), .A3(new_n216), .A4(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n212), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n222));
  XNOR2_X1  g036(.A(G116), .B(G119), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT2), .B(G113), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n222), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n225), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(KEYINPUT66), .A3(new_n223), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n226), .A2(new_n228), .B1(new_n224), .B2(new_n225), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n221), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n231), .A2(KEYINPUT28), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(KEYINPUT72), .ZN(new_n233));
  AND4_X1   g047(.A1(new_n210), .A2(new_n214), .A3(new_n216), .A4(new_n219), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(new_n211), .B2(new_n200), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n229), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n221), .A2(new_n230), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT28), .ZN(new_n239));
  MUX2_X1   g053(.A(KEYINPUT72), .B(new_n233), .S(new_n239), .Z(new_n240));
  INV_X1    g054(.A(G237), .ZN(new_n241));
  INV_X1    g055(.A(G953), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(new_n242), .A3(G210), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n243), .B(G101), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n244), .B(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT29), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(G902), .B1(new_n240), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT30), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n199), .B1(new_n208), .B2(new_n210), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n251), .B1(new_n252), .B2(new_n234), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n212), .A2(KEYINPUT30), .A3(new_n220), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n230), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(new_n236), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(new_n247), .ZN(new_n257));
  INV_X1    g071(.A(new_n232), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT68), .B1(new_n235), .B2(new_n229), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n221), .A2(new_n260), .A3(new_n230), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n231), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT28), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n258), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  OR2_X1    g078(.A1(new_n264), .A2(new_n247), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n248), .B(new_n257), .C1(new_n265), .C2(KEYINPUT71), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n265), .A2(KEYINPUT71), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n250), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G472), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n255), .A2(new_n246), .A3(new_n236), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT67), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT67), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n255), .A2(new_n272), .A3(new_n246), .A4(new_n236), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n271), .A2(KEYINPUT31), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT31), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n274), .A2(new_n276), .B1(new_n247), .B2(new_n264), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT32), .ZN(new_n278));
  NOR2_X1   g092(.A1(G472), .A2(G902), .ZN(new_n279));
  XOR2_X1   g093(.A(new_n279), .B(KEYINPUT69), .Z(new_n280));
  NOR3_X1   g094(.A1(new_n277), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(KEYINPUT73), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n274), .A2(new_n276), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n264), .A2(new_n247), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT70), .ZN(new_n287));
  INV_X1    g101(.A(new_n280), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT70), .B1(new_n277), .B2(new_n280), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n281), .B1(new_n291), .B2(new_n278), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT73), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n269), .B(new_n283), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G217), .ZN(new_n295));
  INV_X1    g109(.A(G902), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n295), .B1(G234), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(G125), .B(G140), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT16), .ZN(new_n300));
  INV_X1    g114(.A(G125), .ZN(new_n301));
  OR3_X1    g115(.A1(new_n301), .A2(KEYINPUT16), .A3(G140), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n192), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT75), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n300), .A2(G146), .A3(new_n302), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  XOR2_X1   g121(.A(KEYINPUT24), .B(G110), .Z(new_n308));
  XNOR2_X1  g122(.A(G119), .B(G128), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n310), .B(KEYINPUT74), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n303), .A2(KEYINPUT75), .A3(new_n192), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT23), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n313), .B1(G119), .B2(new_n215), .ZN(new_n314));
  INV_X1    g128(.A(G119), .ZN(new_n315));
  NOR3_X1   g129(.A1(new_n315), .A2(KEYINPUT23), .A3(G128), .ZN(new_n316));
  OAI22_X1  g130(.A1(new_n314), .A2(new_n316), .B1(G119), .B2(new_n215), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G110), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n307), .A2(new_n311), .A3(new_n312), .A4(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n299), .B(KEYINPUT76), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n192), .ZN(new_n321));
  OAI22_X1  g135(.A1(new_n317), .A2(G110), .B1(new_n309), .B2(new_n308), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n306), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT22), .B(G137), .ZN(new_n325));
  AND3_X1   g139(.A1(new_n242), .A2(G221), .A3(G234), .ZN(new_n326));
  XOR2_X1   g140(.A(new_n325), .B(new_n326), .Z(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n319), .A2(new_n323), .A3(new_n327), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n296), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT25), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n331), .A2(KEYINPUT25), .A3(new_n296), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n298), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n297), .A2(G902), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n331), .B(KEYINPUT77), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n294), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(G214), .B1(G237), .B2(G902), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  XOR2_X1   g157(.A(G110), .B(G122), .Z(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(KEYINPUT8), .ZN(new_n345));
  INV_X1    g159(.A(G107), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(G104), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT3), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(new_n346), .A3(G104), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT79), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n348), .A2(new_n346), .A3(KEYINPUT79), .A4(G104), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n347), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G101), .ZN(new_n354));
  INV_X1    g168(.A(G104), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT3), .B1(new_n355), .B2(G107), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT78), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI211_X1 g172(.A(KEYINPUT78), .B(KEYINPUT3), .C1(new_n355), .C2(G107), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n353), .A2(new_n354), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT81), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT81), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n353), .A2(new_n363), .A3(new_n354), .A4(new_n360), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n355), .A2(G107), .ZN(new_n366));
  OAI21_X1  g180(.A(G101), .B1(new_n366), .B2(new_n347), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n226), .A2(new_n228), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n223), .A2(KEYINPUT5), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n315), .A2(G116), .ZN(new_n371));
  OR2_X1    g185(.A1(new_n371), .A2(KEYINPUT5), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(G113), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n368), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  OR2_X1    g188(.A1(new_n373), .A2(KEYINPUT86), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(KEYINPUT86), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n375), .A2(new_n369), .A3(new_n376), .ZN(new_n377));
  AOI211_X1 g191(.A(new_n345), .B(new_n374), .C1(new_n368), .C2(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(KEYINPUT90), .B(G224), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n242), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT7), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n214), .A2(new_n216), .ZN(new_n382));
  OR2_X1    g196(.A1(new_n382), .A2(G125), .ZN(new_n383));
  XOR2_X1   g197(.A(new_n383), .B(KEYINPUT92), .Z(new_n384));
  NAND2_X1  g198(.A1(new_n199), .A2(G125), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n385), .B(KEYINPUT89), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n381), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n383), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n388), .B1(new_n389), .B2(new_n381), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n378), .A2(new_n390), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n362), .A2(KEYINPUT4), .A3(new_n364), .ZN(new_n392));
  INV_X1    g206(.A(new_n347), .ZN(new_n393));
  AOI21_X1  g207(.A(KEYINPUT79), .B1(new_n366), .B2(new_n348), .ZN(new_n394));
  INV_X1    g208(.A(new_n352), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n359), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n346), .A2(G104), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT78), .B1(new_n398), .B2(KEYINPUT3), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(G101), .B1(new_n396), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT80), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(KEYINPUT4), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n353), .A2(new_n360), .ZN(new_n405));
  INV_X1    g219(.A(new_n403), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(G101), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n230), .B1(new_n392), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT85), .ZN(new_n410));
  INV_X1    g224(.A(new_n344), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n406), .B1(new_n405), .B2(G101), .ZN(new_n412));
  AOI211_X1 g226(.A(new_n354), .B(new_n403), .C1(new_n353), .C2(new_n360), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n362), .A2(KEYINPUT4), .A3(new_n364), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n229), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT85), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n377), .A2(new_n365), .A3(new_n367), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n410), .A2(new_n411), .A3(new_n418), .A4(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(G902), .B1(new_n391), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n419), .B1(new_n416), .B2(new_n417), .ZN(new_n422));
  AOI211_X1 g236(.A(KEYINPUT85), .B(new_n229), .C1(new_n414), .C2(new_n415), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n344), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(new_n420), .A3(KEYINPUT6), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT87), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT87), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n424), .A2(new_n420), .A3(new_n427), .A4(KEYINPUT6), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT88), .B(KEYINPUT6), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n344), .B(new_n430), .C1(new_n422), .C2(new_n423), .ZN(new_n431));
  XOR2_X1   g245(.A(new_n389), .B(new_n380), .Z(new_n432));
  AND4_X1   g246(.A1(KEYINPUT91), .A2(new_n429), .A3(new_n431), .A4(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n431), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n434), .B1(new_n426), .B2(new_n428), .ZN(new_n435));
  AOI21_X1  g249(.A(KEYINPUT91), .B1(new_n435), .B2(new_n432), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n421), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(G210), .B1(G237), .B2(G902), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n438), .B(new_n421), .C1(new_n433), .C2(new_n436), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n343), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  XOR2_X1   g256(.A(KEYINPUT84), .B(G469), .Z(new_n443));
  XNOR2_X1  g257(.A(G110), .B(G140), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n242), .A2(G227), .ZN(new_n445));
  XOR2_X1   g259(.A(new_n444), .B(new_n445), .Z(new_n446));
  OAI21_X1  g260(.A(new_n200), .B1(new_n392), .B2(new_n408), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n365), .A2(new_n382), .A3(new_n367), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT10), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n365), .A2(KEYINPUT10), .A3(new_n382), .A4(new_n367), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n447), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT83), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT83), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n447), .A2(new_n450), .A3(new_n454), .A4(new_n451), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n453), .A2(new_n211), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n211), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n447), .A2(new_n450), .A3(new_n457), .A4(new_n451), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n446), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n458), .A2(new_n446), .ZN(new_n460));
  INV_X1    g274(.A(new_n448), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n382), .B1(new_n365), .B2(new_n367), .ZN(new_n462));
  OR2_X1    g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT82), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT12), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n463), .A2(new_n464), .A3(new_n465), .A4(new_n211), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n211), .B1(new_n461), .B2(new_n462), .ZN(new_n467));
  NAND2_X1  g281(.A1(KEYINPUT82), .A2(KEYINPUT12), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n464), .A2(new_n465), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n460), .A2(new_n466), .A3(new_n470), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n296), .B(new_n443), .C1(new_n459), .C2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n466), .A2(new_n458), .A3(new_n470), .ZN(new_n473));
  INV_X1    g287(.A(new_n446), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n456), .A2(new_n460), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(new_n476), .A3(G469), .ZN(new_n477));
  INV_X1    g291(.A(G469), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(new_n296), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n472), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G221), .ZN(new_n482));
  XOR2_X1   g296(.A(KEYINPUT9), .B(G234), .Z(new_n483));
  AOI21_X1  g297(.A(new_n482), .B1(new_n483), .B2(new_n296), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT14), .ZN(new_n488));
  INV_X1    g302(.A(G116), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n488), .B1(new_n489), .B2(G122), .ZN(new_n490));
  OR2_X1    g304(.A1(new_n490), .A2(KEYINPUT97), .ZN(new_n491));
  OR2_X1    g305(.A1(new_n489), .A2(G122), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(KEYINPUT97), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n488), .A2(new_n489), .A3(G122), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n491), .A2(new_n492), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G107), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n489), .A2(G122), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n346), .ZN(new_n499));
  XNOR2_X1  g313(.A(G128), .B(G143), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n202), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n500), .A2(new_n202), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n496), .B(new_n499), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n498), .B(new_n346), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT96), .B(KEYINPUT13), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n202), .B1(new_n500), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n194), .A2(G128), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n507), .B1(new_n508), .B2(new_n506), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n505), .A2(new_n509), .A3(new_n501), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n483), .A2(G217), .A3(new_n242), .ZN(new_n512));
  XOR2_X1   g326(.A(new_n511), .B(new_n512), .Z(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n296), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT98), .ZN(new_n515));
  INV_X1    g329(.A(G478), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n514), .B(new_n515), .C1(KEYINPUT15), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n514), .A2(new_n515), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT15), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(new_n519), .A3(G478), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n514), .A2(new_n515), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(KEYINPUT99), .ZN(new_n523));
  INV_X1    g337(.A(G475), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n307), .A2(new_n312), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n241), .A2(new_n242), .A3(G214), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(new_n194), .ZN(new_n527));
  INV_X1    g341(.A(new_n209), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(KEYINPUT17), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n528), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n526), .B(G143), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n209), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n525), .B(new_n529), .C1(KEYINPUT17), .C2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n321), .B1(new_n192), .B2(new_n299), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT18), .ZN(new_n536));
  INV_X1    g350(.A(G131), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n531), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n527), .A2(KEYINPUT18), .A3(G131), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n535), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n534), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(G113), .B(G122), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(new_n355), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n534), .A2(new_n543), .A3(new_n540), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n524), .B1(new_n547), .B2(new_n296), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT20), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n533), .A2(KEYINPUT93), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT19), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n299), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n553), .B1(new_n320), .B2(new_n552), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n192), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT93), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n530), .A2(new_n532), .A3(new_n556), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n551), .A2(new_n555), .A3(new_n306), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n540), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT94), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n558), .A2(KEYINPUT94), .A3(new_n540), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(new_n544), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n546), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT95), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT95), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n563), .A2(new_n566), .A3(new_n546), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(G475), .A2(G902), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n550), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n564), .A2(new_n550), .A3(new_n569), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n549), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(G952), .ZN(new_n573));
  AOI211_X1 g387(.A(G953), .B(new_n573), .C1(G234), .C2(G237), .ZN(new_n574));
  XOR2_X1   g388(.A(KEYINPUT21), .B(G898), .Z(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  AOI211_X1 g390(.A(new_n296), .B(new_n242), .C1(G234), .C2(G237), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n574), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n523), .A2(new_n572), .A3(new_n578), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n341), .A2(new_n442), .A3(new_n487), .A4(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(G101), .ZN(G3));
  AOI211_X1 g395(.A(new_n343), .B(new_n578), .C1(new_n440), .C2(new_n441), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n514), .A2(new_n516), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n511), .B(new_n512), .ZN(new_n584));
  XOR2_X1   g398(.A(new_n584), .B(KEYINPUT33), .Z(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n296), .A2(G478), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n583), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n572), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(G472), .B1(new_n277), .B2(G902), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n291), .A2(new_n591), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n487), .A2(new_n339), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n582), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(KEYINPUT34), .B(G104), .Z(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(G6));
  INV_X1    g410(.A(new_n567), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n566), .B1(new_n563), .B2(new_n546), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n569), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n599), .A2(KEYINPUT20), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n600), .A2(new_n570), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n601), .A2(new_n548), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n582), .A2(new_n523), .A3(new_n593), .A4(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(new_n346), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT100), .B(KEYINPUT35), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G9));
  XOR2_X1   g420(.A(new_n324), .B(KEYINPUT101), .Z(new_n607));
  OR2_X1    g421(.A1(new_n328), .A2(KEYINPUT36), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n336), .B1(new_n609), .B2(new_n337), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n592), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n442), .A2(new_n487), .A3(new_n579), .A4(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT102), .B(KEYINPUT37), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G110), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n614), .B(new_n616), .ZN(G12));
  AOI21_X1  g431(.A(new_n287), .B1(new_n286), .B2(new_n288), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n277), .A2(KEYINPUT70), .A3(new_n280), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n278), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n281), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n282), .B1(new_n622), .B2(KEYINPUT73), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n610), .B1(new_n623), .B2(new_n269), .ZN(new_n624));
  INV_X1    g438(.A(new_n523), .ZN(new_n625));
  INV_X1    g439(.A(G900), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n577), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n574), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n549), .B(new_n629), .C1(new_n600), .C2(new_n570), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n442), .A2(new_n624), .A3(new_n487), .A4(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G128), .ZN(G30));
  NAND2_X1  g447(.A1(new_n440), .A2(new_n441), .ZN(new_n634));
  XOR2_X1   g448(.A(new_n634), .B(KEYINPUT38), .Z(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n572), .ZN(new_n637));
  NOR4_X1   g451(.A1(new_n625), .A2(new_n343), .A3(new_n637), .A4(new_n611), .ZN(new_n638));
  AOI22_X1  g452(.A1(new_n271), .A2(new_n273), .B1(new_n247), .B2(new_n238), .ZN(new_n639));
  OAI21_X1  g453(.A(G472), .B1(new_n639), .B2(G902), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n623), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n629), .B(KEYINPUT39), .Z(new_n643));
  NOR2_X1   g457(.A1(new_n486), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n642), .B1(KEYINPUT40), .B2(new_n645), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n636), .B(new_n646), .C1(KEYINPUT40), .C2(new_n645), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G143), .ZN(G45));
  AOI21_X1  g462(.A(new_n571), .B1(new_n599), .B2(KEYINPUT20), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n588), .B(new_n629), .C1(new_n649), .C2(new_n548), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n442), .A2(new_n624), .A3(new_n487), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G146), .ZN(G48));
  OAI21_X1  g467(.A(new_n296), .B1(new_n459), .B2(new_n471), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(G469), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n655), .A2(new_n656), .A3(new_n485), .A4(new_n472), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n655), .A2(new_n472), .ZN(new_n658));
  OAI21_X1  g472(.A(KEYINPUT103), .B1(new_n658), .B2(new_n484), .ZN(new_n659));
  AND4_X1   g473(.A1(new_n339), .A2(new_n294), .A3(new_n657), .A4(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n582), .A2(new_n660), .A3(new_n590), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT41), .B(G113), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G15));
  NAND4_X1  g477(.A1(new_n582), .A2(new_n660), .A3(new_n523), .A4(new_n602), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G116), .ZN(G18));
  AND2_X1   g479(.A1(new_n659), .A2(new_n657), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n442), .A2(new_n624), .A3(new_n579), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G119), .ZN(G21));
  INV_X1    g482(.A(new_n336), .ZN(new_n669));
  INV_X1    g483(.A(new_n338), .ZN(new_n670));
  INV_X1    g484(.A(new_n337), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(KEYINPUT104), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n284), .B1(new_n240), .B2(new_n246), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n288), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n675), .A2(new_n591), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n339), .A2(new_n677), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n673), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  AND4_X1   g493(.A1(new_n572), .A2(new_n679), .A3(new_n659), .A4(new_n657), .ZN(new_n680));
  INV_X1    g494(.A(new_n578), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n680), .A2(new_n442), .A3(new_n681), .A4(new_n523), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G122), .ZN(G24));
  NAND2_X1  g497(.A1(new_n676), .A2(new_n611), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n650), .A2(KEYINPUT105), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n572), .A2(new_n686), .A3(new_n588), .A4(new_n629), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n684), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n442), .A2(new_n666), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G125), .ZN(G27));
  NAND2_X1  g504(.A1(new_n477), .A2(KEYINPUT106), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n475), .A2(new_n692), .A3(G469), .A4(new_n476), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n691), .A2(new_n472), .A3(new_n480), .A4(new_n693), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n694), .A2(new_n485), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n440), .A2(new_n695), .A3(new_n342), .A4(new_n441), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(new_n340), .ZN(new_n697));
  AOI21_X1  g511(.A(KEYINPUT42), .B1(new_n685), .B2(new_n687), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n685), .A2(new_n687), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n673), .A2(new_n678), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n281), .B1(new_n268), .B2(G472), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n278), .B1(new_n277), .B2(new_n280), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(KEYINPUT42), .B1(new_n705), .B2(new_n696), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n699), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(new_n537), .ZN(G33));
  NAND2_X1  g522(.A1(new_n697), .A2(new_n631), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G134), .ZN(G36));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n637), .A2(new_n711), .A3(new_n588), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n637), .A2(KEYINPUT107), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n572), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n713), .A2(new_n715), .A3(new_n588), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n712), .B1(new_n716), .B2(KEYINPUT43), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n592), .A2(new_n610), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n475), .A2(KEYINPUT45), .A3(new_n476), .ZN(new_n722));
  AOI21_X1  g536(.A(KEYINPUT45), .B1(new_n475), .B2(new_n476), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n722), .A2(new_n723), .A3(new_n478), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(new_n479), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT46), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n472), .B1(new_n725), .B2(KEYINPUT46), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n485), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n643), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n721), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n634), .A2(new_n343), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n732), .B1(new_n719), .B2(new_n720), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n731), .B1(KEYINPUT108), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n734), .B1(KEYINPUT108), .B2(new_n733), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT109), .B(G137), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(KEYINPUT110), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n735), .B(new_n737), .ZN(G39));
  XNOR2_X1  g552(.A(new_n729), .B(KEYINPUT47), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n294), .A2(new_n339), .A3(new_n650), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n732), .A2(new_n740), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G140), .ZN(G42));
  NOR4_X1   g559(.A1(new_n716), .A2(new_n484), .A3(new_n343), .A4(new_n701), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n658), .A2(KEYINPUT49), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT112), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n658), .A2(KEYINPUT49), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n746), .A2(new_n749), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  OR3_X1    g566(.A1(new_n636), .A2(new_n752), .A3(new_n641), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n732), .A2(new_n666), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT119), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n641), .A2(new_n672), .A3(new_n628), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(KEYINPUT120), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n759), .A2(new_n572), .A3(new_n588), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n717), .A2(new_n574), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n762), .A2(new_n611), .A3(new_n676), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n666), .A2(new_n679), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n635), .A2(new_n761), .A3(new_n343), .A4(new_n764), .ZN(new_n765));
  OR3_X1    g579(.A1(new_n765), .A2(KEYINPUT118), .A3(KEYINPUT50), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n739), .B1(new_n485), .B2(new_n658), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n761), .A2(new_n679), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n732), .A3(new_n768), .ZN(new_n769));
  XOR2_X1   g583(.A(KEYINPUT118), .B(KEYINPUT50), .Z(new_n770));
  NAND2_X1  g584(.A1(new_n765), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n766), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n760), .A2(new_n763), .A3(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n694), .A2(new_n485), .A3(new_n610), .A4(new_n629), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n777), .B1(new_n623), .B2(new_n640), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n625), .A2(new_n637), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n442), .A3(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n632), .A2(new_n652), .A3(new_n689), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT52), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n624), .A2(new_n487), .ZN(new_n784));
  INV_X1    g598(.A(new_n522), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n630), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n440), .A2(new_n342), .A3(new_n786), .A4(new_n441), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n784), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n696), .ZN(new_n792));
  AOI22_X1  g606(.A1(new_n697), .A2(new_n631), .B1(new_n792), .B2(new_n688), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n664), .A2(new_n661), .A3(new_n667), .A4(new_n682), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n589), .B1(new_n572), .B2(new_n522), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n442), .A2(new_n681), .A3(new_n593), .A4(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n580), .A2(new_n614), .A3(new_n797), .ZN(new_n798));
  NOR4_X1   g612(.A1(new_n794), .A2(new_n795), .A3(new_n707), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n783), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n781), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n805), .B1(new_n782), .B2(new_n803), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n799), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n801), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n802), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n807), .A2(KEYINPUT115), .A3(new_n801), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n776), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT53), .B1(new_n783), .B2(new_n799), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n814), .B1(new_n794), .B2(new_n798), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n795), .A2(new_n801), .A3(new_n707), .ZN(new_n816));
  INV_X1    g630(.A(new_n798), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n817), .A2(KEYINPUT116), .A3(new_n791), .A4(new_n793), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n815), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n819), .A2(new_n806), .A3(new_n820), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n632), .A2(new_n652), .A3(new_n689), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n822), .A2(KEYINPUT52), .A3(new_n780), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n781), .A2(new_n804), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n803), .A3(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n805), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n815), .A2(new_n816), .A3(new_n818), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT117), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n813), .B1(new_n821), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n776), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n812), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n762), .A2(new_n704), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n834), .A2(KEYINPUT121), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(KEYINPUT121), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n835), .A2(KEYINPUT48), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n836), .B1(new_n835), .B2(KEYINPUT48), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n759), .A2(new_n589), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n768), .A2(new_n442), .A3(new_n666), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(G952), .A3(new_n242), .ZN(new_n841));
  NOR4_X1   g655(.A1(new_n837), .A2(new_n838), .A3(new_n839), .A4(new_n841), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n775), .A2(new_n833), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(G952), .A2(G953), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n753), .B1(new_n843), .B2(new_n844), .ZN(G75));
  NOR2_X1   g659(.A1(new_n830), .A2(new_n296), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT56), .B1(new_n846), .B2(G210), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n435), .B(new_n432), .Z(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(KEYINPUT55), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n847), .A2(new_n849), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n242), .A2(G952), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(G51));
  NAND2_X1  g667(.A1(new_n821), .A2(new_n829), .ZN(new_n854));
  INV_X1    g668(.A(new_n813), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT54), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n857), .A2(new_n831), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n479), .B(KEYINPUT57), .Z(new_n859));
  OAI22_X1  g673(.A1(new_n858), .A2(new_n859), .B1(new_n459), .B2(new_n471), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n846), .A2(new_n724), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n852), .B1(new_n860), .B2(new_n861), .ZN(G54));
  INV_X1    g676(.A(new_n852), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n846), .A2(KEYINPUT58), .A3(G475), .ZN(new_n864));
  INV_X1    g678(.A(new_n568), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n866), .B1(new_n865), .B2(new_n864), .ZN(G60));
  NAND2_X1  g681(.A1(G478), .A2(G902), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(KEYINPUT59), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n869), .B1(new_n812), .B2(new_n832), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n586), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n585), .A2(new_n869), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n857), .B2(new_n831), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT122), .B1(new_n873), .B2(new_n852), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n873), .A2(KEYINPUT122), .A3(new_n852), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(G63));
  NAND2_X1  g691(.A1(G217), .A2(G902), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT60), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n670), .B1(new_n830), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n863), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n879), .B1(new_n854), .B2(new_n855), .ZN(new_n882));
  AOI21_X1  g696(.A(KEYINPUT123), .B1(new_n882), .B2(new_n609), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT124), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT61), .ZN(new_n886));
  INV_X1    g700(.A(new_n609), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n830), .A2(new_n887), .A3(new_n879), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT123), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n884), .A2(new_n885), .A3(new_n886), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n885), .A2(new_n886), .ZN(new_n891));
  NAND2_X1  g705(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n863), .B(new_n880), .C1(new_n888), .C2(KEYINPUT123), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n888), .A2(KEYINPUT123), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n891), .B(new_n892), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n890), .A2(new_n895), .ZN(G66));
  AOI21_X1  g710(.A(new_n242), .B1(new_n575), .B2(new_n379), .ZN(new_n897));
  OR2_X1    g711(.A1(new_n795), .A2(new_n798), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n897), .B1(new_n898), .B2(new_n242), .ZN(new_n899));
  INV_X1    g713(.A(G898), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n435), .B1(new_n900), .B2(G953), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n899), .B(new_n901), .ZN(G69));
  NAND2_X1  g716(.A1(G227), .A2(G900), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n709), .A2(new_n699), .A3(new_n706), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT126), .Z(new_n905));
  NAND4_X1  g719(.A1(new_n730), .A2(new_n442), .A3(new_n779), .A4(new_n704), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n906), .A2(new_n822), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n744), .A2(new_n735), .A3(new_n905), .A4(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n242), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n626), .A2(G953), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT127), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n253), .A2(new_n254), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(new_n554), .Z(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  OAI211_X1 g729(.A(G953), .B(new_n903), .C1(new_n912), .C2(new_n915), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n911), .A2(KEYINPUT127), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n911), .A2(KEYINPUT127), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n914), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n903), .A2(G953), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n744), .A2(new_n735), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT62), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n647), .B(new_n822), .C1(KEYINPUT125), .C2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n647), .A2(new_n822), .ZN(new_n924));
  XOR2_X1   g738(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n732), .A2(new_n341), .A3(new_n644), .A4(new_n796), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n921), .A2(new_n923), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n915), .B1(new_n929), .B2(G953), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n919), .A2(new_n920), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n916), .A2(new_n931), .ZN(G72));
  NAND2_X1  g746(.A1(G472), .A2(G902), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT63), .Z(new_n934));
  OAI21_X1  g748(.A(new_n934), .B1(new_n928), .B2(new_n898), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n935), .A2(new_n246), .A3(new_n256), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n934), .B1(new_n908), .B2(new_n898), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n937), .A2(new_n247), .A3(new_n236), .A4(new_n255), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n936), .A2(new_n863), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n810), .A2(new_n811), .ZN(new_n940));
  INV_X1    g754(.A(new_n934), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n271), .A2(new_n273), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n941), .B1(new_n942), .B2(new_n257), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n939), .B1(new_n940), .B2(new_n943), .ZN(G57));
endmodule


