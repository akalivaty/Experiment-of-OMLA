//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 1 0 1 0 1 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT10), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT77), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT76), .ZN(new_n194));
  XNOR2_X1  g008(.A(G104), .B(G107), .ZN(new_n195));
  INV_X1    g009(.A(G101), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n194), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G104), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT3), .B1(new_n198), .B2(G107), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n200));
  INV_X1    g014(.A(G107), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(G104), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(G107), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n199), .A2(new_n202), .A3(new_n196), .A4(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n198), .A2(G107), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n201), .A2(G104), .ZN(new_n206));
  OAI211_X1 g020(.A(KEYINPUT76), .B(G101), .C1(new_n205), .C2(new_n206), .ZN(new_n207));
  AND3_X1   g021(.A1(new_n197), .A2(new_n204), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT1), .B1(new_n209), .B2(G146), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n209), .A2(G146), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(G143), .ZN(new_n213));
  OAI211_X1 g027(.A(G128), .B(new_n210), .C1(new_n211), .C2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(G143), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n209), .A2(G146), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n215), .B(new_n216), .C1(KEYINPUT1), .C2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n193), .B1(new_n208), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n197), .A2(new_n204), .A3(new_n207), .ZN(new_n222));
  NOR3_X1   g036(.A1(new_n222), .A2(KEYINPUT77), .A3(new_n219), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n192), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n199), .A2(new_n202), .A3(new_n203), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT4), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(G101), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT75), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT75), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n225), .A2(new_n229), .A3(new_n226), .A4(G101), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(G143), .B(G146), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(KEYINPUT0), .A3(G128), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT0), .B(G128), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n233), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n225), .A2(G101), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(KEYINPUT4), .A3(new_n204), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n231), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n219), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n214), .A2(KEYINPUT67), .A3(new_n218), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(KEYINPUT10), .A3(new_n208), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n224), .A2(new_n239), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT78), .ZN(new_n246));
  INV_X1    g060(.A(G137), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(KEYINPUT11), .A3(G134), .ZN(new_n248));
  INV_X1    g062(.A(G134), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G137), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G131), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT11), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n253), .B1(new_n249), .B2(G137), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT64), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n247), .A2(G134), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT64), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(new_n257), .A3(new_n253), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n251), .A2(new_n252), .A3(new_n255), .A4(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT65), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n257), .B1(new_n256), .B2(new_n253), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n248), .A2(new_n250), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n264), .A2(KEYINPUT65), .A3(new_n252), .A4(new_n258), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n258), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G131), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT78), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n224), .A2(new_n270), .A3(new_n239), .A4(new_n244), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n246), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n261), .A2(new_n265), .B1(G131), .B2(new_n267), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n224), .A2(new_n273), .A3(new_n239), .A4(new_n244), .ZN(new_n274));
  XNOR2_X1  g088(.A(G110), .B(G140), .ZN(new_n275));
  INV_X1    g089(.A(G227), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(G953), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n275), .B(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  OAI22_X1  g095(.A1(new_n221), .A2(new_n223), .B1(new_n220), .B2(new_n208), .ZN(new_n282));
  AOI21_X1  g096(.A(KEYINPUT12), .B1(new_n282), .B2(new_n269), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n208), .A2(new_n193), .A3(new_n220), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT77), .B1(new_n222), .B2(new_n219), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n284), .A2(new_n285), .B1(new_n219), .B2(new_n222), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT12), .ZN(new_n287));
  NOR3_X1   g101(.A1(new_n286), .A2(new_n287), .A3(new_n273), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n274), .B1(new_n283), .B2(new_n288), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n272), .A2(new_n281), .B1(new_n289), .B2(new_n278), .ZN(new_n290));
  OAI21_X1  g104(.A(G469), .B1(new_n290), .B2(G902), .ZN(new_n291));
  INV_X1    g105(.A(G469), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n279), .B1(new_n272), .B2(new_n274), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n283), .A2(new_n288), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n294), .A2(new_n280), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n292), .B(new_n190), .C1(new_n293), .C2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n191), .B1(new_n291), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT83), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n235), .A2(G125), .ZN(new_n299));
  INV_X1    g113(.A(G953), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G224), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT80), .ZN(new_n302));
  INV_X1    g116(.A(G125), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n302), .B1(new_n219), .B2(new_n303), .ZN(new_n304));
  AOI211_X1 g118(.A(KEYINPUT80), .B(G125), .C1(new_n214), .C2(new_n218), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n299), .B(new_n301), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(KEYINPUT2), .A2(G113), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT66), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT66), .B1(KEYINPUT2), .B2(G113), .ZN(new_n311));
  OAI22_X1  g125(.A1(new_n310), .A2(new_n311), .B1(KEYINPUT2), .B2(G113), .ZN(new_n312));
  INV_X1    g126(.A(G119), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G116), .ZN(new_n314));
  INV_X1    g128(.A(G116), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G119), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n314), .A2(new_n316), .A3(KEYINPUT5), .ZN(new_n318));
  OAI21_X1  g132(.A(G113), .B1(new_n314), .B2(KEYINPUT5), .ZN(new_n319));
  OAI22_X1  g133(.A1(new_n312), .A2(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(new_n222), .ZN(new_n321));
  XNOR2_X1  g135(.A(G110), .B(G122), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(KEYINPUT8), .ZN(new_n323));
  AOI22_X1  g137(.A1(new_n307), .A2(KEYINPUT7), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n312), .B(new_n317), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n231), .A2(new_n325), .A3(new_n238), .ZN(new_n326));
  OR2_X1    g140(.A1(new_n320), .A2(new_n222), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n322), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n219), .A2(new_n303), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT80), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT81), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n219), .A2(new_n302), .A3(new_n303), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT81), .B1(new_n304), .B2(new_n305), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n334), .A3(new_n299), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n301), .A2(KEYINPUT7), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n324), .A2(new_n328), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n190), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n326), .A2(new_n327), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT6), .ZN(new_n341));
  INV_X1    g155(.A(new_n322), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n328), .A2(KEYINPUT6), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n322), .B1(new_n326), .B2(new_n327), .ZN(new_n345));
  OAI211_X1 g159(.A(KEYINPUT79), .B(new_n343), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n345), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT79), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n347), .A2(new_n348), .A3(KEYINPUT6), .A4(new_n328), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n299), .B1(new_n304), .B2(new_n305), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n351), .B(new_n301), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n339), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(G210), .B1(G237), .B2(G902), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n298), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n352), .B1(new_n346), .B2(new_n349), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT82), .B1(new_n357), .B2(new_n339), .ZN(new_n358));
  INV_X1    g172(.A(new_n355), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR3_X1   g174(.A1(new_n357), .A2(KEYINPUT82), .A3(new_n339), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n356), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(G214), .B1(G237), .B2(G902), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT82), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n354), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n365), .A2(new_n298), .A3(new_n359), .A4(new_n358), .ZN(new_n366));
  XNOR2_X1  g180(.A(G113), .B(G122), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n367), .B(new_n198), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n303), .A2(KEYINPUT16), .A3(G140), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(KEYINPUT71), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(G125), .B(G140), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n369), .B1(new_n372), .B2(KEYINPUT16), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT71), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n371), .B(G146), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(G237), .A2(G953), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(G143), .A3(G214), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(G143), .B1(new_n376), .B2(G214), .ZN(new_n379));
  OAI21_X1  g193(.A(G131), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n379), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(new_n252), .A3(new_n377), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G140), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G125), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n303), .A2(G140), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT85), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT19), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n372), .A2(new_n387), .A3(KEYINPUT19), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT86), .B1(new_n392), .B2(new_n212), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT86), .ZN(new_n394));
  AOI211_X1 g208(.A(new_n394), .B(G146), .C1(new_n390), .C2(new_n391), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n375), .B(new_n383), .C1(new_n393), .C2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n381), .A2(new_n377), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT84), .ZN(new_n398));
  OAI211_X1 g212(.A(KEYINPUT18), .B(G131), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(KEYINPUT18), .A2(G131), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n381), .A2(KEYINPUT84), .A3(new_n400), .A4(new_n377), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n372), .B(new_n212), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n368), .B1(new_n396), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT17), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n380), .A2(new_n382), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n385), .A2(new_n386), .A3(KEYINPUT16), .ZN(new_n407));
  OR3_X1    g221(.A1(new_n303), .A2(KEYINPUT16), .A3(G140), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n374), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n212), .B1(new_n409), .B2(new_n370), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n397), .A2(KEYINPUT17), .A3(G131), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n406), .A2(new_n410), .A3(new_n375), .A4(new_n411), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n412), .A2(new_n368), .A3(new_n403), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n404), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(G475), .A2(G902), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT20), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT20), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n418), .B(new_n415), .C1(new_n404), .C2(new_n413), .ZN(new_n419));
  INV_X1    g233(.A(G475), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n368), .B1(new_n412), .B2(new_n403), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n190), .B1(new_n413), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n420), .B1(new_n422), .B2(KEYINPUT87), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT87), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n424), .B(new_n190), .C1(new_n413), .C2(new_n421), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n417), .A2(new_n419), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G122), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G116), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n315), .A2(G122), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n201), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n428), .A2(new_n429), .A3(new_n201), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(KEYINPUT88), .A3(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT88), .ZN(new_n434));
  INV_X1    g248(.A(new_n432), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n434), .B1(new_n435), .B2(new_n430), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n209), .A2(G128), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n217), .A2(G143), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT13), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n249), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  OR2_X1    g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n439), .A2(new_n441), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n433), .A2(new_n436), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n435), .A2(KEYINPUT89), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n315), .A2(KEYINPUT14), .A3(G122), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n428), .A2(new_n429), .ZN(new_n447));
  OAI211_X1 g261(.A(G107), .B(new_n446), .C1(new_n447), .C2(KEYINPUT14), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n439), .A2(G134), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT89), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n432), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n437), .A2(new_n438), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n249), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n450), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n449), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G217), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n188), .A2(new_n457), .A3(G953), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n444), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n433), .A2(new_n436), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n442), .A2(new_n443), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n450), .A2(new_n454), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n464), .A2(new_n452), .A3(new_n445), .A4(new_n448), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n458), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n190), .B1(new_n460), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G478), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(KEYINPUT15), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n459), .B1(new_n444), .B2(new_n456), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n463), .A2(new_n465), .A3(new_n458), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n469), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n190), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n470), .A2(KEYINPUT90), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT90), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n474), .B1(new_n473), .B2(new_n190), .ZN(new_n478));
  AOI211_X1 g292(.A(G902), .B(new_n469), .C1(new_n471), .C2(new_n472), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G952), .ZN(new_n481));
  AOI211_X1 g295(.A(G953), .B(new_n481), .C1(G234), .C2(G237), .ZN(new_n482));
  AOI211_X1 g296(.A(new_n190), .B(new_n300), .C1(G234), .C2(G237), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT21), .B(G898), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n426), .A2(new_n476), .A3(new_n480), .A4(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n362), .A2(new_n363), .A3(new_n366), .A4(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT32), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n376), .A2(G210), .ZN(new_n492));
  XOR2_X1   g306(.A(new_n492), .B(KEYINPUT27), .Z(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT26), .B(G101), .ZN(new_n494));
  XOR2_X1   g308(.A(new_n493), .B(new_n494), .Z(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n269), .A2(new_n236), .ZN(new_n497));
  INV_X1    g311(.A(new_n325), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n252), .B1(new_n256), .B2(new_n250), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n266), .A2(new_n243), .A3(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n497), .A2(KEYINPUT28), .A3(new_n498), .A4(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n235), .B1(new_n266), .B2(new_n268), .ZN(new_n503));
  AOI211_X1 g317(.A(new_n499), .B(new_n219), .C1(new_n261), .C2(new_n265), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n325), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n499), .B1(new_n261), .B2(new_n265), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n269), .A2(new_n236), .B1(new_n507), .B2(new_n243), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT28), .B1(new_n508), .B2(new_n498), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n496), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT30), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n503), .B2(new_n504), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n501), .B(KEYINPUT30), .C1(new_n273), .C2(new_n235), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n513), .A3(new_n325), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT31), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n508), .A2(new_n498), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n514), .A2(new_n515), .A3(new_n495), .A4(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n510), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n514), .A2(new_n495), .A3(new_n516), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT31), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT68), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n519), .A2(KEYINPUT68), .A3(KEYINPUT31), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n518), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(G472), .A2(G902), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n491), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n509), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n528), .A2(new_n495), .A3(new_n505), .A4(new_n502), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT29), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n495), .B1(new_n514), .B2(new_n516), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n190), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n497), .A2(new_n501), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n325), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(KEYINPUT69), .A3(new_n516), .ZN(new_n536));
  OR3_X1    g350(.A1(new_n508), .A2(KEYINPUT69), .A3(new_n498), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(KEYINPUT28), .A3(new_n537), .ZN(new_n538));
  AND4_X1   g352(.A1(KEYINPUT29), .A2(new_n538), .A3(new_n495), .A4(new_n528), .ZN(new_n539));
  OAI21_X1  g353(.A(G472), .B1(new_n533), .B2(new_n539), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n510), .A2(new_n517), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n519), .A2(KEYINPUT68), .A3(KEYINPUT31), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT68), .B1(new_n519), .B2(KEYINPUT31), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(KEYINPUT32), .A3(new_n525), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n527), .A2(new_n540), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n457), .B1(G234), .B2(new_n190), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n410), .A2(new_n375), .ZN(new_n549));
  XOR2_X1   g363(.A(G119), .B(G128), .Z(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT24), .B(G110), .ZN(new_n551));
  OR2_X1    g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(KEYINPUT23), .B1(new_n217), .B2(G119), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT70), .B1(new_n217), .B2(G119), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n313), .A2(G128), .ZN(new_n555));
  OR2_X1    g369(.A1(KEYINPUT70), .A2(KEYINPUT23), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n553), .A2(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(G110), .ZN(new_n558));
  OR2_X1    g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n549), .A2(new_n552), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n557), .A2(new_n558), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n550), .A2(new_n551), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n561), .A2(new_n562), .B1(new_n212), .B2(new_n372), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n563), .A2(KEYINPUT72), .A3(new_n375), .ZN(new_n564));
  AOI21_X1  g378(.A(KEYINPUT72), .B1(new_n563), .B2(new_n375), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n560), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT22), .B(G137), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n300), .A2(G221), .A3(G234), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n569), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n560), .B(new_n571), .C1(new_n564), .C2(new_n565), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n570), .A2(new_n190), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT73), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(KEYINPUT25), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n575), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n570), .A2(new_n190), .A3(new_n572), .A4(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n548), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n547), .A2(G902), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n570), .A2(new_n572), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n546), .A2(KEYINPUT74), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(KEYINPUT74), .B1(new_n546), .B2(new_n584), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n297), .B(new_n490), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(G101), .ZN(G3));
  NAND2_X1  g402(.A1(KEYINPUT91), .A2(G472), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n590), .B1(new_n524), .B2(G902), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n544), .A2(new_n190), .A3(new_n589), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n591), .A2(new_n297), .A3(new_n584), .A4(new_n592), .ZN(new_n593));
  XOR2_X1   g407(.A(new_n593), .B(KEYINPUT92), .Z(new_n594));
  NAND2_X1  g408(.A1(new_n350), .A2(new_n353), .ZN(new_n595));
  INV_X1    g409(.A(new_n339), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n355), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n357), .A2(new_n339), .A3(new_n359), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n363), .B(new_n486), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n417), .A2(new_n419), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n423), .A2(new_n425), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n468), .A2(G902), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT93), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n473), .A2(new_n604), .A3(KEYINPUT33), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT33), .B1(new_n473), .B2(new_n604), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n467), .A2(new_n468), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n602), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n599), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n594), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT34), .B(G104), .Z(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G6));
  NAND3_X1  g428(.A1(new_n417), .A2(KEYINPUT94), .A3(new_n419), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT94), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n616), .B(KEYINPUT20), .C1(new_n414), .C2(new_n416), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n615), .A2(new_n601), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n480), .A2(new_n476), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n618), .A2(KEYINPUT95), .A3(new_n619), .A4(new_n486), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT95), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n619), .A2(new_n615), .A3(new_n601), .A4(new_n617), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n621), .B1(new_n622), .B2(new_n485), .ZN(new_n623));
  INV_X1    g437(.A(new_n363), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n354), .A2(new_n355), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n359), .B1(new_n357), .B2(new_n339), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n620), .A2(new_n623), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n594), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G107), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT96), .B(KEYINPUT35), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  OAI21_X1  g446(.A(new_n566), .B1(KEYINPUT36), .B2(new_n569), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n569), .A2(KEYINPUT36), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n560), .B(new_n634), .C1(new_n564), .C2(new_n565), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n633), .A2(new_n581), .A3(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT97), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n633), .A2(KEYINPUT97), .A3(new_n581), .A4(new_n635), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n579), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n591), .A2(new_n297), .A3(new_n592), .A4(new_n642), .ZN(new_n643));
  OR2_X1    g457(.A1(new_n643), .A2(new_n489), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT37), .B(G110), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G12));
  INV_X1    g460(.A(new_n297), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(new_n641), .ZN(new_n648));
  INV_X1    g462(.A(G900), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n483), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n482), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n622), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n627), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT98), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n627), .A2(new_n654), .A3(KEYINPUT98), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n648), .A2(new_n657), .A3(new_n546), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G128), .ZN(G30));
  XOR2_X1   g474(.A(new_n652), .B(KEYINPUT39), .Z(new_n661));
  NOR2_X1   g475(.A1(new_n647), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT40), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n514), .A2(new_n516), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n495), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n536), .A2(new_n537), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n190), .B(new_n665), .C1(new_n666), .C2(new_n495), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(G472), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n527), .A2(new_n545), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n602), .A2(new_n619), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n624), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n669), .A2(new_n641), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n673), .B(KEYINPUT100), .Z(new_n674));
  NAND3_X1  g488(.A1(new_n362), .A2(new_n366), .A3(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n674), .B1(new_n362), .B2(new_n366), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n663), .A2(new_n672), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G143), .ZN(G45));
  NOR2_X1   g494(.A1(new_n610), .A2(new_n653), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n648), .A2(new_n546), .A3(new_n627), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G146), .ZN(G48));
  OAI21_X1  g497(.A(new_n190), .B1(new_n293), .B2(new_n295), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(G469), .ZN(new_n685));
  INV_X1    g499(.A(new_n191), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n685), .A2(new_n686), .A3(new_n296), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(KEYINPUT101), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT101), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n685), .A2(new_n689), .A3(new_n686), .A4(new_n296), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n688), .A2(new_n611), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n546), .A2(new_n584), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT41), .B(G113), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G15));
  NAND3_X1  g509(.A1(new_n628), .A2(new_n688), .A3(new_n690), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(new_n692), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT102), .B(G116), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G18));
  AND3_X1   g513(.A1(new_n527), .A2(new_n540), .A3(new_n545), .ZN(new_n700));
  INV_X1    g514(.A(new_n296), .ZN(new_n701));
  INV_X1    g515(.A(new_n274), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n273), .B1(new_n245), .B2(KEYINPUT78), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n702), .B1(new_n703), .B2(new_n271), .ZN(new_n704));
  OAI22_X1  g518(.A1(new_n704), .A2(new_n279), .B1(new_n294), .B2(new_n280), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n292), .B1(new_n705), .B2(new_n190), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n701), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n487), .A2(new_n641), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n707), .A2(new_n686), .A3(new_n708), .A4(new_n627), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n700), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G119), .ZN(G21));
  OAI21_X1  g525(.A(G472), .B1(new_n524), .B2(G902), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT103), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI211_X1 g528(.A(KEYINPUT103), .B(G472), .C1(new_n524), .C2(G902), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n495), .B1(new_n538), .B2(new_n528), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n520), .A2(new_n517), .ZN(new_n717));
  OR2_X1    g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n525), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n714), .A2(new_n584), .A3(new_n715), .A4(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n599), .A2(new_n670), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n688), .A2(new_n690), .A3(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(KEYINPUT104), .B(G122), .Z(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G24));
  INV_X1    g539(.A(new_n681), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n363), .B1(new_n597), .B2(new_n598), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n687), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  AOI22_X1  g542(.A1(new_n712), .A2(new_n713), .B1(new_n525), .B2(new_n718), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n728), .A2(new_n729), .A3(new_n642), .A4(new_n715), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G125), .ZN(G27));
  NAND2_X1  g545(.A1(new_n362), .A2(new_n366), .ZN(new_n732));
  NAND2_X1  g546(.A1(G469), .A2(G902), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(KEYINPUT105), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n735), .B1(new_n290), .B2(G469), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n191), .B1(new_n736), .B2(new_n296), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n732), .A2(new_n363), .A3(new_n681), .A4(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT106), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n545), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n544), .A2(KEYINPUT106), .A3(KEYINPUT32), .A4(new_n525), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n741), .A2(new_n527), .A3(new_n540), .A4(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n739), .A2(KEYINPUT42), .A3(new_n584), .A4(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT42), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n624), .B1(new_n362), .B2(new_n366), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n746), .A2(new_n546), .A3(new_n584), .A4(new_n737), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n745), .B1(new_n747), .B2(new_n726), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G131), .ZN(G33));
  INV_X1    g564(.A(new_n747), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n654), .B(KEYINPUT107), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G134), .ZN(G36));
  AND2_X1   g568(.A1(new_n591), .A2(new_n592), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT111), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT43), .B1(new_n426), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n426), .A2(new_n609), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n426), .B(new_n609), .C1(new_n757), .C2(KEYINPUT43), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n641), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n756), .A2(new_n762), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n763), .A2(KEYINPUT44), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n756), .A2(KEYINPUT44), .A3(new_n762), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n746), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT46), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n735), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(G469), .B1(new_n290), .B2(KEYINPUT45), .ZN(new_n771));
  AOI22_X1  g585(.A1(new_n771), .A2(KEYINPUT108), .B1(KEYINPUT45), .B2(new_n290), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT108), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n773), .B(G469), .C1(new_n290), .C2(KEYINPUT45), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n770), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n767), .B1(new_n775), .B2(new_n701), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n771), .A2(KEYINPUT108), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n290), .A2(KEYINPUT45), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n774), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n769), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(KEYINPUT109), .A3(new_n296), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n779), .A2(new_n734), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n768), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n776), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n686), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT110), .ZN(new_n786));
  OR3_X1    g600(.A1(new_n785), .A2(new_n786), .A3(new_n661), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n786), .B1(new_n785), .B2(new_n661), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n766), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(new_n247), .ZN(G39));
  XNOR2_X1  g604(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n785), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n784), .A2(new_n686), .A3(new_n791), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n732), .A2(new_n363), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n795), .A2(new_n546), .A3(new_n584), .A4(new_n726), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n793), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G140), .ZN(G42));
  NAND2_X1  g612(.A1(new_n481), .A2(new_n300), .ZN(new_n799));
  AND4_X1   g613(.A1(new_n470), .A2(new_n618), .A3(new_n475), .A4(new_n652), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n732), .A2(KEYINPUT114), .A3(new_n363), .A4(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n801), .A2(new_n546), .A3(new_n648), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT114), .B1(new_n746), .B2(new_n800), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n752), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n714), .A2(new_n642), .A3(new_n715), .A4(new_n719), .ZN(new_n806));
  OAI22_X1  g620(.A1(new_n747), .A2(new_n805), .B1(new_n806), .B2(new_n738), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n749), .A2(new_n804), .A3(new_n808), .ZN(new_n809));
  OAI22_X1  g623(.A1(new_n700), .A2(new_n709), .B1(new_n643), .B2(new_n489), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n723), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n692), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n688), .A2(new_n690), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n812), .B(new_n813), .C1(new_n611), .C2(new_n628), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n470), .A2(new_n475), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n600), .A2(new_n601), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT113), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n816), .A2(new_n817), .B1(new_n602), .B2(new_n609), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n426), .A2(KEYINPUT113), .A3(new_n815), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n485), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n820), .A2(new_n363), .A3(new_n362), .A4(new_n366), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n593), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n811), .A2(new_n587), .A3(new_n814), .A4(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n809), .A2(new_n824), .ZN(new_n825));
  AOI211_X1 g639(.A(new_n624), .B(new_n670), .C1(new_n625), .C2(new_n626), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n642), .A2(new_n653), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n669), .A2(new_n826), .A3(new_n737), .A4(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n730), .A2(new_n659), .A3(new_n682), .A4(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n730), .A2(new_n659), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT52), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n825), .A2(KEYINPUT53), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n692), .B1(new_n696), .B2(new_n691), .ZN(new_n836));
  NOR4_X1   g650(.A1(new_n836), .A2(new_n723), .A3(new_n810), .A4(new_n822), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n802), .A2(new_n803), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n838), .A2(new_n807), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n837), .A2(new_n587), .A3(new_n749), .A4(new_n839), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n829), .B(KEYINPUT52), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n835), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n834), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n825), .A2(KEYINPUT53), .A3(new_n831), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n825), .A2(KEYINPUT116), .A3(KEYINPUT53), .A4(new_n831), .ZN(new_n848));
  INV_X1    g662(.A(new_n824), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT115), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n849), .A2(new_n850), .A3(new_n749), .A4(new_n839), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT115), .B1(new_n809), .B2(new_n824), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n851), .A2(new_n831), .A3(new_n833), .A4(new_n852), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n847), .A2(new_n848), .B1(new_n853), .B2(new_n835), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n844), .B1(new_n854), .B2(new_n843), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n743), .A2(new_n584), .ZN(new_n857));
  INV_X1    g671(.A(new_n687), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n651), .B1(new_n760), .B2(new_n761), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n746), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(KEYINPUT119), .A2(KEYINPUT48), .ZN(new_n862));
  AND2_X1   g676(.A1(KEYINPUT119), .A2(KEYINPUT48), .ZN(new_n863));
  OR3_X1    g677(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n584), .A2(new_n482), .ZN(new_n865));
  NOR4_X1   g679(.A1(new_n795), .A2(new_n669), .A3(new_n687), .A4(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n610), .ZN(new_n867));
  AOI211_X1 g681(.A(new_n481), .B(G953), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(G472), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(new_n544), .B2(new_n190), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n719), .B1(new_n870), .B2(KEYINPUT103), .ZN(new_n871));
  AOI211_X1 g685(.A(new_n713), .B(new_n869), .C1(new_n544), .C2(new_n190), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n873), .A2(new_n584), .A3(new_n859), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(new_n627), .A3(new_n858), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n861), .A2(new_n863), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n864), .A2(new_n868), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  AOI22_X1  g692(.A1(new_n793), .A2(new_n794), .B1(new_n191), .B2(new_n707), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n873), .A2(new_n584), .A3(new_n859), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n880), .A2(new_n795), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT117), .ZN(new_n883));
  OAI22_X1  g697(.A1(new_n879), .A2(new_n882), .B1(new_n883), .B2(KEYINPUT51), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT51), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n858), .A2(new_n624), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n678), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n874), .A2(new_n887), .A3(KEYINPUT50), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT50), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n624), .B(new_n858), .C1(new_n676), .C2(new_n677), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n889), .B1(new_n880), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n860), .A2(new_n806), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n602), .A2(new_n609), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n893), .B1(new_n866), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n885), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n878), .B1(new_n884), .B2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT118), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n888), .A2(new_n891), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n898), .B1(new_n888), .B2(new_n891), .ZN(new_n900));
  INV_X1    g714(.A(new_n895), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n794), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n791), .B1(new_n784), .B2(new_n686), .ZN(new_n904));
  INV_X1    g718(.A(new_n707), .ZN(new_n905));
  OAI22_X1  g719(.A1(new_n903), .A2(new_n904), .B1(new_n686), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(KEYINPUT117), .A3(new_n881), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT51), .B1(new_n902), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n856), .B1(new_n897), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n900), .A2(new_n901), .ZN(new_n910));
  INV_X1    g724(.A(new_n899), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n879), .A2(new_n883), .A3(new_n882), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n885), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI22_X1  g728(.A1(new_n906), .A2(new_n881), .B1(KEYINPUT117), .B2(new_n885), .ZN(new_n915));
  INV_X1    g729(.A(new_n896), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n877), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n914), .A2(new_n917), .A3(KEYINPUT120), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n909), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n799), .B1(new_n855), .B2(new_n919), .ZN(new_n920));
  NOR4_X1   g734(.A1(new_n583), .A2(new_n759), .A3(new_n191), .A4(new_n624), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT49), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n921), .B1(new_n922), .B2(new_n707), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n905), .A2(KEYINPUT49), .ZN(new_n924));
  OR4_X1    g738(.A1(new_n678), .A2(new_n669), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n920), .A2(new_n925), .ZN(G75));
  NAND2_X1  g740(.A1(new_n481), .A2(G953), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT123), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n834), .A2(new_n842), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n929), .A2(KEYINPUT122), .A3(G210), .A4(G902), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n350), .A2(new_n353), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n931), .A2(new_n357), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT55), .Z(new_n933));
  NOR2_X1   g747(.A1(new_n933), .A2(KEYINPUT56), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n190), .B1(new_n834), .B2(new_n842), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT122), .B1(new_n936), .B2(G210), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n928), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT121), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT56), .B1(new_n936), .B2(G210), .ZN(new_n940));
  INV_X1    g754(.A(new_n933), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n936), .A2(G210), .ZN(new_n943));
  OAI211_X1 g757(.A(KEYINPUT121), .B(new_n933), .C1(new_n943), .C2(KEYINPUT56), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n938), .B1(new_n942), .B2(new_n944), .ZN(G51));
  INV_X1    g759(.A(new_n928), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n734), .B(KEYINPUT57), .Z(new_n947));
  INV_X1    g761(.A(new_n844), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n843), .B1(new_n834), .B2(new_n842), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n705), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n936), .A2(new_n774), .A3(new_n772), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n946), .B1(new_n951), .B2(new_n952), .ZN(G54));
  NAND3_X1  g767(.A1(new_n936), .A2(KEYINPUT58), .A3(G475), .ZN(new_n954));
  INV_X1    g768(.A(new_n414), .ZN(new_n955));
  OR2_X1    g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n954), .A2(new_n955), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n946), .B1(new_n956), .B2(new_n957), .ZN(G60));
  OR2_X1    g772(.A1(new_n605), .A2(new_n606), .ZN(new_n959));
  NAND2_X1  g773(.A1(G478), .A2(G902), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT59), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n959), .B(new_n961), .C1(new_n948), .C2(new_n949), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n928), .ZN(new_n963));
  INV_X1    g777(.A(new_n959), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n847), .A2(new_n848), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n853), .A2(new_n835), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n843), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n961), .B1(new_n967), .B2(new_n948), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n963), .B1(new_n964), .B2(new_n968), .ZN(G63));
  NAND2_X1  g783(.A1(G217), .A2(G902), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT60), .Z(new_n971));
  NAND2_X1  g785(.A1(new_n929), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n633), .A2(new_n635), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n570), .A2(new_n572), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT124), .Z(new_n976));
  AOI21_X1  g790(.A(new_n946), .B1(new_n972), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT61), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n974), .A2(KEYINPUT61), .A3(new_n977), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(G66));
  INV_X1    g796(.A(G224), .ZN(new_n983));
  OAI21_X1  g797(.A(G953), .B1(new_n484), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n849), .B2(G953), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n346), .B(new_n349), .C1(G898), .C2(new_n300), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT125), .Z(new_n987));
  XNOR2_X1  g801(.A(new_n985), .B(new_n987), .ZN(G69));
  NAND2_X1  g802(.A1(new_n787), .A2(new_n788), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n989), .A2(new_n584), .A3(new_n743), .A4(new_n826), .ZN(new_n990));
  INV_X1    g804(.A(new_n789), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n730), .A2(new_n659), .A3(new_n682), .ZN(new_n992));
  AND4_X1   g806(.A1(new_n749), .A2(new_n797), .A3(new_n753), .A4(new_n992), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n990), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n512), .A2(new_n513), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(new_n392), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(G953), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n679), .A2(new_n992), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n999), .A2(KEYINPUT62), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(KEYINPUT126), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n818), .A2(new_n819), .ZN(new_n1002));
  AND3_X1   g816(.A1(new_n662), .A2(new_n746), .A3(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1003), .B1(new_n585), .B2(new_n586), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n797), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1005), .B1(KEYINPUT62), .B2(new_n999), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1001), .A2(new_n991), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(new_n996), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n997), .A2(G227), .ZN(new_n1009));
  AOI211_X1 g823(.A(new_n649), .B(new_n300), .C1(new_n996), .C2(new_n276), .ZN(new_n1010));
  AOI22_X1  g824(.A1(new_n998), .A2(new_n1008), .B1(new_n1009), .B2(new_n1010), .ZN(G72));
  NAND3_X1  g825(.A1(new_n514), .A2(new_n496), .A3(new_n516), .ZN(new_n1012));
  NAND2_X1  g826(.A1(G472), .A2(G902), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1013), .B(KEYINPUT63), .Z(new_n1014));
  NAND3_X1  g828(.A1(new_n665), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n854), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n1001), .A2(new_n1006), .A3(new_n991), .A4(new_n849), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1014), .B(KEYINPUT127), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n665), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n990), .A2(new_n993), .A3(new_n991), .A4(new_n849), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1012), .B1(new_n1020), .B2(new_n1018), .ZN(new_n1021));
  NOR4_X1   g835(.A1(new_n1016), .A2(new_n1019), .A3(new_n946), .A4(new_n1021), .ZN(G57));
endmodule


