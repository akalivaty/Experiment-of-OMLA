//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 1 0 1 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 1 0 1 1 0 0 0 1 1 0 0 0 1 0 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n852, new_n853, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n995,
    new_n996, new_n997;
  XNOR2_X1  g000(.A(KEYINPUT83), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g002(.A1(G228gat), .A2(G233gat), .ZN(new_n204));
  XOR2_X1   g003(.A(KEYINPUT74), .B(G162gat), .Z(new_n205));
  INV_X1    g004(.A(G155gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT2), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G141gat), .ZN(new_n208));
  INV_X1    g007(.A(G148gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  OR2_X1    g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n207), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n212), .A2(KEYINPUT73), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT73), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n210), .A2(new_n218), .A3(new_n211), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n217), .A2(new_n219), .B1(KEYINPUT72), .B2(KEYINPUT2), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n213), .B(KEYINPUT72), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(new_n214), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n216), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n224), .B(KEYINPUT69), .ZN(new_n225));
  XNOR2_X1  g024(.A(G197gat), .B(G204gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT68), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n226), .A2(new_n227), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n225), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G211gat), .B(G218gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n226), .B(new_n227), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(new_n231), .A3(new_n225), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT29), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n223), .B1(new_n236), .B2(KEYINPUT3), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT81), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n204), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n216), .B(new_n240), .C1(new_n220), .C2(new_n222), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT29), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n233), .A2(new_n235), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT82), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  OAI211_X1 g045(.A(KEYINPUT81), .B(new_n223), .C1(new_n236), .C2(KEYINPUT3), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n243), .A2(new_n244), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT82), .ZN(new_n249));
  AND4_X1   g048(.A1(new_n239), .A2(new_n246), .A3(new_n247), .A4(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n223), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n233), .A2(new_n235), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(new_n242), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n251), .B1(new_n253), .B2(new_n240), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT80), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n255), .B1(new_n243), .B2(new_n244), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n243), .A2(new_n244), .A3(new_n255), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n257), .A2(new_n258), .B1(G228gat), .B2(G233gat), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n203), .B1(new_n250), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT84), .ZN(new_n261));
  INV_X1    g060(.A(new_n256), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n262), .A2(new_n258), .A3(new_n237), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(new_n204), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n239), .A2(new_n246), .A3(new_n247), .A4(new_n249), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(new_n202), .A3(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n260), .A2(new_n261), .A3(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n250), .A2(new_n259), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n268), .A2(KEYINPUT84), .A3(new_n202), .ZN(new_n269));
  XNOR2_X1  g068(.A(G78gat), .B(G106gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT78), .ZN(new_n271));
  XOR2_X1   g070(.A(KEYINPUT31), .B(G50gat), .Z(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  XOR2_X1   g072(.A(new_n273), .B(KEYINPUT79), .Z(new_n274));
  NAND3_X1  g073(.A1(new_n267), .A2(new_n269), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G22gat), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n266), .B(new_n273), .C1(new_n268), .C2(new_n276), .ZN(new_n277));
  AND2_X1   g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n279));
  XNOR2_X1  g078(.A(G127gat), .B(G134gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT65), .ZN(new_n281));
  INV_X1    g080(.A(G134gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(G127gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(G113gat), .B(G120gat), .ZN(new_n284));
  OAI221_X1 g083(.A(new_n281), .B1(KEYINPUT65), .B2(new_n283), .C1(KEYINPUT1), .C2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT66), .ZN(new_n286));
  INV_X1    g085(.A(G120gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n286), .B1(new_n287), .B2(G113gat), .ZN(new_n288));
  INV_X1    g087(.A(G113gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n289), .A2(KEYINPUT66), .A3(G120gat), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n288), .B(new_n290), .C1(new_n289), .C2(G120gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT1), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n291), .A2(new_n292), .A3(new_n280), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n285), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n223), .B(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G225gat), .A2(G233gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n279), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n223), .A2(new_n294), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n297), .B1(new_n299), .B2(KEYINPUT4), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n223), .A2(KEYINPUT3), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(new_n241), .A3(new_n294), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT75), .B(KEYINPUT4), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n303), .B1(new_n223), .B2(new_n294), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n300), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n298), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n294), .ZN(new_n307));
  INV_X1    g106(.A(new_n303), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n251), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT4), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n310), .B1(new_n223), .B2(new_n294), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n297), .A2(KEYINPUT5), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n302), .A2(new_n309), .A3(new_n311), .A4(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n306), .A2(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(G1gat), .B(G29gat), .Z(new_n315));
  XNOR2_X1  g114(.A(new_n315), .B(KEYINPUT0), .ZN(new_n316));
  XNOR2_X1  g115(.A(G57gat), .B(G85gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n316), .B(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n313), .A2(new_n318), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT6), .B1(new_n321), .B2(new_n306), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT76), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AOI211_X1 g123(.A(KEYINPUT76), .B(KEYINPUT6), .C1(new_n321), .C2(new_n306), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT77), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n321), .A2(new_n306), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT76), .B1(new_n327), .B2(KEYINPUT6), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT77), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n322), .A2(new_n323), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n328), .A2(new_n329), .A3(new_n330), .A4(new_n320), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n314), .A2(KEYINPUT6), .A3(new_n319), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n326), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(G8gat), .B(G36gat), .Z(new_n334));
  XNOR2_X1  g133(.A(new_n334), .B(KEYINPUT71), .ZN(new_n335));
  XNOR2_X1  g134(.A(G64gat), .B(G92gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G226gat), .A2(G233gat), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n339), .B(KEYINPUT70), .Z(new_n340));
  OAI21_X1  g139(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT23), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(G183gat), .ZN(new_n344));
  INV_X1    g143(.A(G190gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G183gat), .A2(G190gat), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n346), .A2(KEYINPUT24), .A3(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(KEYINPUT24), .ZN(new_n349));
  INV_X1    g148(.A(G169gat), .ZN(new_n350));
  INV_X1    g149(.A(G176gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n343), .A2(KEYINPUT25), .A3(new_n348), .A4(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n343), .A2(new_n348), .A3(new_n353), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT25), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT27), .B(G183gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n345), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT28), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(G169gat), .A2(G176gat), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n352), .A2(KEYINPUT26), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(KEYINPUT26), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n347), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n354), .A2(new_n357), .B1(new_n361), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n340), .B1(new_n367), .B2(KEYINPUT29), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n357), .A2(new_n354), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n361), .A2(new_n366), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n340), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n368), .A2(new_n373), .A3(new_n252), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n252), .B1(new_n368), .B2(new_n373), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n338), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n376), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n378), .A2(new_n337), .A3(new_n374), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n377), .A2(new_n379), .A3(KEYINPUT30), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT30), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n378), .A2(new_n381), .A3(new_n337), .A4(new_n374), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n278), .B1(new_n333), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT36), .ZN(new_n386));
  XNOR2_X1  g185(.A(G15gat), .B(G43gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(G71gat), .B(G99gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n371), .A2(new_n307), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n367), .A2(new_n294), .ZN(new_n391));
  INV_X1    g190(.A(G227gat), .ZN(new_n392));
  INV_X1    g191(.A(G233gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n390), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n389), .B1(new_n395), .B2(KEYINPUT32), .ZN(new_n396));
  INV_X1    g195(.A(new_n395), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n396), .B1(KEYINPUT33), .B2(new_n397), .ZN(new_n398));
  OR2_X1    g197(.A1(new_n389), .A2(KEYINPUT67), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n389), .A2(KEYINPUT67), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(KEYINPUT33), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n395), .A2(KEYINPUT32), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n390), .A2(new_n391), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n404), .B1(new_n392), .B2(new_n393), .ZN(new_n405));
  OR2_X1    g204(.A1(new_n405), .A2(KEYINPUT34), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(KEYINPUT34), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AND2_X1   g207(.A1(new_n403), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n398), .A2(new_n406), .A3(new_n402), .A4(new_n407), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n386), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n403), .A2(new_n408), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n413), .A2(KEYINPUT36), .A3(new_n410), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  OR3_X1    g214(.A1(new_n375), .A2(KEYINPUT37), .A3(new_n376), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT37), .B1(new_n375), .B2(new_n376), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n416), .A2(new_n338), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT38), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n379), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n320), .A2(new_n322), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n416), .A2(new_n419), .A3(new_n338), .A4(new_n417), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n421), .A2(new_n422), .A3(new_n332), .A4(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n302), .A2(new_n311), .A3(new_n309), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n297), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT85), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT85), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n425), .A2(new_n428), .A3(new_n297), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT39), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n319), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OR2_X1    g231(.A1(new_n295), .A2(new_n297), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n427), .A2(KEYINPUT39), .A3(new_n429), .A4(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n432), .A2(KEYINPUT40), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n384), .A2(new_n435), .A3(new_n320), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT40), .B1(new_n432), .B2(new_n434), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n424), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n385), .B(new_n415), .C1(new_n278), .C2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n383), .A2(new_n413), .A3(new_n410), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n440), .B1(new_n275), .B2(new_n277), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n422), .A2(new_n332), .ZN(new_n442));
  XOR2_X1   g241(.A(KEYINPUT86), .B(KEYINPUT35), .Z(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT35), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n326), .A2(new_n331), .A3(new_n332), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n446), .B1(new_n441), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n445), .B1(new_n448), .B2(KEYINPUT87), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT87), .ZN(new_n450));
  AOI211_X1 g249(.A(new_n450), .B(new_n446), .C1(new_n441), .C2(new_n447), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n439), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n453), .B(new_n206), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(G15gat), .B(G22gat), .ZN(new_n456));
  INV_X1    g255(.A(G1gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT16), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(G15gat), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n460), .A2(G22gat), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n276), .A2(G15gat), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n457), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(KEYINPUT93), .ZN(new_n465));
  INV_X1    g264(.A(G8gat), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n459), .B(new_n463), .C1(KEYINPUT93), .C2(G8gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT94), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT94), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  XOR2_X1   g273(.A(G57gat), .B(G64gat), .Z(new_n475));
  OR2_X1    g274(.A1(G71gat), .A2(G78gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(G71gat), .A2(G78gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT9), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n475), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(G57gat), .B(G64gat), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n477), .B(new_n476), .C1(new_n482), .C2(new_n479), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT21), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n474), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT96), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT96), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n474), .A2(new_n488), .A3(new_n485), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n455), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n481), .A2(new_n483), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT21), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(G231gat), .A2(G233gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(G127gat), .ZN(new_n497));
  OR2_X1    g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n497), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G183gat), .B(G211gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n501), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n498), .A2(new_n503), .A3(new_n499), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n487), .A2(new_n489), .A3(new_n455), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n491), .A2(new_n502), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n502), .A2(new_n504), .ZN(new_n507));
  INV_X1    g306(.A(new_n505), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n507), .B1(new_n508), .B2(new_n490), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(G232gat), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n511), .A2(new_n393), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT41), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G190gat), .B(G218gat), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT98), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n515), .B(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  AND2_X1   g319(.A1(G43gat), .A2(G50gat), .ZN(new_n521));
  NOR2_X1   g320(.A1(G43gat), .A2(G50gat), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT15), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR3_X1   g322(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT89), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n527), .B1(new_n525), .B2(new_n526), .ZN(new_n528));
  NAND2_X1  g327(.A1(G29gat), .A2(G36gat), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n523), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G43gat), .B(G50gat), .ZN(new_n531));
  AOI22_X1  g330(.A1(new_n531), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT90), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n521), .A2(new_n522), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT15), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR4_X1   g335(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT90), .A4(KEYINPUT15), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n532), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT91), .ZN(new_n539));
  INV_X1    g338(.A(new_n526), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n539), .B1(new_n540), .B2(new_n524), .ZN(new_n541));
  OR2_X1    g340(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n542));
  OAI211_X1 g341(.A(KEYINPUT91), .B(new_n526), .C1(new_n542), .C2(G36gat), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT92), .B1(new_n538), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n523), .A2(new_n529), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT90), .B1(new_n531), .B2(KEYINPUT15), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n534), .A2(new_n533), .A3(new_n535), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT92), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n541), .A2(new_n543), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n530), .B1(new_n545), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G85gat), .A2(G92gat), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT7), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G99gat), .A2(G106gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT8), .ZN(new_n560));
  INV_X1    g359(.A(G85gat), .ZN(new_n561));
  INV_X1    g360(.A(G92gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n559), .ZN(new_n565));
  NOR2_X1   g364(.A1(G99gat), .A2(G106gat), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT97), .ZN(new_n567));
  NOR3_X1   g366(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(G99gat), .ZN(new_n569));
  INV_X1    g368(.A(G106gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(KEYINPUT97), .B1(new_n571), .B2(new_n559), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n558), .B(new_n564), .C1(new_n568), .C2(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n560), .A2(new_n556), .A3(new_n563), .A4(new_n557), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n567), .B1(new_n565), .B2(new_n566), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n571), .A2(KEYINPUT97), .A3(new_n559), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  OAI22_X1  g377(.A1(new_n553), .A2(new_n578), .B1(new_n514), .B2(new_n513), .ZN(new_n579));
  INV_X1    g378(.A(new_n578), .ZN(new_n580));
  INV_X1    g379(.A(new_n530), .ZN(new_n581));
  NOR3_X1   g380(.A1(new_n538), .A2(new_n544), .A3(KEYINPUT92), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n550), .B1(new_n549), .B2(new_n551), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT17), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n580), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n553), .A2(KEYINPUT17), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n579), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n516), .A2(new_n517), .ZN(new_n589));
  XNOR2_X1  g388(.A(G134gat), .B(G162gat), .ZN(new_n590));
  NOR3_X1   g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n590), .ZN(new_n592));
  AOI22_X1  g391(.A1(new_n584), .A2(new_n580), .B1(KEYINPUT41), .B2(new_n512), .ZN(new_n593));
  AOI211_X1 g392(.A(new_n585), .B(new_n530), .C1(new_n545), .C2(new_n552), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n578), .B1(new_n553), .B2(KEYINPUT17), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n589), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n592), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n520), .B1(new_n591), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n590), .B1(new_n588), .B2(new_n589), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n596), .A2(new_n597), .A3(new_n592), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n600), .A2(new_n519), .A3(new_n601), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(KEYINPUT99), .B1(new_n510), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n506), .A2(new_n509), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n599), .A2(new_n602), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT99), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n580), .A2(KEYINPUT10), .A3(new_n484), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT100), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n568), .A2(new_n572), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n610), .B1(new_n611), .B2(new_n574), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n578), .A2(new_n612), .A3(new_n484), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n573), .B(new_n577), .C1(new_n492), .C2(new_n610), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT10), .ZN(new_n616));
  AOI21_X1  g415(.A(KEYINPUT101), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT101), .ZN(new_n618));
  AOI211_X1 g417(.A(new_n618), .B(KEYINPUT10), .C1(new_n613), .C2(new_n614), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n609), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G230gat), .A2(G233gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n621), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n613), .A2(new_n623), .A3(new_n614), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G120gat), .B(G148gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(G176gat), .B(G204gat), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n626), .B(new_n627), .Z(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n622), .A2(new_n624), .A3(new_n628), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n604), .A2(new_n608), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n584), .A2(new_n473), .ZN(new_n636));
  NAND2_X1  g435(.A1(G229gat), .A2(G233gat), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n469), .B1(new_n553), .B2(KEYINPUT17), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n636), .B(new_n637), .C1(new_n638), .C2(new_n594), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT18), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n637), .B(KEYINPUT13), .Z(new_n642));
  NOR2_X1   g441(.A1(new_n584), .A2(new_n473), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n545), .A2(new_n552), .ZN(new_n644));
  AOI22_X1  g443(.A1(new_n644), .A2(new_n581), .B1(new_n471), .B2(new_n472), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n642), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n584), .A2(new_n585), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n647), .A2(new_n469), .A3(new_n587), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n648), .A2(KEYINPUT18), .A3(new_n636), .A4(new_n637), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n641), .A2(new_n646), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT95), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n651), .B(new_n646), .C1(new_n639), .C2(new_n640), .ZN(new_n652));
  XNOR2_X1  g451(.A(G113gat), .B(G141gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G169gat), .B(G197gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n657), .B(KEYINPUT12), .Z(new_n658));
  NAND2_X1  g457(.A1(new_n652), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n650), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n641), .A2(new_n649), .A3(new_n646), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n661), .A2(new_n652), .A3(new_n658), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n452), .A2(new_n635), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT102), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n452), .A2(new_n635), .A3(new_n666), .A4(new_n663), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n333), .A2(KEYINPUT103), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n333), .A2(KEYINPUT103), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g473(.A(KEYINPUT16), .B(G8gat), .Z(new_n675));
  NAND3_X1  g474(.A1(new_n668), .A2(new_n384), .A3(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT42), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n676), .A2(KEYINPUT104), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT104), .ZN(new_n679));
  INV_X1    g478(.A(new_n676), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n679), .B1(new_n680), .B2(KEYINPUT42), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n466), .B1(new_n668), .B2(new_n384), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n676), .B1(new_n682), .B2(new_n677), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n678), .B1(new_n681), .B2(new_n683), .ZN(G1325gat));
  INV_X1    g483(.A(new_n668), .ZN(new_n685));
  OAI21_X1  g484(.A(G15gat), .B1(new_n685), .B2(new_n415), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n409), .A2(new_n411), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n668), .A2(new_n460), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(G1326gat));
  NAND2_X1  g488(.A1(new_n668), .A2(new_n278), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT43), .B(G22gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  OAI21_X1  g491(.A(new_n415), .B1(new_n438), .B2(new_n278), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n275), .A2(new_n277), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n694), .B1(new_n447), .B2(new_n383), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n440), .ZN(new_n697));
  AND4_X1   g496(.A1(new_n694), .A2(new_n697), .A3(new_n442), .A4(new_n444), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n694), .A2(new_n447), .A3(new_n697), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT35), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n698), .B1(new_n700), .B2(new_n450), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n448), .A2(KEYINPUT87), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n696), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n663), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n510), .A2(new_n633), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n606), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT105), .Z(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(G29gat), .A3(new_n671), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n713), .B1(new_n703), .B2(new_n606), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n452), .A2(KEYINPUT44), .A3(new_n603), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n716), .A2(new_n704), .A3(new_n706), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n672), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(G29gat), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n712), .A2(new_n719), .ZN(G1328gat));
  NOR3_X1   g519(.A1(new_n709), .A2(G36gat), .A3(new_n383), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT46), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n717), .A2(new_n384), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(G36gat), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(G1329gat));
  AND3_X1   g524(.A1(new_n452), .A2(KEYINPUT44), .A3(new_n603), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT44), .B1(new_n452), .B2(new_n603), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n415), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n706), .A2(new_n704), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n728), .A2(G43gat), .A3(new_n729), .A4(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(G43gat), .ZN(new_n732));
  INV_X1    g531(.A(new_n687), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n709), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g535(.A1(new_n728), .A2(new_n278), .A3(new_n730), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G50gat), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n694), .A2(G50gat), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT107), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n705), .A2(new_n708), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT48), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n738), .A2(KEYINPUT48), .A3(new_n741), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(G1331gat));
  NAND4_X1  g545(.A1(new_n604), .A2(new_n704), .A3(new_n608), .A4(new_n632), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n703), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n672), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n384), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n752));
  XOR2_X1   g551(.A(KEYINPUT49), .B(G64gat), .Z(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n751), .B2(new_n753), .ZN(G1333gat));
  NAND2_X1  g553(.A1(new_n748), .A2(new_n729), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n733), .A2(G71gat), .ZN(new_n756));
  AOI22_X1  g555(.A1(new_n755), .A2(G71gat), .B1(new_n748), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(G1334gat));
  NAND2_X1  g558(.A1(new_n748), .A2(new_n278), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g560(.A1(new_n663), .A2(new_n605), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n703), .A2(new_n606), .A3(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(KEYINPUT51), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n700), .A2(new_n450), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n766), .A2(new_n702), .A3(new_n445), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n606), .B1(new_n767), .B2(new_n439), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n768), .A2(KEYINPUT109), .A3(KEYINPUT51), .A4(new_n762), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n452), .A2(KEYINPUT51), .A3(new_n603), .A4(new_n762), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n765), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n769), .A2(new_n772), .A3(KEYINPUT110), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n672), .A2(new_n561), .A3(new_n632), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n763), .A2(new_n633), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n716), .A2(new_n671), .A3(new_n780), .ZN(new_n781));
  OAI22_X1  g580(.A1(new_n777), .A2(new_n778), .B1(new_n561), .B2(new_n781), .ZN(G1336gat));
  NAND3_X1  g581(.A1(new_n384), .A2(new_n562), .A3(new_n632), .ZN(new_n783));
  INV_X1    g582(.A(new_n765), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n784), .B2(new_n773), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n714), .A2(new_n384), .A3(new_n715), .A4(new_n779), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n786), .A2(G92gat), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT52), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n786), .A2(KEYINPUT111), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G92gat), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n786), .A2(KEYINPUT111), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n789), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n783), .B1(new_n775), .B2(new_n776), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n788), .B1(new_n793), .B2(new_n794), .ZN(G1337gat));
  NAND3_X1  g594(.A1(new_n687), .A2(new_n569), .A3(new_n632), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n716), .A2(new_n415), .A3(new_n780), .ZN(new_n797));
  OAI22_X1  g596(.A1(new_n777), .A2(new_n796), .B1(new_n569), .B2(new_n797), .ZN(G1338gat));
  NAND3_X1  g597(.A1(new_n278), .A2(new_n570), .A3(new_n632), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n799), .B1(new_n784), .B2(new_n773), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n714), .A2(new_n278), .A3(new_n715), .A4(new_n779), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(G106gat), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT53), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  OR2_X1    g602(.A1(new_n802), .A2(KEYINPUT53), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n799), .B1(new_n775), .B2(new_n776), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(G1339gat));
  NAND4_X1  g605(.A1(new_n604), .A2(new_n704), .A3(new_n608), .A4(new_n633), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n623), .B(new_n609), .C1(new_n617), .C2(new_n619), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n622), .A2(KEYINPUT54), .A3(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n620), .A2(new_n813), .A3(new_n621), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n629), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n810), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n622), .A2(KEYINPUT54), .A3(new_n811), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n817), .A2(KEYINPUT55), .A3(new_n629), .A4(new_n814), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n816), .A2(new_n631), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n637), .B1(new_n648), .B2(new_n636), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n643), .A2(new_n645), .A3(new_n642), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n657), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n658), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n641), .A2(new_n649), .A3(new_n646), .A4(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n599), .A2(new_n602), .A3(new_n822), .A4(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n809), .B1(new_n819), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n818), .A2(new_n631), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n814), .A2(new_n629), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT55), .B1(new_n828), .B2(new_n817), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n825), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n830), .A2(new_n831), .A3(KEYINPUT112), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n632), .A2(new_n822), .A3(new_n824), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n834), .B1(new_n830), .B2(new_n663), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n826), .B(new_n832), .C1(new_n835), .C2(new_n603), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n808), .B1(new_n836), .B2(new_n510), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n837), .A2(new_n278), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n671), .A2(new_n440), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(G113gat), .B1(new_n841), .B2(new_n663), .ZN(new_n842));
  INV_X1    g641(.A(new_n839), .ZN(new_n843));
  OR3_X1    g642(.A1(new_n837), .A2(KEYINPUT113), .A3(new_n278), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT113), .B1(new_n837), .B2(new_n278), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n704), .A2(new_n289), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n842), .B1(new_n846), .B2(new_n847), .ZN(G1340gat));
  AOI21_X1  g647(.A(G120gat), .B1(new_n841), .B2(new_n632), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n633), .A2(new_n287), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n849), .B1(new_n846), .B2(new_n850), .ZN(G1341gat));
  NOR2_X1   g650(.A1(new_n840), .A2(new_n510), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n852), .A2(KEYINPUT114), .ZN(new_n853));
  AOI21_X1  g652(.A(G127gat), .B1(new_n852), .B2(KEYINPUT114), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n510), .A2(new_n497), .ZN(new_n855));
  AOI22_X1  g654(.A1(new_n853), .A2(new_n854), .B1(new_n846), .B2(new_n855), .ZN(G1342gat));
  NAND2_X1  g655(.A1(new_n832), .A2(new_n826), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n818), .A2(new_n631), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n663), .A3(new_n816), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n603), .B1(new_n859), .B2(new_n833), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n510), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n807), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n694), .A2(new_n687), .ZN(new_n863));
  NOR4_X1   g662(.A1(new_n863), .A2(G134gat), .A3(new_n384), .A4(new_n606), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n862), .A2(new_n672), .A3(new_n864), .ZN(new_n865));
  XOR2_X1   g664(.A(new_n865), .B(KEYINPUT56), .Z(new_n866));
  AND2_X1   g665(.A1(new_n846), .A2(new_n603), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n866), .B1(new_n867), .B2(new_n282), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT115), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT115), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n866), .B(new_n870), .C1(new_n867), .C2(new_n282), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(G1343gat));
  AOI21_X1  g671(.A(new_n694), .B1(new_n861), .B2(new_n807), .ZN(new_n873));
  OAI21_X1  g672(.A(KEYINPUT116), .B1(new_n873), .B2(KEYINPUT57), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n875), .B(new_n876), .C1(new_n837), .C2(new_n694), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n828), .A2(new_n817), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n879));
  AOI21_X1  g678(.A(KEYINPUT55), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n828), .A2(KEYINPUT117), .A3(new_n817), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n827), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n834), .B1(new_n882), .B2(new_n663), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT118), .B1(new_n883), .B2(new_n603), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n878), .A2(new_n879), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n810), .A3(new_n881), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n663), .A3(new_n858), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(new_n833), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(new_n889), .A3(new_n606), .ZN(new_n890));
  INV_X1    g689(.A(new_n857), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n884), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n808), .B1(new_n892), .B2(new_n510), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n278), .A2(KEYINPUT57), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n874), .B(new_n877), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n671), .A2(new_n384), .A3(new_n729), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(G141gat), .B1(new_n897), .B2(new_n704), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n729), .A2(new_n694), .ZN(new_n899));
  XOR2_X1   g698(.A(new_n899), .B(KEYINPUT119), .Z(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n672), .A3(new_n862), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n901), .A2(new_n384), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n208), .A3(new_n663), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n898), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT58), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT58), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n898), .A2(new_n906), .A3(new_n903), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(new_n907), .ZN(G1344gat));
  NAND2_X1  g707(.A1(new_n896), .A2(new_n632), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n883), .A2(new_n603), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n819), .A2(new_n825), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n510), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n807), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n278), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n876), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n873), .A2(KEYINPUT57), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n909), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT59), .B1(new_n917), .B2(new_n209), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n895), .A2(new_n632), .A3(new_n896), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n209), .A2(KEYINPUT59), .ZN(new_n920));
  AND3_X1   g719(.A1(new_n919), .A2(KEYINPUT120), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(KEYINPUT120), .B1(new_n919), .B2(new_n920), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n918), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n902), .A2(new_n209), .A3(new_n632), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(G1345gat));
  OAI21_X1  g724(.A(G155gat), .B1(new_n897), .B2(new_n510), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n902), .A2(new_n206), .A3(new_n605), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1346gat));
  AND2_X1   g727(.A1(new_n895), .A2(new_n896), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n929), .A2(KEYINPUT121), .A3(new_n603), .ZN(new_n930));
  INV_X1    g729(.A(new_n205), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(KEYINPUT121), .B1(new_n929), .B2(new_n603), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n603), .A2(new_n205), .A3(new_n383), .ZN(new_n934));
  OAI22_X1  g733(.A1(new_n932), .A2(new_n933), .B1(new_n901), .B2(new_n934), .ZN(G1347gat));
  NAND3_X1  g734(.A1(new_n671), .A2(new_n384), .A3(new_n687), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n936), .B1(new_n844), .B2(new_n845), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n704), .A2(new_n350), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n837), .A2(new_n672), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n863), .A2(new_n383), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n939), .A2(new_n663), .A3(new_n940), .ZN(new_n941));
  AOI22_X1  g740(.A1(new_n937), .A2(new_n938), .B1(new_n350), .B2(new_n941), .ZN(G1348gat));
  NAND3_X1  g741(.A1(new_n937), .A2(G176gat), .A3(new_n632), .ZN(new_n943));
  OR2_X1    g742(.A1(new_n943), .A2(KEYINPUT122), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n939), .A2(new_n940), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n351), .B1(new_n945), .B2(new_n633), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n943), .A2(KEYINPUT122), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n944), .A2(new_n946), .A3(new_n947), .ZN(G1349gat));
  AND2_X1   g747(.A1(new_n937), .A2(new_n605), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n949), .A2(new_n344), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n605), .A2(new_n358), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n945), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(KEYINPUT60), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT60), .ZN(new_n954));
  OAI221_X1 g753(.A(new_n954), .B1(new_n945), .B2(new_n951), .C1(new_n949), .C2(new_n344), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n953), .A2(new_n955), .ZN(G1350gat));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n937), .A2(new_n603), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n958), .B2(G190gat), .ZN(new_n959));
  AOI211_X1 g758(.A(KEYINPUT61), .B(new_n345), .C1(new_n937), .C2(new_n603), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n603), .A2(new_n345), .ZN(new_n961));
  OAI22_X1  g760(.A1(new_n959), .A2(new_n960), .B1(new_n945), .B2(new_n961), .ZN(G1351gat));
  NAND3_X1  g761(.A1(new_n915), .A2(KEYINPUT125), .A3(new_n916), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n672), .A2(new_n383), .A3(new_n729), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT125), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT57), .B1(new_n913), .B2(new_n278), .ZN(new_n966));
  INV_X1    g765(.A(new_n916), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n963), .A2(new_n964), .A3(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(G197gat), .ZN(new_n970));
  NOR3_X1   g769(.A1(new_n969), .A2(new_n970), .A3(new_n704), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n899), .A2(new_n384), .ZN(new_n972));
  XOR2_X1   g771(.A(new_n972), .B(KEYINPUT123), .Z(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(new_n939), .ZN(new_n974));
  OR2_X1    g773(.A1(new_n974), .A2(KEYINPUT124), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(KEYINPUT124), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n975), .A2(new_n663), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n971), .B1(new_n970), .B2(new_n977), .ZN(G1352gat));
  XOR2_X1   g777(.A(KEYINPUT126), .B(G204gat), .Z(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  NOR3_X1   g779(.A1(new_n974), .A2(new_n633), .A3(new_n980), .ZN(new_n981));
  XNOR2_X1  g780(.A(new_n981), .B(KEYINPUT62), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n980), .B1(new_n969), .B2(new_n633), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(new_n983), .ZN(G1353gat));
  OAI211_X1 g783(.A(new_n605), .B(new_n964), .C1(new_n966), .C2(new_n967), .ZN(new_n985));
  AOI21_X1  g784(.A(KEYINPUT63), .B1(new_n985), .B2(G211gat), .ZN(new_n986));
  INV_X1    g785(.A(new_n986), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n985), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n987), .A2(KEYINPUT127), .A3(new_n988), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n986), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n510), .A2(G211gat), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n975), .A2(new_n976), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n989), .A2(new_n991), .A3(new_n993), .ZN(G1354gat));
  INV_X1    g793(.A(G218gat), .ZN(new_n995));
  NOR3_X1   g794(.A1(new_n969), .A2(new_n995), .A3(new_n606), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n975), .A2(new_n603), .A3(new_n976), .ZN(new_n997));
  AOI21_X1  g796(.A(new_n996), .B1(new_n995), .B2(new_n997), .ZN(G1355gat));
endmodule


