//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 1 1 1 1 0 0 0 1 1 0 0 1 0 0 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 0 1 0 1 1 1 0 0 0 1 1 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT64), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n209));
  INV_X1    g0009(.A(G232), .ZN(new_n210));
  INV_X1    g0010(.A(G97), .ZN(new_n211));
  INV_X1    g0011(.A(G257), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n209), .B1(new_n202), .B2(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n208), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT1), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n208), .A2(G13), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT0), .Z(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n202), .A2(new_n203), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G50), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n218), .B(new_n221), .C1(new_n224), .C2(new_n227), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(G226), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G68), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n202), .ZN(new_n243));
  XOR2_X1   g0043(.A(KEYINPUT66), .B(G50), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n241), .B(new_n245), .Z(G351));
  INV_X1    g0046(.A(G33), .ZN(new_n247));
  AOI21_X1  g0047(.A(G20), .B1(new_n247), .B2(G97), .ZN(new_n248));
  AND3_X1   g0048(.A1(KEYINPUT86), .A2(G33), .A3(G283), .ZN(new_n249));
  AOI21_X1  g0049(.A(KEYINPUT86), .B1(G33), .B2(G283), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G116), .ZN(new_n253));
  AOI22_X1  g0053(.A1(new_n252), .A2(new_n222), .B1(G20), .B2(new_n253), .ZN(new_n254));
  AND3_X1   g0054(.A1(new_n251), .A2(KEYINPUT20), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(KEYINPUT20), .B1(new_n251), .B2(new_n254), .ZN(new_n256));
  INV_X1    g0056(.A(G13), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G1), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(KEYINPUT71), .A3(G20), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G13), .A3(G20), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT71), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  OAI22_X1  g0064(.A1(new_n255), .A2(new_n256), .B1(G116), .B2(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n252), .A2(new_n222), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT73), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n264), .A2(KEYINPUT73), .A3(new_n266), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n253), .B1(new_n260), .B2(G33), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n265), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G200), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G1), .A3(G13), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n276), .A2(G274), .ZN(new_n277));
  INV_X1    g0077(.A(G45), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(G1), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT88), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n279), .B(new_n280), .C1(KEYINPUT5), .C2(new_n281), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n260), .B(G45), .C1(new_n281), .C2(KEYINPUT5), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT88), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n281), .A2(KEYINPUT5), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n277), .A2(new_n282), .A3(new_n284), .A4(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n285), .ZN(new_n287));
  OAI211_X1 g0087(.A(G270), .B(new_n276), .C1(new_n287), .C2(new_n283), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  AND2_X1   g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NOR2_X1   g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G303), .ZN(new_n293));
  OAI211_X1 g0093(.A(G264), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n294));
  INV_X1    g0094(.A(G1698), .ZN(new_n295));
  OAI211_X1 g0095(.A(G257), .B(new_n295), .C1(new_n290), .C2(new_n291), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n293), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n276), .B1(new_n297), .B2(KEYINPUT90), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT90), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n293), .A2(new_n299), .A3(new_n294), .A4(new_n296), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n289), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n273), .B(KEYINPUT91), .C1(new_n274), .C2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT91), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n297), .A2(KEYINPUT90), .ZN(new_n304));
  INV_X1    g0104(.A(new_n276), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n304), .A2(new_n300), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n289), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n274), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT73), .B1(new_n264), .B2(new_n266), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n252), .A2(new_n222), .ZN(new_n310));
  AOI211_X1 g0110(.A(new_n268), .B(new_n310), .C1(new_n259), .C2(new_n263), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n272), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n251), .A2(new_n254), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT20), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n251), .A2(KEYINPUT20), .A3(new_n254), .ZN(new_n316));
  INV_X1    g0116(.A(new_n264), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n315), .A2(new_n316), .B1(new_n253), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n303), .B1(new_n308), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n301), .A2(G190), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n302), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n306), .A2(new_n307), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n323), .A2(new_n319), .A3(G169), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT21), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n323), .A2(new_n319), .A3(KEYINPUT21), .A4(G169), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n306), .A2(G179), .A3(new_n307), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n319), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n326), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n322), .A2(new_n330), .ZN(new_n331));
  XOR2_X1   g0131(.A(KEYINPUT8), .B(G58), .Z(new_n332));
  NAND2_X1  g0132(.A1(new_n223), .A2(G33), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(G20), .A2(G33), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n332), .A2(new_n334), .B1(G150), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n204), .A2(G20), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n266), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT68), .ZN(new_n339));
  INV_X1    g0139(.A(new_n261), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n340), .A2(new_n310), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n223), .A2(G1), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n342), .A2(new_n201), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n341), .A2(new_n343), .B1(new_n201), .B2(new_n340), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n338), .A2(KEYINPUT68), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT9), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n347), .B(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n351), .A2(new_n276), .A3(G274), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n276), .A2(new_n350), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n353), .B1(G226), .B2(new_n355), .ZN(new_n356));
  OR2_X1    g0156(.A1(KEYINPUT3), .A2(G33), .ZN(new_n357));
  NAND2_X1  g0157(.A1(KEYINPUT3), .A2(G33), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G1698), .ZN(new_n360));
  INV_X1    g0160(.A(G223), .ZN(new_n361));
  INV_X1    g0161(.A(G77), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n360), .A2(new_n361), .B1(new_n362), .B2(new_n359), .ZN(new_n363));
  AOI21_X1  g0163(.A(G1698), .B1(new_n357), .B2(new_n358), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n363), .B1(G222), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n356), .B1(new_n365), .B2(new_n276), .ZN(new_n366));
  INV_X1    g0166(.A(G190), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(G200), .B2(new_n366), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n349), .A2(new_n369), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n370), .B(KEYINPUT10), .ZN(new_n371));
  INV_X1    g0171(.A(G169), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n347), .B1(new_n372), .B2(new_n366), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(G179), .B2(new_n366), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G226), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n295), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n210), .A2(G1698), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n377), .B(new_n378), .C1(new_n290), .C2(new_n291), .ZN(new_n379));
  NAND2_X1  g0179(.A1(G33), .A2(G97), .ZN(new_n380));
  AND3_X1   g0180(.A1(new_n379), .A2(KEYINPUT74), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT74), .B1(new_n379), .B2(new_n380), .ZN(new_n382));
  NOR3_X1   g0182(.A1(new_n381), .A2(new_n382), .A3(new_n276), .ZN(new_n383));
  INV_X1    g0183(.A(G238), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n352), .B1(new_n354), .B2(new_n384), .ZN(new_n385));
  NOR4_X1   g0185(.A1(new_n383), .A2(KEYINPUT75), .A3(KEYINPUT13), .A4(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT75), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n379), .A2(new_n380), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT74), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n276), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n379), .A2(KEYINPUT74), .A3(new_n380), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n385), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT13), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n387), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n386), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT76), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n392), .B2(new_n393), .ZN(new_n397));
  OAI211_X1 g0197(.A(KEYINPUT76), .B(KEYINPUT13), .C1(new_n383), .C2(new_n385), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(G200), .B1(new_n395), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT13), .B1(new_n383), .B2(new_n385), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n390), .A2(new_n391), .ZN(new_n402));
  INV_X1    g0202(.A(new_n385), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(new_n393), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n401), .A2(G190), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT77), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n401), .A2(new_n404), .A3(KEYINPUT77), .A4(G190), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n203), .A2(G20), .ZN(new_n410));
  INV_X1    g0210(.A(new_n335), .ZN(new_n411));
  OAI221_X1 g0211(.A(new_n410), .B1(new_n333), .B2(new_n362), .C1(new_n411), .C2(new_n201), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n310), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n413), .B(KEYINPUT11), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT12), .B1(new_n264), .B2(G68), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT12), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n258), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n415), .B1(new_n410), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  AOI211_X1 g0219(.A(new_n203), .B(new_n342), .C1(new_n269), .C2(new_n270), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n400), .A2(new_n409), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT78), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n400), .A2(new_n409), .A3(KEYINPUT78), .A4(new_n421), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n421), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n397), .B(new_n398), .C1(new_n386), .C2(new_n394), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT14), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n428), .A2(new_n429), .A3(G169), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n401), .A2(G179), .A3(new_n404), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n429), .B1(new_n428), .B2(G169), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n427), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n426), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT81), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n364), .A2(new_n436), .A3(G223), .ZN(new_n437));
  OAI211_X1 g0237(.A(G223), .B(new_n295), .C1(new_n290), .C2(new_n291), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT81), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(G87), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n247), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n292), .A2(new_n295), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n442), .B1(new_n443), .B2(G226), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n276), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n352), .B1(new_n354), .B2(new_n210), .ZN(new_n446));
  OAI21_X1  g0246(.A(G169), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n446), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n359), .A2(G226), .A3(G1698), .ZN(new_n449));
  INV_X1    g0249(.A(new_n442), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n451), .B1(new_n437), .B2(new_n439), .ZN(new_n452));
  OAI211_X1 g0252(.A(G179), .B(new_n448), .C1(new_n452), .C2(new_n276), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT82), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n447), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n454), .B1(new_n447), .B2(new_n453), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT18), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G58), .A2(G68), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n225), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G20), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT79), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n335), .A2(G159), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n223), .B1(new_n225), .B2(new_n460), .ZN(new_n466));
  INV_X1    g0266(.A(new_n464), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT79), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT7), .ZN(new_n470));
  NOR3_X1   g0270(.A1(new_n359), .A2(new_n470), .A3(G20), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT7), .B1(new_n292), .B2(new_n223), .ZN(new_n472));
  OAI21_X1  g0272(.A(G68), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n469), .A2(new_n473), .A3(KEYINPUT16), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT16), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n470), .B1(new_n359), .B2(G20), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n292), .A2(KEYINPUT7), .A3(new_n223), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n203), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n462), .A2(new_n464), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n474), .A2(new_n480), .A3(new_n310), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT80), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT80), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n474), .A2(new_n480), .A3(new_n483), .A4(new_n310), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n332), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(new_n342), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n487), .A2(new_n341), .B1(new_n340), .B2(new_n486), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n458), .A2(new_n459), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n447), .A2(new_n453), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(KEYINPUT82), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n455), .ZN(new_n493));
  INV_X1    g0293(.A(new_n488), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n494), .B1(new_n482), .B2(new_n484), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT18), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n274), .B1(new_n445), .B2(new_n446), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n448), .B1(new_n452), .B2(new_n276), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n497), .B1(new_n498), .B2(G190), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n485), .A2(new_n488), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT17), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n495), .A2(KEYINPUT17), .A3(new_n499), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n490), .A2(new_n496), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n353), .B1(G244), .B2(new_n355), .ZN(new_n505));
  INV_X1    g0305(.A(G107), .ZN(new_n506));
  OAI22_X1  g0306(.A1(new_n360), .A2(new_n384), .B1(new_n506), .B2(new_n359), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT69), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n364), .A2(new_n508), .A3(G232), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n364), .A2(G232), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT69), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n507), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n505), .B1(new_n512), .B2(new_n276), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G200), .ZN(new_n514));
  XNOR2_X1  g0314(.A(KEYINPUT15), .B(G87), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT70), .ZN(new_n516));
  XNOR2_X1  g0316(.A(new_n515), .B(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n517), .A2(new_n333), .ZN(new_n518));
  OAI22_X1  g0318(.A1(new_n486), .A2(new_n411), .B1(new_n223), .B2(new_n362), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n310), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n264), .A2(G77), .ZN(new_n521));
  XNOR2_X1  g0321(.A(new_n521), .B(KEYINPUT72), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n342), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n271), .A2(G77), .A3(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(G190), .B(new_n505), .C1(new_n512), .C2(new_n276), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n514), .A2(new_n523), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n513), .A2(new_n372), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n525), .A2(new_n520), .A3(new_n522), .ZN(new_n529));
  INV_X1    g0329(.A(G179), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n530), .B(new_n505), .C1(new_n512), .C2(new_n276), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n528), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  NOR4_X1   g0333(.A1(new_n375), .A2(new_n435), .A3(new_n504), .A4(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n260), .A2(G33), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n266), .A2(G107), .A3(new_n261), .A4(new_n535), .ZN(new_n536));
  OR3_X1    g0336(.A1(new_n261), .A2(KEYINPUT25), .A3(G107), .ZN(new_n537));
  OAI21_X1  g0337(.A(KEYINPUT25), .B1(new_n261), .B2(G107), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT93), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT93), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n536), .A2(new_n541), .A3(new_n537), .A4(new_n538), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT23), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n223), .B2(G107), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n506), .A2(KEYINPUT23), .A3(G20), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n247), .A2(new_n253), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n223), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT92), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n551), .A2(new_n223), .A3(G87), .ZN(new_n552));
  OAI21_X1  g0352(.A(KEYINPUT22), .B1(new_n292), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT22), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n441), .A2(KEYINPUT92), .A3(G20), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n359), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n550), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n310), .B1(new_n557), .B2(KEYINPUT24), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n547), .A2(new_n549), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n292), .A2(KEYINPUT22), .A3(new_n552), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n554), .B1(new_n359), .B2(new_n555), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT24), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n543), .B1(new_n558), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(G264), .B(new_n276), .C1(new_n287), .C2(new_n283), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(G257), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n568));
  OAI211_X1 g0368(.A(G250), .B(new_n295), .C1(new_n290), .C2(new_n291), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G33), .A2(G294), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n567), .B1(new_n305), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n286), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n372), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n530), .A3(new_n286), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n565), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n562), .A2(new_n563), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n557), .A2(KEYINPUT24), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n577), .A2(new_n578), .A3(new_n310), .ZN(new_n579));
  AOI21_X1  g0379(.A(G200), .B1(new_n572), .B2(new_n286), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n571), .A2(new_n305), .ZN(new_n581));
  AND4_X1   g0381(.A1(new_n367), .A2(new_n581), .A3(new_n286), .A4(new_n566), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n579), .B(new_n543), .C1(new_n580), .C2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n576), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT94), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT94), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n576), .A2(new_n583), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT6), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n211), .A2(new_n506), .ZN(new_n590));
  NOR2_X1   g0390(.A1(G97), .A2(G107), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n506), .A2(KEYINPUT84), .A3(KEYINPUT6), .A4(G97), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT84), .ZN(new_n594));
  NAND2_X1  g0394(.A1(KEYINPUT6), .A2(G97), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n594), .B1(new_n595), .B2(G107), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n592), .A2(new_n593), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G20), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT83), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n411), .B2(new_n362), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n335), .A2(KEYINPUT83), .A3(G77), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n598), .A2(KEYINPUT85), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n506), .B1(new_n476), .B2(new_n477), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n597), .A2(G20), .B1(new_n600), .B2(new_n601), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(KEYINPUT85), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n310), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n340), .A2(new_n211), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n266), .A2(new_n261), .A3(new_n535), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n610), .B1(new_n611), .B2(new_n211), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  OAI211_X1 g0413(.A(G250), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT87), .ZN(new_n615));
  XNOR2_X1  g0415(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n364), .A2(KEYINPUT4), .A3(G244), .ZN(new_n617));
  OAI211_X1 g0417(.A(G244), .B(new_n295), .C1(new_n290), .C2(new_n291), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT4), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OR2_X1    g0420(.A1(new_n249), .A2(new_n250), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n617), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n305), .B1(new_n616), .B2(new_n622), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n276), .B(G257), .C1(new_n283), .C2(new_n287), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n286), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n623), .A2(new_n367), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(G200), .B1(new_n623), .B2(new_n626), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n609), .B(new_n613), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n623), .A2(new_n626), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n372), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n623), .A2(new_n530), .A3(new_n626), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n604), .B1(new_n607), .B2(KEYINPUT85), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n598), .A2(new_n602), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT85), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n266), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n631), .B(new_n632), .C1(new_n637), .C2(new_n612), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n359), .A2(G244), .A3(G1698), .ZN(new_n639));
  INV_X1    g0439(.A(new_n548), .ZN(new_n640));
  OAI211_X1 g0440(.A(G238), .B(new_n295), .C1(new_n290), .C2(new_n291), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n305), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n260), .A2(G45), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(G250), .ZN(new_n645));
  OAI21_X1  g0445(.A(KEYINPUT89), .B1(new_n305), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT89), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n276), .A2(new_n647), .A3(G250), .A4(new_n644), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n646), .A2(new_n648), .B1(new_n279), .B2(new_n277), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n643), .A2(new_n649), .A3(new_n530), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n517), .A2(new_n317), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT19), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n223), .B1(new_n380), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n591), .A2(new_n441), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n652), .B1(new_n333), .B2(new_n211), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n223), .A2(G68), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n655), .B(new_n656), .C1(new_n292), .C2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n310), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n651), .B(new_n659), .C1(new_n611), .C2(new_n517), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n643), .A2(new_n649), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n650), .B(new_n660), .C1(new_n661), .C2(G169), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n643), .A2(new_n649), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(G200), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n341), .A2(G87), .A3(new_n535), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n651), .A2(new_n659), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n643), .A2(new_n649), .A3(G190), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n664), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n629), .A2(new_n638), .A3(new_n669), .ZN(new_n670));
  AND4_X1   g0470(.A1(new_n331), .A2(new_n534), .A3(new_n588), .A4(new_n670), .ZN(G372));
  AND2_X1   g0471(.A1(new_n502), .A2(new_n503), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n532), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n426), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n673), .B1(new_n675), .B2(new_n434), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n459), .B1(new_n489), .B2(new_n491), .ZN(new_n677));
  INV_X1    g0477(.A(new_n491), .ZN(new_n678));
  NOR3_X1   g0478(.A1(new_n495), .A2(KEYINPUT18), .A3(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n371), .B1(new_n676), .B2(new_n681), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n682), .A2(new_n374), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n638), .A2(new_n629), .A3(new_n669), .A4(new_n583), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT95), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n583), .A2(new_n662), .A3(new_n668), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n687), .A2(KEYINPUT95), .A3(new_n638), .A4(new_n629), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n326), .A2(new_n327), .A3(new_n329), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n576), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n686), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n609), .A2(new_n613), .ZN(new_n692));
  AOI21_X1  g0492(.A(G169), .B1(new_n623), .B2(new_n626), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n614), .B(KEYINPUT87), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n694), .A2(new_n621), .A3(new_n617), .A4(new_n620), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n625), .B1(new_n695), .B2(new_n305), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n693), .B1(new_n530), .B2(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n669), .A2(KEYINPUT26), .A3(new_n692), .A4(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(KEYINPUT96), .ZN(new_n699));
  INV_X1    g0499(.A(new_n638), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT96), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n700), .A2(new_n701), .A3(KEYINPUT26), .A4(new_n669), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT26), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n662), .A2(new_n668), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n703), .B1(new_n638), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n699), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n691), .A2(new_n662), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n534), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n683), .A2(new_n708), .ZN(G369));
  NAND2_X1  g0509(.A1(new_n258), .A2(new_n223), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n710), .A2(KEYINPUT27), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(KEYINPUT27), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n711), .A2(G213), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G343), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT97), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n714), .B(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(new_n273), .ZN(new_n718));
  MUX2_X1   g0518(.A(new_n331), .B(new_n330), .S(new_n718), .Z(new_n719));
  XNOR2_X1  g0519(.A(KEYINPUT98), .B(G330), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n716), .A2(new_n565), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n588), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(new_n576), .B2(new_n717), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n330), .A2(new_n717), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n588), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n576), .A2(new_n716), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n725), .A2(new_n731), .ZN(G399));
  INV_X1    g0532(.A(new_n219), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G41), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n591), .A2(new_n441), .A3(new_n253), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n734), .A2(new_n260), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n736), .B1(new_n227), .B2(new_n734), .ZN(new_n737));
  XOR2_X1   g0537(.A(new_n737), .B(KEYINPUT28), .Z(new_n738));
  AND2_X1   g0538(.A1(new_n629), .A2(new_n638), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n690), .A2(new_n739), .A3(new_n687), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n662), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n705), .A2(new_n698), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n717), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT29), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n707), .A2(new_n717), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n745), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT30), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n661), .A2(new_n572), .A3(new_n623), .A4(new_n626), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n301), .A2(G179), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n661), .A2(G179), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n752), .A2(new_n323), .A3(new_n630), .A4(new_n573), .ZN(new_n753));
  AND2_X1   g0553(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n754), .A2(KEYINPUT99), .ZN(new_n755));
  AND3_X1   g0555(.A1(new_n572), .A2(new_n643), .A3(new_n649), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n328), .A2(new_n696), .A3(KEYINPUT30), .A4(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(new_n754), .B2(KEYINPUT99), .ZN(new_n758));
  OAI211_X1 g0558(.A(KEYINPUT31), .B(new_n716), .C1(new_n755), .C2(new_n758), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n331), .A2(new_n588), .A3(new_n670), .A4(new_n717), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n751), .A2(new_n753), .A3(new_n757), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n716), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT31), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n759), .A2(new_n760), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n747), .B1(new_n720), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n738), .B1(new_n766), .B2(G1), .ZN(G364));
  NOR2_X1   g0567(.A1(new_n257), .A2(G20), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n260), .B1(new_n768), .B2(G45), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n734), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n721), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(new_n720), .B2(new_n719), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n223), .B1(KEYINPUT101), .B2(new_n372), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n372), .A2(KEYINPUT101), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n222), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n223), .A2(new_n530), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n367), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n223), .A2(G179), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G190), .A2(G200), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G159), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n781), .A2(new_n201), .B1(new_n786), .B2(KEYINPUT32), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n779), .A2(G190), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n782), .A2(G190), .A3(G200), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n789), .A2(new_n203), .B1(new_n790), .B2(new_n441), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n367), .A2(G200), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n223), .B1(new_n793), .B2(new_n530), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT102), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G97), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n778), .A2(new_n793), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n359), .B1(new_n797), .B2(new_n202), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n778), .A2(new_n783), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n798), .B1(G77), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n782), .A2(new_n367), .A3(G200), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n786), .A2(KEYINPUT32), .B1(G107), .B2(new_n803), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n792), .A2(new_n796), .A3(new_n801), .A4(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G322), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n797), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G311), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n292), .B1(new_n799), .B2(new_n808), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n807), .B(new_n809), .C1(G329), .C2(new_n785), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n780), .A2(G326), .ZN(new_n811));
  XNOR2_X1  g0611(.A(KEYINPUT33), .B(G317), .ZN(new_n812));
  INV_X1    g0612(.A(new_n790), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n788), .A2(new_n812), .B1(new_n813), .B2(G303), .ZN(new_n814));
  INV_X1    g0614(.A(new_n794), .ZN(new_n815));
  AOI22_X1  g0615(.A1(G294), .A2(new_n815), .B1(new_n803), .B2(G283), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n810), .A2(new_n811), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n777), .B1(new_n805), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(G13), .A2(G33), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(G20), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n776), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n219), .A2(new_n292), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(new_n278), .B2(new_n227), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n245), .B2(new_n278), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n219), .A2(G116), .ZN(new_n827));
  INV_X1    g0627(.A(G355), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT100), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n359), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(new_n829), .B2(new_n828), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n827), .B1(new_n219), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n823), .B1(new_n826), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n771), .ZN(new_n834));
  NOR3_X1   g0634(.A1(new_n818), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n821), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n835), .B1(new_n719), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n773), .A2(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT103), .Z(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(G396));
  OAI22_X1  g0640(.A1(new_n799), .A2(new_n253), .B1(new_n784), .B2(new_n808), .ZN(new_n841));
  INV_X1    g0641(.A(new_n797), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n359), .B(new_n841), .C1(G294), .C2(new_n842), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n780), .A2(G303), .B1(new_n813), .B2(G107), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n802), .A2(new_n441), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(G283), .B2(new_n788), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n843), .A2(new_n796), .A3(new_n844), .A4(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(G132), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n359), .B1(new_n784), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G68), .B2(new_n803), .ZN(new_n850));
  AOI22_X1  g0650(.A1(G58), .A2(new_n815), .B1(new_n813), .B2(G50), .ZN(new_n851));
  AOI22_X1  g0651(.A1(G143), .A2(new_n842), .B1(new_n800), .B2(G159), .ZN(new_n852));
  INV_X1    g0652(.A(G137), .ZN(new_n853));
  INV_X1    g0653(.A(G150), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n852), .B1(new_n781), .B2(new_n853), .C1(new_n854), .C2(new_n789), .ZN(new_n855));
  XNOR2_X1  g0655(.A(KEYINPUT104), .B(KEYINPUT34), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n850), .B(new_n851), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n855), .A2(new_n856), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n847), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n776), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n776), .A2(new_n819), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n834), .B1(new_n362), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n716), .A2(new_n529), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n527), .A2(new_n532), .A3(new_n863), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n716), .A2(new_n531), .A3(new_n528), .A4(new_n529), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT105), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n865), .A2(KEYINPUT105), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n864), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n860), .B(new_n862), .C1(new_n869), .C2(new_n820), .ZN(new_n870));
  OR2_X1    g0670(.A1(new_n865), .A2(KEYINPUT105), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n527), .A2(new_n532), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n871), .A2(new_n866), .B1(new_n872), .B2(new_n863), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n746), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n873), .A2(new_n716), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n707), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n765), .A2(new_n720), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n771), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n877), .A2(new_n878), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n870), .B1(new_n880), .B2(new_n881), .ZN(G384));
  NOR2_X1   g0682(.A1(new_n768), .A2(new_n260), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n761), .A2(KEYINPUT31), .A3(new_n716), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT31), .B1(new_n761), .B2(new_n716), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n873), .B1(new_n887), .B2(new_n760), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n427), .A2(new_n716), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n426), .A2(new_n434), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n889), .B1(new_n426), .B2(new_n434), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(KEYINPUT110), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n469), .A2(new_n473), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n475), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(new_n310), .A3(new_n474), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n488), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n713), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n504), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT37), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n897), .A2(new_n491), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n500), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n899), .B1(new_n903), .B2(KEYINPUT108), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT108), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n500), .A2(new_n905), .A3(new_n902), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n901), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n901), .B1(new_n493), .B2(new_n495), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n485), .A2(new_n488), .A3(new_n499), .ZN(new_n909));
  INV_X1    g0709(.A(new_n713), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n495), .A2(new_n910), .ZN(new_n911));
  NOR3_X1   g0711(.A1(new_n908), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  OAI211_X1 g0712(.A(KEYINPUT38), .B(new_n900), .C1(new_n907), .C2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT38), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n489), .A2(new_n713), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n672), .B2(new_n680), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n489), .A2(new_n491), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(new_n915), .A3(new_n500), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n909), .A2(new_n911), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT37), .B1(new_n458), .B2(new_n489), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n918), .A2(KEYINPUT37), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n914), .B1(new_n916), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n913), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT110), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n888), .B(new_n924), .C1(new_n890), .C2(new_n891), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n893), .A2(KEYINPUT40), .A3(new_n923), .A4(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT111), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n925), .A2(KEYINPUT40), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n929), .A2(KEYINPUT111), .A3(new_n923), .A4(new_n893), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n903), .A2(KEYINPUT108), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(new_n906), .A3(new_n898), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n912), .B1(new_n933), .B2(KEYINPUT37), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n504), .A2(new_n899), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n914), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n892), .B1(new_n936), .B2(new_n913), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n931), .B1(KEYINPUT40), .B2(new_n937), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n938), .B(KEYINPUT112), .Z(new_n939));
  NAND2_X1  g0739(.A1(new_n887), .A2(new_n760), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n534), .A2(new_n940), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n941), .B(KEYINPUT113), .Z(new_n942));
  OR2_X1    g0742(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n939), .A2(new_n942), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n943), .A2(new_n944), .A3(new_n720), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT39), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n923), .A2(new_n946), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n434), .A2(new_n716), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n936), .A2(KEYINPUT39), .A3(new_n913), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n947), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n936), .A2(new_n913), .ZN(new_n952));
  INV_X1    g0752(.A(new_n889), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n435), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n426), .A2(new_n434), .A3(new_n889), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n532), .A2(new_n716), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(KEYINPUT107), .B1(new_n876), .B2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT107), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n960), .B(new_n957), .C1(new_n707), .C2(new_n875), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n952), .B(new_n956), .C1(new_n959), .C2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n681), .A2(new_n910), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n951), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(KEYINPUT109), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT109), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n951), .A2(new_n962), .A3(new_n966), .A4(new_n963), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n747), .A2(new_n534), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n683), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n968), .B(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n883), .B1(new_n945), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n945), .B2(new_n971), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n597), .A2(KEYINPUT35), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n597), .A2(KEYINPUT35), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n974), .A2(G116), .A3(new_n224), .A4(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT36), .ZN(new_n977));
  AND3_X1   g0777(.A1(new_n227), .A2(G77), .A3(new_n460), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n203), .A2(G50), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT106), .Z(new_n980));
  OAI211_X1 g0780(.A(G1), .B(new_n257), .C1(new_n978), .C2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n973), .A2(new_n977), .A3(new_n981), .ZN(G367));
  NAND2_X1  g0782(.A1(new_n692), .A2(new_n716), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n739), .A2(new_n983), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n984), .A2(new_n576), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n716), .B1(new_n985), .B2(new_n638), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n700), .A2(new_n716), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n729), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n986), .B1(KEYINPUT42), .B2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT114), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n989), .A2(KEYINPUT42), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n990), .B2(new_n991), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n717), .A2(new_n666), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(new_n704), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n992), .A2(new_n994), .B1(KEYINPUT43), .B2(new_n997), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n999), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n988), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1002), .B1(new_n725), .B2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n725), .A2(new_n1003), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1000), .A2(new_n1005), .A3(new_n1001), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n734), .B(KEYINPUT41), .Z(new_n1007));
  NAND2_X1  g0807(.A1(new_n731), .A2(new_n988), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(KEYINPUT115), .B(KEYINPUT45), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1003), .B1(new_n729), .B2(new_n730), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1011), .A2(KEYINPUT116), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(KEYINPUT116), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1012), .A2(KEYINPUT44), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(KEYINPUT44), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(KEYINPUT117), .B2(new_n725), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n728), .B1(new_n724), .B2(new_n727), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n721), .B(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n725), .A2(KEYINPUT117), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1018), .A2(new_n766), .A3(new_n1020), .A4(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1007), .B1(new_n1023), .B2(new_n766), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1004), .B(new_n1006), .C1(new_n1024), .C2(new_n770), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n822), .B1(new_n219), .B2(new_n517), .C1(new_n824), .C2(new_n236), .ZN(new_n1026));
  AND2_X1   g0826(.A1(new_n1026), .A2(new_n771), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n797), .A2(new_n854), .B1(new_n799), .B2(new_n201), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n292), .B(new_n1028), .C1(G137), .C2(new_n785), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n795), .A2(G68), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n788), .A2(G159), .B1(new_n780), .B2(G143), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n802), .A2(new_n362), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(G58), .B2(new_n813), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n788), .A2(G294), .B1(new_n803), .B2(G97), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n506), .B2(new_n794), .C1(new_n808), .C2(new_n781), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G303), .A2(new_n842), .B1(new_n785), .B2(G317), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT46), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n790), .B2(new_n253), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n359), .B1(new_n800), .B2(G283), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n813), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1037), .A2(new_n1039), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1034), .B1(new_n1036), .B2(new_n1042), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT47), .Z(new_n1044));
  OAI221_X1 g0844(.A(new_n1027), .B1(new_n777), .B2(new_n1044), .C1(new_n997), .C2(new_n836), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1025), .A2(new_n1045), .ZN(G387));
  NAND2_X1  g0846(.A1(new_n1020), .A2(new_n770), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G303), .A2(new_n800), .B1(new_n842), .B2(G317), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n781), .B2(new_n806), .C1(new_n808), .C2(new_n789), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT48), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G283), .A2(new_n815), .B1(new_n813), .B2(G294), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT49), .Z(new_n1055));
  AOI21_X1  g0855(.A(new_n359), .B1(new_n785), .B2(G326), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n253), .B2(new_n802), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n517), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n795), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n797), .A2(new_n201), .B1(new_n784), .B2(new_n854), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n292), .B(new_n1061), .C1(G68), .C2(new_n800), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n788), .A2(new_n332), .B1(new_n803), .B2(G97), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n780), .A2(G159), .B1(new_n813), .B2(G77), .ZN(new_n1064));
  AND4_X1   g0864(.A1(new_n1060), .A2(new_n1062), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n776), .B1(new_n1058), .B2(new_n1065), .ZN(new_n1066));
  NOR3_X1   g0866(.A1(new_n233), .A2(new_n278), .A3(new_n359), .ZN(new_n1067));
  OR3_X1    g0867(.A1(new_n486), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1068));
  OAI21_X1  g0868(.A(KEYINPUT50), .B1(new_n486), .B2(G50), .ZN(new_n1069));
  AOI21_X1  g0869(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n735), .B1(new_n1071), .B2(new_n292), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n219), .B1(new_n1067), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n823), .B1(G107), .B2(new_n733), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n834), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1066), .B(new_n1075), .C1(new_n724), .C2(new_n836), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n766), .A2(new_n1020), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n766), .A2(new_n1020), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT118), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n734), .B(new_n1077), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1047), .B(new_n1076), .C1(new_n1080), .C2(new_n1081), .ZN(G393));
  OR2_X1    g0882(.A1(new_n1017), .A2(new_n725), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1017), .A2(new_n725), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n1077), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1086), .A2(new_n734), .A3(new_n1023), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1083), .A2(new_n1084), .A3(new_n770), .ZN(new_n1088));
  AND3_X1   g0888(.A1(new_n241), .A2(new_n219), .A3(new_n292), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n822), .B1(new_n219), .B2(new_n211), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n771), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(G159), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n781), .A2(new_n854), .B1(new_n1092), .B2(new_n797), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT51), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n795), .A2(G77), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n845), .B1(G50), .B2(new_n788), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n785), .A2(G143), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n292), .B1(new_n800), .B2(new_n332), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n813), .A2(G68), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n780), .A2(G317), .B1(new_n842), .B2(G311), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT52), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n292), .B1(new_n784), .B2(new_n806), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(G294), .B2(new_n800), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n788), .A2(G303), .B1(new_n803), .B2(G107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(G116), .A2(new_n815), .B1(new_n813), .B2(G283), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n1098), .A2(new_n1103), .B1(new_n1105), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1091), .B1(new_n776), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n988), .B2(new_n836), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1087), .A2(new_n1088), .A3(new_n1113), .ZN(G390));
  INV_X1    g0914(.A(KEYINPUT119), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n956), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n869), .A2(new_n717), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n662), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n684), .A2(new_n685), .B1(new_n689), .B2(new_n576), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1118), .B1(new_n1119), .B2(new_n688), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1117), .B1(new_n1120), .B2(new_n706), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n960), .B1(new_n1121), .B2(new_n957), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n876), .A2(KEYINPUT107), .A3(new_n958), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1116), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1115), .B1(new_n1124), .B2(new_n949), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n947), .A2(new_n950), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n956), .B1(new_n959), .B2(new_n961), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1127), .A2(KEYINPUT119), .A3(new_n948), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1125), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n878), .A2(new_n873), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n956), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n958), .B1(new_n743), .B2(new_n873), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n956), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1133), .A2(new_n923), .A3(new_n948), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1129), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1134), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n947), .A2(new_n950), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1127), .A2(new_n948), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1137), .B1(new_n1138), .B2(new_n1115), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1136), .B1(new_n1139), .B2(new_n1128), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n956), .A2(G330), .A3(new_n888), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1135), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1142), .A2(new_n769), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1126), .A2(new_n819), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n861), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n771), .B1(new_n332), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(G128), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n1147), .A2(new_n781), .B1(new_n789), .B2(new_n853), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(G50), .B2(new_n803), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT54), .B(G143), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n799), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n359), .B1(new_n797), .B2(new_n848), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1151), .B(new_n1152), .C1(G125), .C2(new_n785), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n795), .A2(G159), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n790), .A2(new_n854), .ZN(new_n1155));
  XOR2_X1   g0955(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n1156));
  XNOR2_X1  g0956(.A(new_n1155), .B(new_n1156), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1149), .A2(new_n1153), .A3(new_n1154), .A4(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1096), .B1(new_n253), .B2(new_n797), .ZN(new_n1159));
  XOR2_X1   g0959(.A(new_n1159), .B(KEYINPUT121), .Z(new_n1160));
  INV_X1    g0960(.A(G283), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n506), .A2(new_n789), .B1(new_n781), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(G294), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n292), .B1(new_n784), .B2(new_n1163), .C1(new_n211), .C2(new_n799), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n203), .A2(new_n802), .B1(new_n790), .B2(new_n441), .ZN(new_n1165));
  OR3_X1    g0965(.A1(new_n1162), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1158), .B1(new_n1160), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1146), .B1(new_n1167), .B2(new_n776), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1143), .B1(new_n1144), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1141), .B1(new_n1130), .B2(new_n956), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n959), .B2(new_n961), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n888), .A2(G330), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1132), .B1(new_n1116), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n1131), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n534), .A2(G330), .A3(new_n940), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n969), .A2(new_n1176), .A3(new_n683), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1175), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1142), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1177), .B1(new_n1171), .B2(new_n1174), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1135), .B(new_n1181), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1180), .A2(new_n734), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1169), .A2(new_n1183), .ZN(G378));
  OAI21_X1  g0984(.A(G330), .B1(new_n937), .B2(KEYINPUT40), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n931), .A2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n713), .B1(new_n345), .B2(new_n346), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT55), .Z(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n375), .B(new_n1190), .ZN(new_n1191));
  XOR2_X1   g0991(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n375), .B(new_n1189), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1192), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1193), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1187), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1197), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n931), .A2(new_n1186), .A3(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1198), .A2(new_n968), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n965), .A2(new_n967), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1197), .B(new_n1185), .C1(new_n928), .C2(new_n930), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1199), .B1(new_n931), .B2(new_n1186), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1202), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1201), .A2(new_n1205), .A3(KEYINPUT123), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1182), .A2(new_n1178), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT123), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1198), .A2(new_n968), .A3(new_n1208), .A4(new_n1200), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1206), .A2(new_n1207), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT57), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n734), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1211), .B1(new_n1201), .B2(new_n1205), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1213), .B1(new_n1214), .B2(new_n1207), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1212), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1206), .A2(new_n770), .A3(new_n1209), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n771), .B1(G50), .B2(new_n1145), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n359), .A2(G41), .ZN(new_n1219));
  AOI211_X1 g1019(.A(G50), .B(new_n1219), .C1(new_n247), .C2(new_n281), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1219), .B1(new_n1161), .B2(new_n784), .C1(new_n506), .C2(new_n797), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n1059), .B2(new_n800), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n813), .A2(G77), .B1(new_n803), .B2(G58), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n788), .A2(G97), .B1(new_n780), .B2(G116), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1222), .A2(new_n1030), .A3(new_n1223), .A4(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT58), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1220), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n795), .A2(G150), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n797), .A2(new_n1147), .B1(new_n799), .B2(new_n853), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(G132), .B2(new_n788), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1150), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n780), .A2(G125), .B1(new_n813), .B2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1228), .A2(new_n1230), .A3(new_n1232), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1233), .A2(KEYINPUT59), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(KEYINPUT59), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n803), .A2(G159), .ZN(new_n1236));
  AOI211_X1 g1036(.A(G33), .B(G41), .C1(new_n785), .C2(G124), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1227), .B1(new_n1226), .B2(new_n1225), .C1(new_n1234), .C2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1218), .B1(new_n1239), .B2(new_n776), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n1197), .B2(new_n820), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1217), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1216), .A2(new_n1242), .ZN(G375));
  AOI21_X1  g1043(.A(new_n834), .B1(new_n203), .B2(new_n861), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n359), .B1(new_n785), .B2(G303), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n1245), .B1(new_n506), .B2(new_n799), .C1(new_n1161), .C2(new_n797), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n781), .A2(new_n1163), .B1(new_n790), .B2(new_n211), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n789), .A2(new_n253), .ZN(new_n1248));
  NOR4_X1   g1048(.A1(new_n1246), .A2(new_n1247), .A3(new_n1032), .A4(new_n1248), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n789), .A2(new_n1150), .B1(new_n1092), .B2(new_n790), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n781), .A2(new_n848), .B1(new_n802), .B2(new_n202), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n359), .B1(new_n797), .B2(new_n853), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n799), .A2(new_n854), .B1(new_n784), .B2(new_n1147), .ZN(new_n1253));
  NOR4_X1   g1053(.A1(new_n1250), .A2(new_n1251), .A3(new_n1252), .A4(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n795), .A2(G50), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1249), .A2(new_n1060), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n1244), .B1(new_n777), .B2(new_n1256), .C1(new_n956), .C2(new_n820), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n1175), .B2(new_n770), .ZN(new_n1259));
  OR2_X1    g1059(.A1(new_n1181), .A2(new_n1007), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1177), .A2(new_n1171), .A3(new_n1174), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1259), .B1(new_n1260), .B2(new_n1262), .ZN(G381));
  INV_X1    g1063(.A(G390), .ZN(new_n1264));
  INV_X1    g1064(.A(G384), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  OR4_X1    g1066(.A1(G396), .A2(new_n1266), .A3(G393), .A4(G381), .ZN(new_n1267));
  OR4_X1    g1067(.A1(G387), .A2(new_n1267), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1068(.A(G378), .ZN(new_n1269));
  INV_X1    g1069(.A(G343), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(G213), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(new_n1271), .B(KEYINPUT124), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1269), .A2(new_n1216), .A3(new_n1242), .A4(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(G407), .A2(G213), .A3(new_n1273), .ZN(G409));
  NAND3_X1  g1074(.A1(new_n1216), .A2(G378), .A3(new_n1242), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1201), .A2(new_n1205), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n770), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1241), .B(new_n1277), .C1(new_n1210), .C2(new_n1007), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1269), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1275), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1272), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1262), .A2(new_n1179), .A3(KEYINPUT60), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT60), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1261), .B1(new_n1181), .B2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1282), .A2(new_n1284), .A3(new_n734), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1285), .A2(G384), .A3(new_n1259), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(G384), .B1(new_n1285), .B2(new_n1259), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1280), .A2(new_n1281), .A3(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT63), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(G390), .A2(new_n1025), .A3(new_n1045), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT126), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(G393), .B(new_n839), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(G387), .A2(new_n1264), .ZN(new_n1297));
  AOI22_X1  g1097(.A1(new_n1295), .A2(new_n1296), .B1(new_n1297), .B2(new_n1293), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT61), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1297), .A2(KEYINPUT126), .A3(new_n1293), .A4(new_n1296), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1299), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1288), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1304), .A2(G2897), .A3(new_n1272), .A4(new_n1286), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1272), .A2(G2897), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1306), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1305), .A2(KEYINPUT125), .A3(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(KEYINPUT125), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1303), .A2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1272), .B1(new_n1275), .B2(new_n1279), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1312), .A2(KEYINPUT63), .A3(new_n1289), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1292), .A2(new_n1302), .A3(new_n1311), .A4(new_n1313), .ZN(new_n1314));
  AND2_X1   g1114(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1300), .B1(new_n1312), .B2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT62), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1290), .A2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1312), .A2(KEYINPUT62), .A3(new_n1289), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1316), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1299), .A2(new_n1301), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT127), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1299), .A2(KEYINPUT127), .A3(new_n1301), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1314), .B1(new_n1320), .B2(new_n1325), .ZN(G405));
  INV_X1    g1126(.A(new_n1275), .ZN(new_n1327));
  AOI21_X1  g1127(.A(G378), .B1(new_n1216), .B2(new_n1242), .ZN(new_n1328));
  OR3_X1    g1128(.A1(new_n1327), .A2(new_n1289), .A3(new_n1328), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1289), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n1321), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1329), .A2(new_n1301), .A3(new_n1299), .A4(new_n1330), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(G402));
endmodule


