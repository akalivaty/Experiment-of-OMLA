

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n618, n619, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781;

  INV_X1 U373 ( .A(n658), .ZN(n356) );
  INV_X1 U374 ( .A(KEYINPUT60), .ZN(n354) );
  INV_X1 U375 ( .A(KEYINPUT56), .ZN(n358) );
  XNOR2_X1 U376 ( .A(n431), .B(n430), .ZN(n777) );
  XNOR2_X1 U377 ( .A(n351), .B(n350), .ZN(n778) );
  INV_X1 U378 ( .A(KEYINPUT111), .ZN(n350) );
  XNOR2_X1 U379 ( .A(n627), .B(n360), .ZN(n384) );
  NOR2_X1 U380 ( .A1(n624), .A2(n623), .ZN(n625) );
  INV_X1 U381 ( .A(n408), .ZN(n360) );
  INV_X1 U382 ( .A(n608), .ZN(n586) );
  XNOR2_X1 U383 ( .A(n463), .B(KEYINPUT38), .ZN(n434) );
  INV_X1 U384 ( .A(KEYINPUT109), .ZN(n353) );
  NAND2_X1 U385 ( .A1(n363), .A2(n362), .ZN(n592) );
  INV_X1 U386 ( .A(n693), .ZN(n363) );
  XOR2_X1 U387 ( .A(G131), .B(G140), .Z(n525) );
  INV_X1 U388 ( .A(KEYINPUT4), .ZN(n474) );
  BUF_X1 U389 ( .A(n433), .Z(n463) );
  INV_X2 U390 ( .A(n748), .ZN(n364) );
  XNOR2_X2 U391 ( .A(n653), .B(KEYINPUT68), .ZN(n654) );
  NAND2_X1 U392 ( .A1(n479), .A2(n477), .ZN(n655) );
  BUF_X2 U393 ( .A(n738), .Z(n743) );
  AND2_X1 U394 ( .A1(n619), .A2(n412), .ZN(n351) );
  NAND2_X2 U395 ( .A1(n481), .A2(n480), .ZN(n489) );
  NAND2_X1 U396 ( .A1(n452), .A2(n352), .ZN(n650) );
  XNOR2_X1 U397 ( .A(n616), .B(n353), .ZN(n352) );
  XNOR2_X1 U398 ( .A(n355), .B(n354), .ZN(G60) );
  NAND2_X1 U399 ( .A1(n462), .A2(n364), .ZN(n355) );
  XNOR2_X1 U400 ( .A(n357), .B(n356), .ZN(G57) );
  NAND2_X1 U401 ( .A1(n371), .A2(n364), .ZN(n357) );
  XNOR2_X1 U402 ( .A(n359), .B(n358), .ZN(G51) );
  NAND2_X1 U403 ( .A1(n369), .A2(n364), .ZN(n359) );
  XNOR2_X2 U404 ( .A(n737), .B(KEYINPUT59), .ZN(n416) );
  INV_X1 U405 ( .A(n384), .ZN(n636) );
  NAND2_X1 U406 ( .A1(n365), .A2(n384), .ZN(n383) );
  XNOR2_X2 U407 ( .A(n655), .B(KEYINPUT86), .ZN(n767) );
  NAND2_X2 U408 ( .A1(n688), .A2(n685), .ZN(n646) );
  XNOR2_X2 U409 ( .A(n419), .B(n418), .ZN(n688) );
  XNOR2_X1 U410 ( .A(G131), .B(KEYINPUT75), .ZN(n556) );
  XNOR2_X1 U411 ( .A(G143), .B(G104), .ZN(n532) );
  NAND2_X1 U412 ( .A1(n597), .A2(n598), .ZN(n672) );
  XNOR2_X1 U413 ( .A(KEYINPUT91), .B(KEYINPUT0), .ZN(n361) );
  XOR2_X1 U414 ( .A(n694), .B(KEYINPUT98), .Z(n362) );
  NOR2_X1 U415 ( .A1(n585), .A2(n597), .ZN(n685) );
  XNOR2_X1 U416 ( .A(n580), .B(n579), .ZN(n693) );
  NOR2_X1 U417 ( .A1(n745), .A2(G902), .ZN(n580) );
  XNOR2_X1 U418 ( .A(n374), .B(n600), .ZN(n757) );
  AND2_X1 U419 ( .A1(n685), .A2(n362), .ZN(n390) );
  NAND2_X1 U420 ( .A1(n586), .A2(n366), .ZN(n386) );
  XNOR2_X1 U421 ( .A(n499), .B(KEYINPUT19), .ZN(n628) );
  INV_X1 U422 ( .A(G119), .ZN(n444) );
  XNOR2_X1 U423 ( .A(n747), .B(n746), .ZN(n367) );
  NOR2_X1 U424 ( .A1(n757), .A2(n652), .ZN(n373) );
  NAND2_X1 U425 ( .A1(n429), .A2(n426), .ZN(n374) );
  NOR2_X1 U426 ( .A1(n641), .A2(n642), .ZN(n507) );
  NOR2_X1 U427 ( .A1(n659), .A2(n413), .ZN(n426) );
  BUF_X1 U428 ( .A(n779), .Z(n402) );
  AND2_X1 U429 ( .A1(n581), .A2(n427), .ZN(n659) );
  NOR2_X1 U430 ( .A1(n459), .A2(n699), .ZN(n612) );
  NAND2_X1 U431 ( .A1(n486), .A2(n485), .ZN(n480) );
  XNOR2_X1 U432 ( .A(n457), .B(KEYINPUT22), .ZN(n590) );
  AND2_X1 U433 ( .A1(n394), .A2(n395), .ZN(n635) );
  AND2_X1 U434 ( .A1(n380), .A2(n470), .ZN(n596) );
  INV_X1 U435 ( .A(n704), .ZN(n380) );
  NOR2_X1 U436 ( .A1(n386), .A2(KEYINPUT33), .ZN(n385) );
  AND2_X1 U437 ( .A1(n618), .A2(n407), .ZN(n452) );
  INV_X1 U438 ( .A(n386), .ZN(n365) );
  INV_X1 U439 ( .A(n592), .ZN(n366) );
  XNOR2_X1 U440 ( .A(n733), .B(n732), .ZN(n734) );
  XNOR2_X1 U441 ( .A(n544), .B(n435), .ZN(n546) );
  XNOR2_X1 U442 ( .A(n764), .B(n473), .ZN(n559) );
  INV_X1 U443 ( .A(n500), .ZN(n389) );
  XNOR2_X1 U444 ( .A(n541), .B(KEYINPUT10), .ZN(n575) );
  XNOR2_X1 U445 ( .A(KEYINPUT69), .B(G101), .ZN(n473) );
  XNOR2_X2 U446 ( .A(G128), .B(G110), .ZN(n571) );
  XNOR2_X2 U447 ( .A(KEYINPUT5), .B(KEYINPUT99), .ZN(n455) );
  NOR2_X1 U448 ( .A1(G953), .A2(G237), .ZN(n560) );
  NOR2_X1 U449 ( .A1(n367), .A2(n748), .ZN(G66) );
  NAND2_X1 U450 ( .A1(n738), .A2(G210), .ZN(n728) );
  XNOR2_X2 U451 ( .A(n503), .B(KEYINPUT65), .ZN(n738) );
  XNOR2_X1 U452 ( .A(n728), .B(n370), .ZN(n369) );
  INV_X1 U453 ( .A(n729), .ZN(n370) );
  XNOR2_X1 U454 ( .A(n657), .B(n372), .ZN(n371) );
  INV_X1 U455 ( .A(n417), .ZN(n372) );
  NAND2_X1 U456 ( .A1(n375), .A2(n373), .ZN(n440) );
  NAND2_X1 U457 ( .A1(n377), .A2(n376), .ZN(n375) );
  NAND2_X1 U458 ( .A1(n767), .A2(n441), .ZN(n376) );
  NAND2_X1 U459 ( .A1(n378), .A2(KEYINPUT76), .ZN(n377) );
  INV_X1 U460 ( .A(n767), .ZN(n378) );
  NAND2_X1 U461 ( .A1(n421), .A2(n379), .ZN(n422) );
  NAND2_X1 U462 ( .A1(n424), .A2(n379), .ZN(n423) );
  XNOR2_X1 U463 ( .A(n379), .B(G119), .ZN(G21) );
  XNOR2_X2 U464 ( .A(n502), .B(n389), .ZN(n379) );
  NAND2_X1 U465 ( .A1(n470), .A2(n390), .ZN(n457) );
  AND2_X1 U466 ( .A1(n470), .A2(n624), .ZN(n593) );
  XNOR2_X2 U467 ( .A(n391), .B(n361), .ZN(n470) );
  NAND2_X1 U468 ( .A1(n382), .A2(n381), .ZN(n387) );
  NAND2_X1 U469 ( .A1(n385), .A2(n384), .ZN(n381) );
  NAND2_X1 U470 ( .A1(n383), .A2(KEYINPUT33), .ZN(n382) );
  NAND2_X1 U471 ( .A1(n365), .A2(n384), .ZN(n587) );
  NOR2_X1 U472 ( .A1(n636), .A2(n592), .ZN(n594) );
  NAND2_X1 U473 ( .A1(n470), .A2(n387), .ZN(n469) );
  NAND2_X1 U474 ( .A1(n388), .A2(n494), .ZN(n493) );
  OR2_X1 U475 ( .A1(n388), .A2(n498), .ZN(n497) );
  XNOR2_X1 U476 ( .A(n388), .B(n727), .ZN(n729) );
  XNOR2_X2 U477 ( .A(n547), .B(n546), .ZN(n388) );
  NAND2_X1 U478 ( .A1(n628), .A2(n555), .ZN(n391) );
  XNOR2_X1 U479 ( .A(n506), .B(n505), .ZN(n479) );
  NAND2_X1 U480 ( .A1(n508), .A2(n507), .ZN(n506) );
  NAND2_X2 U481 ( .A1(n458), .A2(n497), .ZN(n433) );
  BUF_X1 U482 ( .A(n767), .Z(n392) );
  XNOR2_X1 U483 ( .A(n587), .B(KEYINPUT33), .ZN(n393) );
  NOR2_X1 U484 ( .A1(n610), .A2(n672), .ZN(n394) );
  AND2_X1 U485 ( .A1(n396), .A2(n645), .ZN(n395) );
  INV_X1 U486 ( .A(n644), .ZN(n396) );
  INV_X1 U487 ( .A(n624), .ZN(n397) );
  NOR2_X1 U488 ( .A1(n672), .A2(n610), .ZN(n611) );
  XNOR2_X1 U489 ( .A(n648), .B(n649), .ZN(n779) );
  BUF_X1 U490 ( .A(n749), .Z(n398) );
  BUF_X1 U491 ( .A(n656), .Z(n399) );
  BUF_X1 U492 ( .A(n646), .Z(n400) );
  BUF_X1 U493 ( .A(n688), .Z(n401) );
  XNOR2_X1 U494 ( .A(n400), .B(KEYINPUT41), .ZN(n403) );
  NOR2_X2 U495 ( .A1(n656), .A2(G902), .ZN(n567) );
  NOR2_X2 U496 ( .A1(n627), .A2(n592), .ZN(n616) );
  NAND2_X1 U497 ( .A1(n678), .A2(n640), .ZN(n641) );
  AND2_X1 U498 ( .A1(n777), .A2(n666), .ZN(n421) );
  INV_X1 U499 ( .A(n681), .ZN(n478) );
  XNOR2_X1 U500 ( .A(KEYINPUT15), .B(G902), .ZN(n652) );
  INV_X1 U501 ( .A(KEYINPUT46), .ZN(n509) );
  XOR2_X1 U502 ( .A(KEYINPUT95), .B(KEYINPUT81), .Z(n549) );
  AND2_X1 U503 ( .A1(n777), .A2(n405), .ZN(n424) );
  INV_X1 U504 ( .A(KEYINPUT8), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n765), .B(G146), .ZN(n565) );
  XNOR2_X1 U506 ( .A(n448), .B(KEYINPUT78), .ZN(n447) );
  INV_X1 U507 ( .A(KEYINPUT79), .ZN(n448) );
  INV_X1 U508 ( .A(KEYINPUT112), .ZN(n418) );
  XNOR2_X1 U509 ( .A(n533), .B(n528), .ZN(n460) );
  XNOR2_X1 U510 ( .A(n531), .B(n442), .ZN(n533) );
  XNOR2_X1 U511 ( .A(n464), .B(KEYINPUT77), .ZN(n504) );
  NOR2_X1 U512 ( .A1(n757), .A2(n491), .ZN(n464) );
  NAND2_X1 U513 ( .A1(n492), .A2(KEYINPUT2), .ZN(n491) );
  NOR2_X1 U514 ( .A1(n456), .A2(n414), .ZN(n485) );
  INV_X1 U515 ( .A(n463), .ZN(n644) );
  XNOR2_X1 U516 ( .A(n578), .B(n577), .ZN(n579) );
  INV_X1 U517 ( .A(KEYINPUT25), .ZN(n577) );
  NOR2_X1 U518 ( .A1(G902), .A2(n741), .ZN(n523) );
  NOR2_X1 U519 ( .A1(G952), .A2(n769), .ZN(n748) );
  INV_X1 U520 ( .A(n455), .ZN(n557) );
  INV_X1 U521 ( .A(KEYINPUT48), .ZN(n505) );
  OR2_X1 U522 ( .A1(G237), .A2(G902), .ZN(n551) );
  XOR2_X1 U523 ( .A(KEYINPUT97), .B(KEYINPUT21), .Z(n538) );
  INV_X1 U524 ( .A(n559), .ZN(n472) );
  XOR2_X1 U525 ( .A(KEYINPUT103), .B(KEYINPUT11), .Z(n530) );
  XNOR2_X1 U526 ( .A(n532), .B(n443), .ZN(n442) );
  INV_X1 U527 ( .A(KEYINPUT12), .ZN(n443) );
  XOR2_X1 U528 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n527) );
  XNOR2_X1 U529 ( .A(G113), .B(G122), .ZN(n526) );
  INV_X1 U530 ( .A(n575), .ZN(n568) );
  NAND2_X1 U531 ( .A1(n550), .A2(n496), .ZN(n495) );
  INV_X1 U532 ( .A(G472), .ZN(n471) );
  XOR2_X1 U533 ( .A(KEYINPUT7), .B(G122), .Z(n515) );
  XNOR2_X1 U534 ( .A(G116), .B(G107), .ZN(n514) );
  XOR2_X1 U535 ( .A(KEYINPUT9), .B(KEYINPUT104), .Z(n520) );
  XNOR2_X1 U536 ( .A(n542), .B(G134), .ZN(n517) );
  XNOR2_X1 U537 ( .A(n511), .B(n525), .ZN(n461) );
  XNOR2_X1 U538 ( .A(KEYINPUT16), .B(G122), .ZN(n540) );
  XNOR2_X1 U539 ( .A(n437), .B(n436), .ZN(n435) );
  XNOR2_X1 U540 ( .A(n406), .B(n543), .ZN(n437) );
  XNOR2_X1 U541 ( .A(n447), .B(n545), .ZN(n436) );
  NAND2_X1 U542 ( .A1(G234), .A2(G237), .ZN(n553) );
  NOR2_X1 U543 ( .A1(n484), .A2(n672), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n454), .B(n404), .ZN(n745) );
  XNOR2_X1 U545 ( .A(n574), .B(n575), .ZN(n454) );
  INV_X1 U546 ( .A(n504), .ZN(n720) );
  XNOR2_X1 U547 ( .A(n634), .B(KEYINPUT108), .ZN(n459) );
  NAND2_X1 U548 ( .A1(n411), .A2(n480), .ZN(n651) );
  NAND2_X1 U549 ( .A1(n450), .A2(n699), .ZN(n678) );
  INV_X1 U550 ( .A(KEYINPUT35), .ZN(n430) );
  XNOR2_X1 U551 ( .A(n501), .B(KEYINPUT32), .ZN(n500) );
  NAND2_X1 U552 ( .A1(n584), .A2(n583), .ZN(n502) );
  INV_X1 U553 ( .A(KEYINPUT80), .ZN(n501) );
  OR2_X2 U554 ( .A1(n597), .A2(n598), .ZN(n675) );
  XOR2_X1 U555 ( .A(n410), .B(n572), .Z(n404) );
  AND2_X1 U556 ( .A1(n666), .A2(KEYINPUT44), .ZN(n405) );
  INV_X1 U557 ( .A(n652), .ZN(n496) );
  XNOR2_X1 U558 ( .A(KEYINPUT17), .B(KEYINPUT93), .ZN(n406) );
  XOR2_X1 U559 ( .A(KEYINPUT82), .B(n606), .Z(n407) );
  XOR2_X1 U560 ( .A(KEYINPUT67), .B(KEYINPUT1), .Z(n408) );
  XOR2_X1 U561 ( .A(n571), .B(KEYINPUT24), .Z(n410) );
  AND2_X1 U562 ( .A1(n488), .A2(n487), .ZN(n411) );
  AND2_X1 U563 ( .A1(n585), .A2(n597), .ZN(n412) );
  AND2_X1 U564 ( .A1(n599), .A2(n687), .ZN(n413) );
  XOR2_X1 U565 ( .A(KEYINPUT72), .B(KEYINPUT39), .Z(n414) );
  XOR2_X1 U566 ( .A(KEYINPUT36), .B(KEYINPUT89), .Z(n415) );
  XNOR2_X1 U567 ( .A(KEYINPUT62), .B(n399), .ZN(n417) );
  INV_X1 U568 ( .A(KEYINPUT44), .ZN(n467) );
  INV_X1 U569 ( .A(KEYINPUT76), .ZN(n441) );
  NAND2_X1 U570 ( .A1(n420), .A2(n645), .ZN(n419) );
  XNOR2_X1 U571 ( .A(n433), .B(n643), .ZN(n420) );
  NAND2_X1 U572 ( .A1(n422), .A2(n467), .ZN(n425) );
  NAND2_X1 U573 ( .A1(n425), .A2(n423), .ZN(n429) );
  NOR2_X1 U574 ( .A1(n699), .A2(n428), .ZN(n427) );
  INV_X1 U575 ( .A(n363), .ZN(n428) );
  XNOR2_X1 U576 ( .A(n635), .B(n415), .ZN(n450) );
  NAND2_X1 U577 ( .A1(n468), .A2(n412), .ZN(n431) );
  XNOR2_X1 U578 ( .A(n449), .B(n509), .ZN(n508) );
  INV_X1 U579 ( .A(n655), .ZN(n492) );
  XNOR2_X1 U580 ( .A(n646), .B(KEYINPUT41), .ZN(n438) );
  XNOR2_X1 U581 ( .A(n469), .B(n588), .ZN(n468) );
  NAND2_X1 U582 ( .A1(n779), .A2(n781), .ZN(n449) );
  NAND2_X1 U583 ( .A1(n458), .A2(n497), .ZN(n432) );
  XNOR2_X1 U584 ( .A(n697), .B(KEYINPUT6), .ZN(n608) );
  AND2_X2 U585 ( .A1(n493), .A2(n495), .ZN(n458) );
  NAND2_X1 U586 ( .A1(n438), .A2(n647), .ZN(n648) );
  NAND2_X1 U587 ( .A1(n403), .A2(n393), .ZN(n716) );
  NAND2_X1 U588 ( .A1(n708), .A2(n403), .ZN(n709) );
  XNOR2_X2 U589 ( .A(n439), .B(n751), .ZN(n547) );
  XNOR2_X1 U590 ( .A(n439), .B(n461), .ZN(n476) );
  XNOR2_X2 U591 ( .A(n510), .B(n559), .ZN(n439) );
  NAND2_X1 U592 ( .A1(n440), .A2(n654), .ZN(n466) );
  XNOR2_X2 U593 ( .A(n534), .B(n535), .ZN(n597) );
  XNOR2_X1 U594 ( .A(n460), .B(n763), .ZN(n737) );
  XNOR2_X2 U595 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X2 U596 ( .A(KEYINPUT3), .B(KEYINPUT92), .ZN(n445) );
  XNOR2_X2 U597 ( .A(n749), .B(KEYINPUT71), .ZN(n510) );
  XNOR2_X2 U598 ( .A(n446), .B(n539), .ZN(n562) );
  XNOR2_X1 U599 ( .A(n614), .B(n615), .ZN(n618) );
  XNOR2_X2 U600 ( .A(n562), .B(n540), .ZN(n751) );
  NOR2_X1 U601 ( .A1(n608), .A2(n623), .ZN(n609) );
  INV_X4 U602 ( .A(G953), .ZN(n769) );
  XOR2_X2 U603 ( .A(n524), .B(G478), .Z(n598) );
  NAND2_X1 U604 ( .A1(n573), .A2(G217), .ZN(n519) );
  XNOR2_X2 U605 ( .A(n518), .B(n451), .ZN(n573) );
  XNOR2_X2 U606 ( .A(n489), .B(KEYINPUT40), .ZN(n781) );
  BUF_X1 U607 ( .A(n434), .Z(n456) );
  NOR2_X1 U608 ( .A1(n682), .A2(n478), .ZN(n477) );
  XNOR2_X1 U609 ( .A(n558), .B(n561), .ZN(n475) );
  XNOR2_X1 U610 ( .A(n475), .B(n472), .ZN(n564) );
  XOR2_X2 U611 ( .A(G146), .B(G125), .Z(n541) );
  NAND2_X1 U612 ( .A1(n650), .A2(n414), .ZN(n488) );
  XNOR2_X1 U613 ( .A(n739), .B(n416), .ZN(n462) );
  NOR2_X2 U614 ( .A1(n590), .A2(n586), .ZN(n584) );
  NAND2_X1 U615 ( .A1(n465), .A2(n504), .ZN(n503) );
  XNOR2_X1 U616 ( .A(n466), .B(KEYINPUT66), .ZN(n465) );
  XNOR2_X2 U617 ( .A(n567), .B(n471), .ZN(n697) );
  XNOR2_X2 U618 ( .A(n513), .B(n512), .ZN(n627) );
  XNOR2_X2 U619 ( .A(n474), .B(KEYINPUT64), .ZN(n764) );
  NOR2_X1 U620 ( .A1(n731), .A2(G902), .ZN(n513) );
  XNOR2_X1 U621 ( .A(n476), .B(n565), .ZN(n731) );
  INV_X1 U622 ( .A(n482), .ZN(n481) );
  NAND2_X1 U623 ( .A1(n488), .A2(n483), .ZN(n482) );
  INV_X1 U624 ( .A(n487), .ZN(n484) );
  INV_X1 U625 ( .A(n650), .ZN(n486) );
  NAND2_X1 U626 ( .A1(n434), .A2(n414), .ZN(n487) );
  XNOR2_X2 U627 ( .A(G143), .B(G128), .ZN(n542) );
  XNOR2_X1 U628 ( .A(n566), .B(n565), .ZN(n656) );
  XNOR2_X2 U629 ( .A(n490), .B(G107), .ZN(n749) );
  XNOR2_X2 U630 ( .A(G104), .B(G110), .ZN(n490) );
  NOR2_X1 U631 ( .A1(n550), .A2(n496), .ZN(n494) );
  INV_X1 U632 ( .A(n550), .ZN(n498) );
  NAND2_X1 U633 ( .A1(n432), .A2(n645), .ZN(n499) );
  XNOR2_X1 U634 ( .A(n735), .B(n734), .ZN(n736) );
  INV_X1 U635 ( .A(n562), .ZN(n563) );
  XNOR2_X1 U636 ( .A(n564), .B(n563), .ZN(n566) );
  AND2_X1 U637 ( .A1(n554), .A2(n604), .ZN(n555) );
  INV_X1 U638 ( .A(KEYINPUT38), .ZN(n643) );
  XNOR2_X1 U639 ( .A(n745), .B(n744), .ZN(n746) );
  OR2_X1 U640 ( .A1(n675), .A2(n651), .ZN(n681) );
  INV_X1 U641 ( .A(KEYINPUT63), .ZN(n658) );
  XNOR2_X1 U642 ( .A(n517), .B(G137), .ZN(n765) );
  AND2_X1 U643 ( .A1(G227), .A2(n769), .ZN(n511) );
  XNOR2_X1 U644 ( .A(KEYINPUT70), .B(G469), .ZN(n512) );
  INV_X1 U645 ( .A(n636), .ZN(n699) );
  XNOR2_X1 U646 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U647 ( .A(n517), .B(n516), .ZN(n522) );
  NAND2_X1 U648 ( .A1(G234), .A2(n769), .ZN(n518) );
  XNOR2_X1 U649 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U650 ( .A(n522), .B(n521), .ZN(n741) );
  XNOR2_X1 U651 ( .A(n523), .B(KEYINPUT105), .ZN(n524) );
  INV_X1 U652 ( .A(n598), .ZN(n585) );
  XNOR2_X1 U653 ( .A(KEYINPUT13), .B(G475), .ZN(n535) );
  XOR2_X1 U654 ( .A(n525), .B(n568), .Z(n763) );
  XNOR2_X1 U655 ( .A(n527), .B(n526), .ZN(n528) );
  NAND2_X1 U656 ( .A1(G214), .A2(n560), .ZN(n529) );
  XNOR2_X1 U657 ( .A(n530), .B(n529), .ZN(n531) );
  NOR2_X1 U658 ( .A1(G902), .A2(n737), .ZN(n534) );
  NAND2_X1 U659 ( .A1(n652), .A2(G234), .ZN(n536) );
  XNOR2_X1 U660 ( .A(n536), .B(KEYINPUT20), .ZN(n576) );
  NAND2_X1 U661 ( .A1(n576), .A2(G221), .ZN(n537) );
  XNOR2_X1 U662 ( .A(n538), .B(n537), .ZN(n694) );
  XNOR2_X1 U663 ( .A(G116), .B(G113), .ZN(n539) );
  XOR2_X1 U664 ( .A(n542), .B(n541), .Z(n544) );
  XNOR2_X1 U665 ( .A(KEYINPUT94), .B(KEYINPUT18), .ZN(n543) );
  NAND2_X1 U666 ( .A1(G224), .A2(n769), .ZN(n545) );
  NAND2_X1 U667 ( .A1(G210), .A2(n551), .ZN(n548) );
  XNOR2_X1 U668 ( .A(n549), .B(n548), .ZN(n550) );
  NAND2_X1 U669 ( .A1(G214), .A2(n551), .ZN(n645) );
  XNOR2_X1 U670 ( .A(G898), .B(KEYINPUT96), .ZN(n755) );
  NOR2_X1 U671 ( .A1(n769), .A2(n755), .ZN(n752) );
  NAND2_X1 U672 ( .A1(n752), .A2(G902), .ZN(n552) );
  NAND2_X1 U673 ( .A1(G952), .A2(n769), .ZN(n602) );
  NAND2_X1 U674 ( .A1(n552), .A2(n602), .ZN(n554) );
  XNOR2_X1 U675 ( .A(KEYINPUT14), .B(n553), .ZN(n604) );
  INV_X1 U676 ( .A(n604), .ZN(n713) );
  XNOR2_X1 U677 ( .A(n557), .B(n556), .ZN(n558) );
  NAND2_X1 U678 ( .A1(n560), .A2(G210), .ZN(n561) );
  XNOR2_X1 U679 ( .A(KEYINPUT88), .B(n584), .ZN(n581) );
  XOR2_X2 U680 ( .A(KEYINPUT23), .B(G140), .Z(n570) );
  XNOR2_X1 U681 ( .A(G119), .B(G137), .ZN(n569) );
  XNOR2_X1 U682 ( .A(n570), .B(n569), .ZN(n572) );
  NAND2_X1 U683 ( .A1(G221), .A2(n573), .ZN(n574) );
  NAND2_X1 U684 ( .A1(n576), .A2(G217), .ZN(n578) );
  NOR2_X1 U685 ( .A1(n636), .A2(n363), .ZN(n582) );
  XNOR2_X1 U686 ( .A(KEYINPUT106), .B(n582), .ZN(n583) );
  XNOR2_X1 U687 ( .A(KEYINPUT73), .B(KEYINPUT34), .ZN(n588) );
  INV_X1 U688 ( .A(n697), .ZN(n624) );
  NAND2_X1 U689 ( .A1(n693), .A2(n624), .ZN(n589) );
  NOR2_X1 U690 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U691 ( .A1(n591), .A2(n636), .ZN(n666) );
  NAND2_X1 U692 ( .A1(n616), .A2(n593), .ZN(n662) );
  NAND2_X1 U693 ( .A1(n397), .A2(n594), .ZN(n704) );
  XNOR2_X1 U694 ( .A(KEYINPUT100), .B(KEYINPUT31), .ZN(n595) );
  XNOR2_X1 U695 ( .A(n596), .B(n595), .ZN(n676) );
  NAND2_X1 U696 ( .A1(n662), .A2(n676), .ZN(n599) );
  NAND2_X1 U697 ( .A1(n672), .A2(n675), .ZN(n687) );
  XNOR2_X1 U698 ( .A(KEYINPUT87), .B(KEYINPUT45), .ZN(n600) );
  NOR2_X1 U699 ( .A1(n694), .A2(n363), .ZN(n607) );
  NOR2_X1 U700 ( .A1(G900), .A2(n769), .ZN(n601) );
  NAND2_X1 U701 ( .A1(n601), .A2(G902), .ZN(n603) );
  NAND2_X1 U702 ( .A1(n603), .A2(n602), .ZN(n605) );
  NAND2_X1 U703 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U704 ( .A1(n607), .A2(n407), .ZN(n623) );
  XNOR2_X1 U705 ( .A(n609), .B(KEYINPUT107), .ZN(n610) );
  NAND2_X1 U706 ( .A1(n611), .A2(n645), .ZN(n634) );
  XNOR2_X1 U707 ( .A(n612), .B(KEYINPUT43), .ZN(n613) );
  NOR2_X1 U708 ( .A1(n396), .A2(n613), .ZN(n682) );
  XOR2_X1 U709 ( .A(KEYINPUT110), .B(KEYINPUT30), .Z(n615) );
  NAND2_X1 U710 ( .A1(n697), .A2(n645), .ZN(n614) );
  NOR2_X1 U711 ( .A1(n644), .A2(n650), .ZN(n619) );
  INV_X1 U712 ( .A(KEYINPUT47), .ZN(n631) );
  AND2_X1 U713 ( .A1(n631), .A2(n687), .ZN(n621) );
  XNOR2_X1 U714 ( .A(n621), .B(KEYINPUT74), .ZN(n622) );
  NOR2_X1 U715 ( .A1(KEYINPUT85), .A2(n622), .ZN(n629) );
  XOR2_X1 U716 ( .A(KEYINPUT28), .B(n625), .Z(n626) );
  NOR2_X1 U717 ( .A1(n627), .A2(n626), .ZN(n647) );
  NAND2_X1 U718 ( .A1(n647), .A2(n628), .ZN(n670) );
  NOR2_X1 U719 ( .A1(n629), .A2(n670), .ZN(n630) );
  NOR2_X1 U720 ( .A1(n778), .A2(n630), .ZN(n633) );
  NAND2_X1 U721 ( .A1(KEYINPUT85), .A2(n631), .ZN(n632) );
  NAND2_X1 U722 ( .A1(n633), .A2(n632), .ZN(n642) );
  INV_X1 U723 ( .A(KEYINPUT85), .ZN(n637) );
  NAND2_X1 U724 ( .A1(n637), .A2(n670), .ZN(n638) );
  NAND2_X1 U725 ( .A1(n638), .A2(n687), .ZN(n639) );
  NAND2_X1 U726 ( .A1(n639), .A2(KEYINPUT47), .ZN(n640) );
  XOR2_X1 U727 ( .A(KEYINPUT113), .B(KEYINPUT42), .Z(n649) );
  INV_X1 U728 ( .A(n645), .ZN(n684) );
  NAND2_X1 U729 ( .A1(KEYINPUT2), .A2(n496), .ZN(n653) );
  NAND2_X1 U730 ( .A1(n738), .A2(G472), .ZN(n657) );
  XOR2_X1 U731 ( .A(G101), .B(n659), .Z(G3) );
  NOR2_X1 U732 ( .A1(n672), .A2(n662), .ZN(n660) );
  XOR2_X1 U733 ( .A(KEYINPUT114), .B(n660), .Z(n661) );
  XNOR2_X1 U734 ( .A(G104), .B(n661), .ZN(G6) );
  NOR2_X1 U735 ( .A1(n675), .A2(n662), .ZN(n664) );
  XNOR2_X1 U736 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n663) );
  XNOR2_X1 U737 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U738 ( .A(G107), .B(n665), .ZN(G9) );
  XNOR2_X1 U739 ( .A(G110), .B(n666), .ZN(G12) );
  NOR2_X1 U740 ( .A1(n675), .A2(n670), .ZN(n668) );
  XNOR2_X1 U741 ( .A(KEYINPUT29), .B(KEYINPUT115), .ZN(n667) );
  XNOR2_X1 U742 ( .A(n668), .B(n667), .ZN(n669) );
  XOR2_X1 U743 ( .A(G128), .B(n669), .Z(G30) );
  NOR2_X1 U744 ( .A1(n672), .A2(n670), .ZN(n671) );
  XOR2_X1 U745 ( .A(G146), .B(n671), .Z(G48) );
  NOR2_X1 U746 ( .A1(n676), .A2(n672), .ZN(n673) );
  XOR2_X1 U747 ( .A(KEYINPUT116), .B(n673), .Z(n674) );
  XNOR2_X1 U748 ( .A(G113), .B(n674), .ZN(G15) );
  NOR2_X1 U749 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U750 ( .A(G116), .B(n677), .Z(G18) );
  INV_X1 U751 ( .A(n678), .ZN(n679) );
  XNOR2_X1 U752 ( .A(G125), .B(n679), .ZN(n680) );
  XNOR2_X1 U753 ( .A(n680), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U754 ( .A(G134), .B(n681), .ZN(G36) );
  XNOR2_X1 U755 ( .A(G140), .B(n682), .ZN(n683) );
  XNOR2_X1 U756 ( .A(n683), .B(KEYINPUT117), .ZN(G42) );
  NAND2_X1 U757 ( .A1(n456), .A2(n684), .ZN(n686) );
  NAND2_X1 U758 ( .A1(n686), .A2(n685), .ZN(n690) );
  NAND2_X1 U759 ( .A1(n401), .A2(n687), .ZN(n689) );
  NAND2_X1 U760 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U761 ( .A(KEYINPUT121), .B(n691), .Z(n692) );
  NAND2_X1 U762 ( .A1(n692), .A2(n393), .ZN(n710) );
  NAND2_X1 U763 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U764 ( .A(KEYINPUT49), .B(n695), .ZN(n696) );
  NOR2_X1 U765 ( .A1(n397), .A2(n696), .ZN(n698) );
  XOR2_X1 U766 ( .A(KEYINPUT118), .B(n698), .Z(n702) );
  NOR2_X1 U767 ( .A1(n699), .A2(n366), .ZN(n700) );
  XNOR2_X1 U768 ( .A(KEYINPUT50), .B(n700), .ZN(n701) );
  NOR2_X1 U769 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U770 ( .A(n703), .B(KEYINPUT119), .ZN(n705) );
  NAND2_X1 U771 ( .A1(n705), .A2(n704), .ZN(n707) );
  XOR2_X1 U772 ( .A(KEYINPUT51), .B(KEYINPUT120), .Z(n706) );
  XNOR2_X1 U773 ( .A(n707), .B(n706), .ZN(n708) );
  NAND2_X1 U774 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U775 ( .A(KEYINPUT52), .B(n711), .Z(n712) );
  NOR2_X1 U776 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U777 ( .A1(n714), .A2(G952), .ZN(n715) );
  NAND2_X1 U778 ( .A1(n716), .A2(n715), .ZN(n722) );
  XNOR2_X1 U779 ( .A(KEYINPUT84), .B(KEYINPUT2), .ZN(n718) );
  NOR2_X1 U780 ( .A1(n757), .A2(n392), .ZN(n717) );
  NOR2_X1 U781 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U782 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U783 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U784 ( .A1(n769), .A2(n723), .ZN(n724) );
  XOR2_X1 U785 ( .A(KEYINPUT53), .B(n724), .Z(G75) );
  XOR2_X1 U786 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n726) );
  XNOR2_X1 U787 ( .A(KEYINPUT90), .B(KEYINPUT83), .ZN(n725) );
  XNOR2_X1 U788 ( .A(n726), .B(n725), .ZN(n727) );
  NAND2_X1 U789 ( .A1(n743), .A2(G469), .ZN(n735) );
  BUF_X1 U790 ( .A(n731), .Z(n733) );
  XOR2_X1 U791 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n732) );
  NOR2_X1 U792 ( .A1(n748), .A2(n736), .ZN(G54) );
  NAND2_X1 U793 ( .A1(n738), .A2(G475), .ZN(n739) );
  NAND2_X1 U794 ( .A1(n743), .A2(G478), .ZN(n740) );
  XNOR2_X1 U795 ( .A(n741), .B(n740), .ZN(n742) );
  NOR2_X1 U796 ( .A1(n742), .A2(n748), .ZN(G63) );
  NAND2_X1 U797 ( .A1(n743), .A2(G217), .ZN(n747) );
  XOR2_X1 U798 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n744) );
  XOR2_X1 U799 ( .A(n398), .B(G101), .Z(n750) );
  XNOR2_X1 U800 ( .A(n751), .B(n750), .ZN(n753) );
  NOR2_X1 U801 ( .A1(n753), .A2(n752), .ZN(n761) );
  NAND2_X1 U802 ( .A1(G953), .A2(G224), .ZN(n754) );
  XNOR2_X1 U803 ( .A(KEYINPUT61), .B(n754), .ZN(n756) );
  NAND2_X1 U804 ( .A1(n756), .A2(n755), .ZN(n759) );
  OR2_X1 U805 ( .A1(n757), .A2(G953), .ZN(n758) );
  NAND2_X1 U806 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U807 ( .A(n761), .B(n760), .ZN(n762) );
  XNOR2_X1 U808 ( .A(KEYINPUT124), .B(n762), .ZN(G69) );
  XNOR2_X1 U809 ( .A(n764), .B(n763), .ZN(n766) );
  XNOR2_X1 U810 ( .A(n766), .B(n765), .ZN(n771) );
  XOR2_X1 U811 ( .A(n392), .B(KEYINPUT125), .Z(n768) );
  XNOR2_X1 U812 ( .A(n771), .B(n768), .ZN(n770) );
  NAND2_X1 U813 ( .A1(n770), .A2(n769), .ZN(n775) );
  XNOR2_X1 U814 ( .A(G227), .B(n771), .ZN(n772) );
  NAND2_X1 U815 ( .A1(n772), .A2(G900), .ZN(n773) );
  NAND2_X1 U816 ( .A1(n773), .A2(G953), .ZN(n774) );
  NAND2_X1 U817 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U818 ( .A(KEYINPUT126), .B(n776), .ZN(G72) );
  XNOR2_X1 U819 ( .A(n777), .B(G122), .ZN(G24) );
  XOR2_X1 U820 ( .A(n778), .B(G143), .Z(G45) );
  XOR2_X1 U821 ( .A(n402), .B(G137), .Z(n780) );
  XNOR2_X1 U822 ( .A(KEYINPUT127), .B(n780), .ZN(G39) );
  XNOR2_X1 U823 ( .A(n781), .B(G131), .ZN(G33) );
endmodule

