

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577;

  AND2_X1 U321 ( .A1(G230GAT), .A2(G233GAT), .ZN(n289) );
  XNOR2_X1 U322 ( .A(KEYINPUT113), .B(KEYINPUT46), .ZN(n394) );
  XNOR2_X1 U323 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U324 ( .A(n362), .B(n289), .ZN(n364) );
  XNOR2_X1 U325 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U326 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U327 ( .A(n376), .B(n375), .ZN(n401) );
  XOR2_X1 U328 ( .A(KEYINPUT92), .B(n451), .Z(n504) );
  XNOR2_X1 U329 ( .A(n443), .B(G190GAT), .ZN(n444) );
  XNOR2_X1 U330 ( .A(n445), .B(n444), .ZN(G1351GAT) );
  XNOR2_X1 U331 ( .A(G36GAT), .B(G190GAT), .ZN(n290) );
  XNOR2_X1 U332 ( .A(n290), .B(KEYINPUT79), .ZN(n342) );
  XOR2_X1 U333 ( .A(KEYINPUT74), .B(G92GAT), .Z(n292) );
  XNOR2_X1 U334 ( .A(G99GAT), .B(G85GAT), .ZN(n291) );
  XNOR2_X1 U335 ( .A(n292), .B(n291), .ZN(n370) );
  XNOR2_X1 U336 ( .A(n342), .B(n370), .ZN(n310) );
  XOR2_X1 U337 ( .A(KEYINPUT78), .B(KEYINPUT11), .Z(n294) );
  XNOR2_X1 U338 ( .A(G218GAT), .B(KEYINPUT66), .ZN(n293) );
  XNOR2_X1 U339 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U340 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n296) );
  XNOR2_X1 U341 ( .A(KEYINPUT76), .B(KEYINPUT10), .ZN(n295) );
  XNOR2_X1 U342 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U343 ( .A(n298), .B(n297), .Z(n308) );
  XOR2_X1 U344 ( .A(KEYINPUT64), .B(KEYINPUT77), .Z(n300) );
  XNOR2_X1 U345 ( .A(G162GAT), .B(G106GAT), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n306) );
  XOR2_X1 U347 ( .A(G29GAT), .B(G134GAT), .Z(n311) );
  XOR2_X1 U348 ( .A(G43GAT), .B(G50GAT), .Z(n302) );
  XNOR2_X1 U349 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n380) );
  XOR2_X1 U351 ( .A(n311), .B(n380), .Z(n304) );
  NAND2_X1 U352 ( .A1(G232GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U353 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U354 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U355 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U356 ( .A(n310), .B(n309), .Z(n543) );
  INV_X1 U357 ( .A(n543), .ZN(n460) );
  XOR2_X1 U358 ( .A(KEYINPUT4), .B(KEYINPUT91), .Z(n313) );
  XOR2_X1 U359 ( .A(G120GAT), .B(G148GAT), .Z(n362) );
  XNOR2_X1 U360 ( .A(n311), .B(n362), .ZN(n312) );
  XNOR2_X1 U361 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U362 ( .A(n314), .B(KEYINPUT1), .Z(n320) );
  XNOR2_X1 U363 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n315) );
  XNOR2_X1 U364 ( .A(n315), .B(KEYINPUT83), .ZN(n433) );
  XOR2_X1 U365 ( .A(n433), .B(G57GAT), .Z(n317) );
  NAND2_X1 U366 ( .A1(G225GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U367 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n318), .B(G85GAT), .ZN(n319) );
  XNOR2_X1 U369 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U370 ( .A(KEYINPUT89), .B(KEYINPUT5), .Z(n322) );
  XNOR2_X1 U371 ( .A(KEYINPUT6), .B(KEYINPUT90), .ZN(n321) );
  XNOR2_X1 U372 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U373 ( .A(n324), .B(n323), .Z(n329) );
  XOR2_X1 U374 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n326) );
  XNOR2_X1 U375 ( .A(G141GAT), .B(G162GAT), .ZN(n325) );
  XNOR2_X1 U376 ( .A(n326), .B(n325), .ZN(n413) );
  XNOR2_X1 U377 ( .A(G1GAT), .B(G127GAT), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n327), .B(G155GAT), .ZN(n359) );
  XNOR2_X1 U379 ( .A(n413), .B(n359), .ZN(n328) );
  XNOR2_X1 U380 ( .A(n329), .B(n328), .ZN(n451) );
  XOR2_X1 U381 ( .A(KEYINPUT21), .B(G218GAT), .Z(n331) );
  XNOR2_X1 U382 ( .A(KEYINPUT88), .B(KEYINPUT87), .ZN(n330) );
  XNOR2_X1 U383 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U384 ( .A(G197GAT), .B(n332), .Z(n423) );
  XNOR2_X1 U385 ( .A(G8GAT), .B(G183GAT), .ZN(n333) );
  XNOR2_X1 U386 ( .A(n333), .B(G211GAT), .ZN(n358) );
  XOR2_X1 U387 ( .A(G176GAT), .B(G64GAT), .Z(n366) );
  XOR2_X1 U388 ( .A(n358), .B(n366), .Z(n335) );
  XNOR2_X1 U389 ( .A(G204GAT), .B(G92GAT), .ZN(n334) );
  XNOR2_X1 U390 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U391 ( .A(n423), .B(n336), .ZN(n346) );
  XOR2_X1 U392 ( .A(KEYINPUT95), .B(KEYINPUT93), .Z(n338) );
  NAND2_X1 U393 ( .A1(G226GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U395 ( .A(n339), .B(KEYINPUT94), .Z(n344) );
  XOR2_X1 U396 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n341) );
  XNOR2_X1 U397 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n341), .B(n340), .ZN(n434) );
  XNOR2_X1 U399 ( .A(n434), .B(n342), .ZN(n343) );
  XNOR2_X1 U400 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U401 ( .A(n346), .B(n345), .Z(n508) );
  INV_X1 U402 ( .A(n508), .ZN(n407) );
  XOR2_X1 U403 ( .A(KEYINPUT12), .B(KEYINPUT80), .Z(n348) );
  NAND2_X1 U404 ( .A1(G231GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U405 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U406 ( .A(n349), .B(KEYINPUT81), .Z(n353) );
  XNOR2_X1 U407 ( .A(G15GAT), .B(G22GAT), .ZN(n350) );
  XNOR2_X1 U408 ( .A(n350), .B(KEYINPUT70), .ZN(n378) );
  XNOR2_X1 U409 ( .A(G71GAT), .B(G57GAT), .ZN(n351) );
  XNOR2_X1 U410 ( .A(n351), .B(KEYINPUT13), .ZN(n363) );
  XNOR2_X1 U411 ( .A(n378), .B(n363), .ZN(n352) );
  XNOR2_X1 U412 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U413 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n355) );
  XNOR2_X1 U414 ( .A(G78GAT), .B(G64GAT), .ZN(n354) );
  XNOR2_X1 U415 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U416 ( .A(n357), .B(n356), .Z(n361) );
  XNOR2_X1 U417 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U418 ( .A(n361), .B(n360), .Z(n572) );
  XOR2_X1 U419 ( .A(n572), .B(KEYINPUT112), .Z(n559) );
  XOR2_X1 U420 ( .A(n365), .B(KEYINPUT75), .Z(n368) );
  XNOR2_X1 U421 ( .A(n366), .B(KEYINPUT72), .ZN(n367) );
  XNOR2_X1 U422 ( .A(n368), .B(n367), .ZN(n376) );
  XNOR2_X1 U423 ( .A(G106GAT), .B(G78GAT), .ZN(n369) );
  XNOR2_X1 U424 ( .A(n369), .B(G204GAT), .ZN(n410) );
  XOR2_X1 U425 ( .A(n410), .B(n370), .Z(n374) );
  XOR2_X1 U426 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n372) );
  XNOR2_X1 U427 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n371) );
  XNOR2_X1 U428 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U429 ( .A(n401), .B(KEYINPUT41), .ZN(n551) );
  XNOR2_X1 U430 ( .A(G113GAT), .B(G29GAT), .ZN(n377) );
  XNOR2_X1 U431 ( .A(n377), .B(G36GAT), .ZN(n379) );
  XOR2_X1 U432 ( .A(n379), .B(n378), .Z(n385) );
  XOR2_X1 U433 ( .A(n380), .B(KEYINPUT30), .Z(n382) );
  NAND2_X1 U434 ( .A1(G229GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U435 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U436 ( .A(G169GAT), .B(n383), .ZN(n384) );
  XNOR2_X1 U437 ( .A(n385), .B(n384), .ZN(n393) );
  XOR2_X1 U438 ( .A(G8GAT), .B(G1GAT), .Z(n387) );
  XNOR2_X1 U439 ( .A(G141GAT), .B(G197GAT), .ZN(n386) );
  XNOR2_X1 U440 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U441 ( .A(KEYINPUT69), .B(KEYINPUT29), .Z(n389) );
  XNOR2_X1 U442 ( .A(KEYINPUT71), .B(KEYINPUT68), .ZN(n388) );
  XNOR2_X1 U443 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U444 ( .A(n391), .B(n390), .Z(n392) );
  XOR2_X1 U445 ( .A(n393), .B(n392), .Z(n534) );
  NAND2_X1 U446 ( .A1(n551), .A2(n534), .ZN(n395) );
  NOR2_X1 U447 ( .A1(n559), .A2(n396), .ZN(n397) );
  XNOR2_X1 U448 ( .A(n397), .B(KEYINPUT114), .ZN(n398) );
  NAND2_X1 U449 ( .A1(n398), .A2(n460), .ZN(n399) );
  XNOR2_X1 U450 ( .A(n399), .B(KEYINPUT47), .ZN(n405) );
  XOR2_X1 U451 ( .A(KEYINPUT36), .B(n543), .Z(n575) );
  NOR2_X1 U452 ( .A1(n575), .A2(n572), .ZN(n400) );
  XNOR2_X1 U453 ( .A(KEYINPUT45), .B(n400), .ZN(n402) );
  NAND2_X1 U454 ( .A1(n402), .A2(n401), .ZN(n403) );
  NOR2_X1 U455 ( .A1(n403), .A2(n534), .ZN(n404) );
  NOR2_X1 U456 ( .A1(n405), .A2(n404), .ZN(n406) );
  XNOR2_X1 U457 ( .A(n406), .B(KEYINPUT48), .ZN(n517) );
  NOR2_X1 U458 ( .A1(n407), .A2(n517), .ZN(n408) );
  XOR2_X1 U459 ( .A(KEYINPUT54), .B(n408), .Z(n409) );
  NOR2_X1 U460 ( .A1(n504), .A2(n409), .ZN(n565) );
  XOR2_X1 U461 ( .A(G155GAT), .B(n410), .Z(n412) );
  NAND2_X1 U462 ( .A1(G228GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U463 ( .A(n412), .B(n411), .ZN(n416) );
  XNOR2_X1 U464 ( .A(G22GAT), .B(n413), .ZN(n414) );
  XNOR2_X1 U465 ( .A(n414), .B(G211GAT), .ZN(n415) );
  XOR2_X1 U466 ( .A(n416), .B(n415), .Z(n421) );
  XOR2_X1 U467 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n418) );
  XNOR2_X1 U468 ( .A(G148GAT), .B(KEYINPUT24), .ZN(n417) );
  XNOR2_X1 U469 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U470 ( .A(G50GAT), .B(n419), .ZN(n420) );
  XNOR2_X1 U471 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U472 ( .A(n423), .B(n422), .ZN(n454) );
  NAND2_X1 U473 ( .A1(n565), .A2(n454), .ZN(n424) );
  XNOR2_X1 U474 ( .A(n424), .B(KEYINPUT55), .ZN(n557) );
  XOR2_X1 U475 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n426) );
  XNOR2_X1 U476 ( .A(G120GAT), .B(G183GAT), .ZN(n425) );
  XNOR2_X1 U477 ( .A(n426), .B(n425), .ZN(n442) );
  XOR2_X1 U478 ( .A(G127GAT), .B(G190GAT), .Z(n428) );
  XNOR2_X1 U479 ( .A(G43GAT), .B(G15GAT), .ZN(n427) );
  XNOR2_X1 U480 ( .A(n428), .B(n427), .ZN(n430) );
  XOR2_X1 U481 ( .A(G134GAT), .B(G99GAT), .Z(n429) );
  XNOR2_X1 U482 ( .A(n430), .B(n429), .ZN(n438) );
  XNOR2_X1 U483 ( .A(KEYINPUT86), .B(G176GAT), .ZN(n431) );
  XNOR2_X1 U484 ( .A(n431), .B(G71GAT), .ZN(n432) );
  XOR2_X1 U485 ( .A(n432), .B(KEYINPUT20), .Z(n436) );
  XNOR2_X1 U486 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U487 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U488 ( .A(n438), .B(n437), .ZN(n440) );
  NAND2_X1 U489 ( .A1(G227GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U490 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U491 ( .A(n442), .B(n441), .Z(n456) );
  INV_X1 U492 ( .A(n456), .ZN(n556) );
  NAND2_X1 U493 ( .A1(n557), .A2(n556), .ZN(n548) );
  NOR2_X1 U494 ( .A1(n460), .A2(n548), .ZN(n445) );
  XNOR2_X1 U495 ( .A(KEYINPUT58), .B(KEYINPUT125), .ZN(n443) );
  XOR2_X1 U496 ( .A(KEYINPUT34), .B(KEYINPUT98), .Z(n466) );
  NAND2_X1 U497 ( .A1(n534), .A2(n401), .ZN(n477) );
  XNOR2_X1 U498 ( .A(n508), .B(KEYINPUT27), .ZN(n453) );
  NOR2_X1 U499 ( .A1(n454), .A2(n556), .ZN(n446) );
  XNOR2_X1 U500 ( .A(n446), .B(KEYINPUT26), .ZN(n564) );
  NAND2_X1 U501 ( .A1(n453), .A2(n564), .ZN(n450) );
  NAND2_X1 U502 ( .A1(n556), .A2(n508), .ZN(n447) );
  NAND2_X1 U503 ( .A1(n454), .A2(n447), .ZN(n448) );
  XOR2_X1 U504 ( .A(KEYINPUT25), .B(n448), .Z(n449) );
  NAND2_X1 U505 ( .A1(n450), .A2(n449), .ZN(n452) );
  NAND2_X1 U506 ( .A1(n452), .A2(n451), .ZN(n459) );
  NAND2_X1 U507 ( .A1(n504), .A2(n453), .ZN(n531) );
  XNOR2_X1 U508 ( .A(KEYINPUT67), .B(KEYINPUT28), .ZN(n455) );
  XNOR2_X1 U509 ( .A(n455), .B(n454), .ZN(n512) );
  NOR2_X1 U510 ( .A1(n531), .A2(n512), .ZN(n518) );
  NAND2_X1 U511 ( .A1(n456), .A2(n518), .ZN(n457) );
  XNOR2_X1 U512 ( .A(KEYINPUT96), .B(n457), .ZN(n458) );
  NAND2_X1 U513 ( .A1(n459), .A2(n458), .ZN(n475) );
  XOR2_X1 U514 ( .A(KEYINPUT16), .B(KEYINPUT82), .Z(n462) );
  INV_X1 U515 ( .A(n572), .ZN(n541) );
  NAND2_X1 U516 ( .A1(n541), .A2(n460), .ZN(n461) );
  XNOR2_X1 U517 ( .A(n462), .B(n461), .ZN(n463) );
  NAND2_X1 U518 ( .A1(n475), .A2(n463), .ZN(n464) );
  XOR2_X1 U519 ( .A(KEYINPUT97), .B(n464), .Z(n491) );
  NOR2_X1 U520 ( .A1(n477), .A2(n491), .ZN(n472) );
  NAND2_X1 U521 ( .A1(n472), .A2(n504), .ZN(n465) );
  XNOR2_X1 U522 ( .A(n466), .B(n465), .ZN(n467) );
  XOR2_X1 U523 ( .A(G1GAT), .B(n467), .Z(G1324GAT) );
  XOR2_X1 U524 ( .A(G8GAT), .B(KEYINPUT99), .Z(n469) );
  NAND2_X1 U525 ( .A1(n472), .A2(n508), .ZN(n468) );
  XNOR2_X1 U526 ( .A(n469), .B(n468), .ZN(G1325GAT) );
  XOR2_X1 U527 ( .A(G15GAT), .B(KEYINPUT35), .Z(n471) );
  NAND2_X1 U528 ( .A1(n472), .A2(n556), .ZN(n470) );
  XNOR2_X1 U529 ( .A(n471), .B(n470), .ZN(G1326GAT) );
  NAND2_X1 U530 ( .A1(n512), .A2(n472), .ZN(n473) );
  XNOR2_X1 U531 ( .A(n473), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U532 ( .A1(n541), .A2(n575), .ZN(n474) );
  NAND2_X1 U533 ( .A1(n475), .A2(n474), .ZN(n476) );
  XOR2_X1 U534 ( .A(KEYINPUT37), .B(n476), .Z(n502) );
  NOR2_X1 U535 ( .A1(n502), .A2(n477), .ZN(n479) );
  XNOR2_X1 U536 ( .A(KEYINPUT100), .B(KEYINPUT38), .ZN(n478) );
  XNOR2_X1 U537 ( .A(n479), .B(n478), .ZN(n487) );
  NAND2_X1 U538 ( .A1(n487), .A2(n504), .ZN(n482) );
  XNOR2_X1 U539 ( .A(G29GAT), .B(KEYINPUT101), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n480), .B(KEYINPUT39), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n482), .B(n481), .ZN(G1328GAT) );
  NAND2_X1 U542 ( .A1(n508), .A2(n487), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n483), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U544 ( .A(KEYINPUT40), .B(KEYINPUT102), .Z(n485) );
  NAND2_X1 U545 ( .A1(n487), .A2(n556), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U547 ( .A(G43GAT), .B(n486), .Z(G1330GAT) );
  XOR2_X1 U548 ( .A(G50GAT), .B(KEYINPUT103), .Z(n489) );
  NAND2_X1 U549 ( .A1(n487), .A2(n512), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n489), .B(n488), .ZN(G1331GAT) );
  INV_X1 U551 ( .A(n534), .ZN(n566) );
  NAND2_X1 U552 ( .A1(n551), .A2(n566), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n490), .B(KEYINPUT104), .ZN(n503) );
  NOR2_X1 U554 ( .A1(n503), .A2(n491), .ZN(n498) );
  NAND2_X1 U555 ( .A1(n498), .A2(n504), .ZN(n495) );
  XOR2_X1 U556 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n493) );
  XNOR2_X1 U557 ( .A(G57GAT), .B(KEYINPUT106), .ZN(n492) );
  XNOR2_X1 U558 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U559 ( .A(n495), .B(n494), .ZN(G1332GAT) );
  NAND2_X1 U560 ( .A1(n508), .A2(n498), .ZN(n496) );
  XNOR2_X1 U561 ( .A(n496), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U562 ( .A1(n556), .A2(n498), .ZN(n497) );
  XNOR2_X1 U563 ( .A(n497), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n500) );
  NAND2_X1 U565 ( .A1(n498), .A2(n512), .ZN(n499) );
  XNOR2_X1 U566 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U567 ( .A(G78GAT), .B(n501), .Z(G1335GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n506) );
  NOR2_X1 U569 ( .A1(n503), .A2(n502), .ZN(n513) );
  NAND2_X1 U570 ( .A1(n513), .A2(n504), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U572 ( .A(G85GAT), .B(n507), .ZN(G1336GAT) );
  NAND2_X1 U573 ( .A1(n508), .A2(n513), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n509), .B(KEYINPUT110), .ZN(n510) );
  XNOR2_X1 U575 ( .A(G92GAT), .B(n510), .ZN(G1337GAT) );
  NAND2_X1 U576 ( .A1(n556), .A2(n513), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n511), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT111), .B(KEYINPUT44), .Z(n515) );
  NAND2_X1 U579 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U581 ( .A(G106GAT), .B(n516), .ZN(G1339GAT) );
  NAND2_X1 U582 ( .A1(n518), .A2(n556), .ZN(n519) );
  NOR2_X1 U583 ( .A1(n517), .A2(n519), .ZN(n528) );
  NAND2_X1 U584 ( .A1(n528), .A2(n534), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n520), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT117), .B(KEYINPUT116), .Z(n522) );
  XNOR2_X1 U587 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n522), .B(n521), .ZN(n525) );
  NAND2_X1 U589 ( .A1(n551), .A2(n528), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n523), .B(KEYINPUT115), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(G1341GAT) );
  NAND2_X1 U592 ( .A1(n559), .A2(n528), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n526), .B(KEYINPUT50), .ZN(n527) );
  XNOR2_X1 U594 ( .A(G127GAT), .B(n527), .ZN(G1342GAT) );
  XOR2_X1 U595 ( .A(G134GAT), .B(KEYINPUT51), .Z(n530) );
  NAND2_X1 U596 ( .A1(n528), .A2(n543), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n530), .B(n529), .ZN(G1343GAT) );
  XOR2_X1 U598 ( .A(G141GAT), .B(KEYINPUT119), .Z(n536) );
  NOR2_X1 U599 ( .A1(n517), .A2(n531), .ZN(n532) );
  NAND2_X1 U600 ( .A1(n564), .A2(n532), .ZN(n533) );
  XOR2_X1 U601 ( .A(KEYINPUT118), .B(n533), .Z(n544) );
  NAND2_X1 U602 ( .A1(n534), .A2(n544), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(G1344GAT) );
  XNOR2_X1 U604 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n540) );
  XOR2_X1 U605 ( .A(KEYINPUT120), .B(KEYINPUT52), .Z(n538) );
  NAND2_X1 U606 ( .A1(n544), .A2(n551), .ZN(n537) );
  XNOR2_X1 U607 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U608 ( .A(n540), .B(n539), .ZN(G1345GAT) );
  NAND2_X1 U609 ( .A1(n544), .A2(n541), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n542), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n546) );
  NAND2_X1 U612 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(G162GAT), .B(n547), .ZN(G1347GAT) );
  NOR2_X1 U615 ( .A1(n566), .A2(n548), .ZN(n550) );
  XNOR2_X1 U616 ( .A(G169GAT), .B(KEYINPUT123), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(G1348GAT) );
  AND2_X1 U618 ( .A1(n551), .A2(n556), .ZN(n552) );
  AND2_X1 U619 ( .A1(n557), .A2(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(G176GAT), .B(n555), .ZN(G1349GAT) );
  AND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n560), .B(KEYINPUT124), .ZN(n561) );
  XNOR2_X1 U626 ( .A(G183GAT), .B(n561), .ZN(G1350GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT59), .B(KEYINPUT126), .Z(n563) );
  XNOR2_X1 U628 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n568) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n574) );
  NOR2_X1 U631 ( .A1(n566), .A2(n574), .ZN(n567) );
  XOR2_X1 U632 ( .A(n568), .B(n567), .Z(G1352GAT) );
  NOR2_X1 U633 ( .A1(n401), .A2(n574), .ZN(n570) );
  XNOR2_X1 U634 ( .A(KEYINPUT61), .B(KEYINPUT127), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XOR2_X1 U636 ( .A(G204GAT), .B(n571), .Z(G1353GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n574), .ZN(n573) );
  XOR2_X1 U638 ( .A(G211GAT), .B(n573), .Z(G1354GAT) );
  NOR2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U640 ( .A(KEYINPUT62), .B(n576), .Z(n577) );
  XNOR2_X1 U641 ( .A(G218GAT), .B(n577), .ZN(G1355GAT) );
endmodule

