//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 0 1 1 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n566, new_n568, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1173, new_n1174;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT67), .Z(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(new_n466), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n473), .A2(KEYINPUT3), .A3(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n475), .A2(G137), .A3(new_n476), .A4(new_n465), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n473), .A2(new_n474), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n478), .A2(G101), .A3(new_n476), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n471), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT69), .ZN(G160));
  NAND2_X1  g056(.A1(new_n475), .A2(new_n465), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT70), .Z(new_n485));
  NOR2_X1   g060(.A1(new_n482), .A2(new_n476), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  INV_X1    g062(.A(G100), .ZN(new_n488));
  AND3_X1   g063(.A1(new_n488), .A2(new_n476), .A3(KEYINPUT71), .ZN(new_n489));
  AOI21_X1  g064(.A(KEYINPUT71), .B1(new_n488), .B2(new_n476), .ZN(new_n490));
  OAI221_X1 g065(.A(G2104), .B1(G112), .B2(new_n476), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n485), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  XOR2_X1   g067(.A(new_n492), .B(KEYINPUT72), .Z(G162));
  AND2_X1   g068(.A1(KEYINPUT4), .A2(G138), .ZN(new_n494));
  AND3_X1   g069(.A1(new_n475), .A2(new_n465), .A3(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(G102), .A2(G2104), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n476), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n475), .A2(G126), .A3(new_n465), .ZN(new_n498));
  NAND2_X1  g073(.A1(G114), .A2(G2104), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n465), .A2(new_n467), .A3(G138), .A4(new_n476), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n497), .A2(new_n501), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n504), .B1(new_n500), .B2(G2105), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(KEYINPUT73), .A3(new_n497), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  AND3_X1   g091(.A1(new_n516), .A2(KEYINPUT74), .A3(KEYINPUT5), .ZN(new_n517));
  AOI21_X1  g092(.A(KEYINPUT74), .B1(new_n516), .B2(KEYINPUT5), .ZN(new_n518));
  OAI211_X1 g093(.A(new_n513), .B(new_n515), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT75), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n521), .B1(new_n514), .B2(G543), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n516), .A2(KEYINPUT74), .A3(KEYINPUT5), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n522), .A2(new_n523), .B1(new_n514), .B2(G543), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT75), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n524), .A2(new_n525), .A3(new_n513), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  XOR2_X1   g102(.A(KEYINPUT76), .B(G88), .Z(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(G75), .A2(G543), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n531));
  INV_X1    g106(.A(G62), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n513), .A2(G543), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n533), .A2(G651), .B1(G50), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n529), .A2(new_n535), .ZN(G303));
  INV_X1    g111(.A(G303), .ZN(G166));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n520), .A2(new_n526), .ZN(new_n540));
  INV_X1    g115(.A(G89), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT78), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n543), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n524), .A2(G63), .A3(G651), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(KEYINPUT77), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(KEYINPUT77), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n547), .A2(new_n548), .B1(G51), .B2(new_n534), .ZN(new_n549));
  AND3_X1   g124(.A1(new_n544), .A2(new_n545), .A3(new_n549), .ZN(G168));
  NAND2_X1  g125(.A1(new_n527), .A2(G90), .ZN(new_n551));
  NAND2_X1  g126(.A1(G77), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G64), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n531), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n554), .A2(G651), .B1(G52), .B2(new_n534), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n551), .A2(new_n555), .ZN(G301));
  INV_X1    g131(.A(G301), .ZN(G171));
  NAND2_X1  g132(.A1(G68), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G56), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n531), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G651), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT79), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n527), .A2(G81), .B1(G43), .B2(new_n534), .ZN(new_n563));
  AND2_X1   g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  AND3_X1   g140(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G36), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT80), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(G188));
  NAND2_X1  g146(.A1(new_n534), .A2(G53), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT9), .ZN(new_n573));
  INV_X1    g148(.A(G91), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n574), .B2(new_n540), .ZN(new_n575));
  INV_X1    g150(.A(G651), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n531), .B(KEYINPUT81), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G65), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n576), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G299));
  NAND3_X1  g157(.A1(new_n544), .A2(new_n545), .A3(new_n549), .ZN(G286));
  INV_X1    g158(.A(G74), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n531), .A2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(new_n534), .B2(G49), .ZN(new_n586));
  INV_X1    g161(.A(G87), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n540), .B2(new_n587), .ZN(G288));
  INV_X1    g163(.A(KEYINPUT82), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n524), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n590), .B2(new_n576), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n520), .A2(G86), .A3(new_n526), .ZN(new_n592));
  OAI211_X1 g167(.A(G61), .B(new_n515), .C1(new_n517), .C2(new_n518), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n595), .A2(KEYINPUT82), .A3(G651), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n534), .A2(G48), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n591), .A2(new_n592), .A3(new_n596), .A4(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(new_n527), .A2(G85), .ZN(new_n599));
  NAND2_X1  g174(.A1(G72), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G60), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n531), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(G47), .B2(new_n534), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n599), .A2(new_n603), .ZN(G290));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NOR2_X1   g180(.A1(G301), .A2(new_n605), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n577), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT84), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n576), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(new_n608), .B2(new_n607), .ZN(new_n610));
  XOR2_X1   g185(.A(KEYINPUT83), .B(KEYINPUT10), .Z(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n540), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n534), .A2(G54), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR3_X1   g190(.A1(new_n540), .A2(new_n612), .A3(new_n611), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g192(.A1(new_n610), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n606), .B1(new_n618), .B2(new_n605), .ZN(G284));
  AOI21_X1  g194(.A(new_n606), .B1(new_n618), .B2(new_n605), .ZN(G321));
  MUX2_X1   g195(.A(G286), .B(G299), .S(new_n605), .Z(G297));
  MUX2_X1   g196(.A(G286), .B(G299), .S(new_n605), .Z(G280));
  XNOR2_X1  g197(.A(KEYINPUT85), .B(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n618), .B1(G860), .B2(new_n623), .ZN(G148));
  NAND2_X1  g199(.A1(new_n562), .A2(new_n563), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(new_n605), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n618), .A2(new_n623), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT86), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n626), .B1(new_n628), .B2(new_n605), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND4_X1  g205(.A1(new_n478), .A2(new_n476), .A3(new_n465), .A4(new_n467), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2100), .ZN(new_n634));
  MUX2_X1   g209(.A(G99), .B(G111), .S(G2105), .Z(new_n635));
  AOI22_X1  g210(.A1(new_n486), .A2(G123), .B1(G2104), .B2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(G135), .ZN(new_n637));
  INV_X1    g212(.A(new_n483), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(G2096), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n634), .A2(new_n641), .ZN(G156));
  INV_X1    g217(.A(KEYINPUT14), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT15), .B(G2435), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2427), .ZN(new_n646));
  INV_X1    g221(.A(G2430), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n643), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n647), .B2(new_n646), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n649), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n649), .A2(new_n655), .ZN(new_n657));
  AND3_X1   g232(.A1(new_n656), .A2(G14), .A3(new_n657), .ZN(G401));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2072), .B(G2078), .Z(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  NOR3_X1   g238(.A1(new_n660), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT18), .ZN(new_n665));
  INV_X1    g240(.A(new_n661), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(KEYINPUT17), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n662), .B1(new_n668), .B2(new_n659), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n669), .B1(new_n660), .B2(new_n667), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n660), .A2(new_n663), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n666), .B1(new_n671), .B2(KEYINPUT17), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n665), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(new_n640), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G2100), .ZN(G227));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT88), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G1971), .B(G1976), .Z(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT20), .Z(new_n684));
  NAND2_X1  g259(.A1(new_n677), .A2(new_n678), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n685), .A2(new_n682), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT89), .Z(new_n687));
  NAND3_X1  g262(.A1(new_n679), .A2(new_n682), .A3(new_n685), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n684), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n691), .B(new_n694), .ZN(G229));
  MUX2_X1   g270(.A(G23), .B(G288), .S(G16), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT92), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT33), .B(G1976), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT93), .Z(new_n699));
  XOR2_X1   g274(.A(new_n697), .B(new_n699), .Z(new_n700));
  NOR2_X1   g275(.A1(G6), .A2(G16), .ZN(new_n701));
  INV_X1    g276(.A(G305), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(G16), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT32), .B(G1981), .Z(new_n704));
  XOR2_X1   g279(.A(new_n703), .B(new_n704), .Z(new_n705));
  NOR2_X1   g280(.A1(G16), .A2(G22), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G166), .B2(G16), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1971), .ZN(new_n708));
  NOR3_X1   g283(.A1(new_n700), .A2(new_n705), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT34), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(new_n710), .ZN(new_n712));
  MUX2_X1   g287(.A(G24), .B(G290), .S(G16), .Z(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G1986), .ZN(new_n714));
  NOR2_X1   g289(.A1(G25), .A2(G29), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n483), .A2(G131), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n486), .A2(G119), .ZN(new_n717));
  INV_X1    g292(.A(G95), .ZN(new_n718));
  AND3_X1   g293(.A1(new_n718), .A2(new_n476), .A3(KEYINPUT90), .ZN(new_n719));
  AOI21_X1  g294(.A(KEYINPUT90), .B1(new_n718), .B2(new_n476), .ZN(new_n720));
  OAI221_X1 g295(.A(G2104), .B1(G107), .B2(new_n476), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n716), .A2(new_n717), .A3(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n715), .B1(new_n723), .B2(G29), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT35), .B(G1991), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT91), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n724), .B(new_n726), .Z(new_n727));
  NOR2_X1   g302(.A1(new_n713), .A2(G1986), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n711), .A2(new_n712), .A3(new_n714), .A4(new_n729), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT36), .Z(new_n731));
  NOR2_X1   g306(.A1(G4), .A2(G16), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n618), .B2(G16), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G1348), .ZN(new_n734));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G35), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G162), .B2(new_n735), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT29), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G2090), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n734), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(G5), .A2(G16), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G171), .B2(G16), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT100), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G1961), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT24), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n746), .A2(G34), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(G34), .ZN(new_n748));
  AOI21_X1  g323(.A(G29), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G160), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n749), .B1(new_n750), .B2(G29), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT97), .Z(new_n752));
  INV_X1    g327(.A(G2084), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n745), .A2(new_n754), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n741), .B(new_n755), .C1(new_n740), .C2(new_n739), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n483), .A2(G139), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT96), .B(KEYINPUT25), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n465), .A2(new_n467), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n763), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n764));
  OAI221_X1 g339(.A(new_n757), .B1(new_n761), .B2(new_n762), .C1(new_n476), .C2(new_n764), .ZN(new_n765));
  MUX2_X1   g340(.A(G33), .B(new_n765), .S(G29), .Z(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(G2072), .Z(new_n767));
  XOR2_X1   g342(.A(KEYINPUT31), .B(G11), .Z(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT30), .B(G28), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n768), .B1(new_n735), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n639), .B2(new_n735), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n735), .A2(G32), .ZN(new_n772));
  NAND3_X1  g347(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT98), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(KEYINPUT26), .ZN(new_n775));
  AOI22_X1  g350(.A1(G129), .A2(new_n486), .B1(new_n483), .B2(G141), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n774), .A2(KEYINPUT26), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n478), .A2(G105), .A3(new_n476), .ZN(new_n778));
  AND4_X1   g353(.A1(new_n775), .A2(new_n776), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n772), .B1(new_n779), .B2(new_n735), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT27), .B(G1996), .Z(new_n781));
  AOI21_X1  g356(.A(new_n771), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n767), .B(new_n782), .C1(new_n780), .C2(new_n781), .ZN(new_n783));
  NOR2_X1   g358(.A1(G16), .A2(G19), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n564), .B2(G16), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1341), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n735), .A2(G26), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT28), .Z(new_n789));
  NAND2_X1  g364(.A1(new_n486), .A2(G128), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(KEYINPUT95), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(KEYINPUT95), .ZN(new_n792));
  MUX2_X1   g367(.A(G104), .B(G116), .S(G2105), .Z(new_n793));
  AOI22_X1  g368(.A1(new_n791), .A2(new_n792), .B1(G2104), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n483), .A2(G140), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT94), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n789), .B1(new_n797), .B2(G29), .ZN(new_n798));
  INV_X1    g373(.A(G2067), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(G16), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(G20), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT23), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n581), .B2(new_n801), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1956), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n800), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n735), .A2(G27), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G164), .B2(new_n735), .ZN(new_n808));
  INV_X1    g383(.A(G2078), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n787), .A2(new_n806), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n756), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(KEYINPUT99), .B1(G16), .B2(G21), .ZN(new_n813));
  NOR2_X1   g388(.A1(G286), .A2(new_n801), .ZN(new_n814));
  MUX2_X1   g389(.A(new_n813), .B(KEYINPUT99), .S(new_n814), .Z(new_n815));
  INV_X1    g390(.A(G1966), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n752), .A2(new_n753), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT101), .Z(new_n819));
  NAND2_X1  g394(.A1(new_n815), .A2(new_n816), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n812), .A2(new_n817), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n731), .A2(new_n821), .ZN(G311));
  INV_X1    g397(.A(G311), .ZN(G150));
  NAND2_X1  g398(.A1(new_n618), .A2(G559), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT38), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n527), .A2(G93), .ZN(new_n826));
  NAND2_X1  g401(.A1(G80), .A2(G543), .ZN(new_n827));
  INV_X1    g402(.A(G67), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n531), .B2(new_n828), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n829), .A2(G651), .B1(G55), .B2(new_n534), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(KEYINPUT102), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n826), .A2(new_n830), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT102), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n564), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n625), .A2(new_n834), .A3(new_n833), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n825), .B(new_n838), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n839), .A2(KEYINPUT39), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(KEYINPUT39), .ZN(new_n841));
  XOR2_X1   g416(.A(KEYINPUT103), .B(G860), .Z(new_n842));
  NAND3_X1  g417(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n831), .A2(new_n842), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT37), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(G145));
  XNOR2_X1  g421(.A(G162), .B(new_n750), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n639), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n797), .B(new_n506), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n722), .B(new_n632), .ZN(new_n850));
  MUX2_X1   g425(.A(G106), .B(G118), .S(G2105), .Z(new_n851));
  AOI22_X1  g426(.A1(new_n486), .A2(G130), .B1(G2104), .B2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(G142), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n852), .B1(new_n853), .B2(new_n638), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n850), .B(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n849), .B(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n779), .B(new_n765), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n848), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT104), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n848), .A2(new_n858), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n861), .A2(G37), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n860), .A2(KEYINPUT40), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(KEYINPUT40), .B1(new_n860), .B2(new_n862), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(G395));
  XNOR2_X1  g440(.A(new_n628), .B(new_n838), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n581), .B1(new_n610), .B2(new_n617), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT41), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n610), .A2(new_n581), .A3(new_n617), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n870), .ZN(new_n872));
  OAI21_X1  g447(.A(KEYINPUT41), .B1(new_n872), .B2(new_n867), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n866), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n702), .B(G303), .ZN(new_n875));
  XNOR2_X1  g450(.A(G290), .B(G288), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n875), .B(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n877), .A2(KEYINPUT105), .A3(KEYINPUT42), .ZN(new_n878));
  XNOR2_X1  g453(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n878), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n628), .A2(new_n838), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n628), .A2(new_n838), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n881), .B(new_n882), .C1(new_n867), .C2(new_n872), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n874), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(KEYINPUT106), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n874), .A2(new_n883), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n885), .B1(new_n886), .B2(new_n880), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n884), .A2(KEYINPUT106), .ZN(new_n888));
  OAI21_X1  g463(.A(G868), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n833), .A2(new_n605), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(G295));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n890), .ZN(G331));
  INV_X1    g467(.A(KEYINPUT43), .ZN(new_n893));
  INV_X1    g468(.A(G37), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n873), .A2(new_n871), .ZN(new_n895));
  NAND2_X1  g470(.A1(G168), .A2(G171), .ZN(new_n896));
  NAND2_X1  g471(.A1(G286), .A2(G301), .ZN(new_n897));
  AOI22_X1  g472(.A1(new_n896), .A2(new_n897), .B1(new_n836), .B2(new_n837), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT107), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n896), .A2(new_n836), .A3(new_n837), .A4(new_n897), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n902), .B1(new_n898), .B2(new_n899), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n895), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n896), .A2(new_n897), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n838), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n902), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n872), .A2(new_n867), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n904), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n894), .B1(new_n911), .B2(new_n877), .ZN(new_n912));
  INV_X1    g487(.A(new_n877), .ZN(new_n913));
  OAI211_X1 g488(.A(KEYINPUT108), .B(KEYINPUT41), .C1(new_n872), .C2(new_n867), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n907), .B(new_n914), .C1(new_n895), .C2(KEYINPUT108), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n906), .A2(KEYINPUT107), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n916), .A2(new_n909), .A3(new_n900), .A4(new_n902), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n913), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n893), .B1(new_n912), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n916), .A2(new_n900), .A3(new_n902), .ZN(new_n920));
  AOI22_X1  g495(.A1(new_n920), .A2(new_n895), .B1(new_n908), .B2(new_n909), .ZN(new_n921));
  AOI21_X1  g496(.A(G37), .B1(new_n921), .B2(new_n913), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n911), .A2(new_n877), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(KEYINPUT43), .A3(new_n923), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n919), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR3_X1   g502(.A1(new_n912), .A2(KEYINPUT109), .A3(new_n918), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT109), .ZN(new_n929));
  INV_X1    g504(.A(new_n918), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n929), .B1(new_n922), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT43), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n922), .A2(new_n893), .A3(new_n923), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT44), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT110), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT109), .B1(new_n912), .B2(new_n918), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n922), .A2(new_n930), .A3(new_n929), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n893), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT110), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n939), .A2(new_n940), .A3(new_n934), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n927), .B1(new_n936), .B2(new_n941), .ZN(G397));
  AOI21_X1  g517(.A(G1384), .B1(new_n509), .B2(new_n497), .ZN(new_n943));
  XNOR2_X1  g518(.A(KEYINPUT111), .B(KEYINPUT45), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G40), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n480), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n797), .B(new_n799), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n779), .B(G1996), .ZN(new_n952));
  OR2_X1    g527(.A1(new_n723), .A2(new_n726), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n723), .A2(new_n726), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n951), .A2(new_n952), .A3(new_n953), .A4(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(G290), .B(G1986), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n950), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT62), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT122), .ZN(new_n959));
  INV_X1    g534(.A(new_n948), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT50), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n960), .B1(new_n943), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(G1384), .B1(new_n508), .B2(new_n510), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n962), .B(new_n753), .C1(new_n963), .C2(new_n961), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n948), .B1(new_n943), .B2(KEYINPUT45), .ZN(new_n965));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n509), .A2(KEYINPUT73), .A3(new_n497), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT73), .B1(new_n509), .B2(new_n497), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n966), .B(new_n945), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT117), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n511), .A2(KEYINPUT117), .A3(new_n966), .A4(new_n945), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n965), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI211_X1 g548(.A(G168), .B(new_n964), .C1(new_n973), .C2(G1966), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(G8), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n964), .B1(new_n973), .B2(G1966), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(G286), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT51), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n981), .B1(new_n974), .B2(G8), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n959), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n981), .B1(new_n977), .B2(G286), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n985), .A2(new_n975), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n986), .A2(KEYINPUT122), .A3(new_n982), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n958), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n980), .A2(new_n959), .A3(new_n983), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT122), .B1(new_n986), .B2(new_n982), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n989), .A2(new_n990), .A3(KEYINPUT62), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n960), .B1(new_n943), .B2(KEYINPUT45), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(new_n963), .B2(new_n945), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G1971), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n992), .B(KEYINPUT112), .C1(new_n963), .C2(new_n945), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n506), .A2(new_n966), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n948), .B1(new_n999), .B2(KEYINPUT50), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1000), .B1(KEYINPUT50), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n740), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n998), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(G303), .A2(G8), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1005), .B(KEYINPUT55), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1004), .A2(G8), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT82), .B1(new_n595), .B2(G651), .ZN(new_n1009));
  AOI211_X1 g584(.A(new_n589), .B(new_n576), .C1(new_n593), .C2(new_n594), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(KEYINPUT114), .B(G86), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n520), .A2(new_n526), .A3(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1013), .A2(KEYINPUT115), .A3(new_n597), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT115), .B1(new_n1013), .B2(new_n597), .ZN(new_n1016));
  OAI21_X1  g591(.A(G1981), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OR2_X1    g592(.A1(G305), .A2(G1981), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n1017), .A2(KEYINPUT49), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT49), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1020));
  INV_X1    g595(.A(G8), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1021), .B1(new_n943), .B2(new_n948), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n1019), .A2(new_n1020), .A3(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n586), .B(G1976), .C1(new_n540), .C2(new_n587), .ZN(new_n1025));
  INV_X1    g600(.A(G1976), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT52), .B1(G288), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1022), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1029), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1028), .B1(new_n1030), .B2(KEYINPUT113), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n948), .A2(new_n506), .A3(new_n966), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1032), .A2(G8), .A3(new_n1025), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT113), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G288), .A2(new_n1026), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1033), .A2(new_n1034), .A3(new_n1029), .A4(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1031), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1024), .A2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n999), .A2(new_n961), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1039), .B1(new_n1001), .B2(new_n961), .ZN(new_n1040));
  OR3_X1    g615(.A1(new_n1040), .A2(G2090), .A3(new_n960), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1021), .B1(new_n998), .B2(new_n1041), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1008), .B(new_n1038), .C1(new_n1007), .C2(new_n1042), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n809), .A2(KEYINPUT53), .ZN(new_n1044));
  INV_X1    g619(.A(G1961), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n962), .B1(new_n963), .B2(new_n961), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n973), .A2(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(G2078), .B1(new_n995), .B2(new_n997), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1047), .B1(new_n1048), .B2(KEYINPUT53), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(G171), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1043), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n988), .A2(new_n991), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT126), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT126), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n988), .A2(new_n1054), .A3(new_n991), .A4(new_n1051), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT49), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1017), .A2(new_n1018), .A3(KEYINPUT49), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(new_n1060), .A3(new_n1022), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT116), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1061), .A2(new_n1062), .A3(new_n1031), .A4(new_n1036), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1032), .A2(G8), .A3(new_n1025), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT52), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1066), .A2(new_n1034), .B1(new_n1033), .B2(new_n1027), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1035), .ZN(new_n1068));
  NOR4_X1   g643(.A1(new_n1065), .A2(new_n1068), .A3(KEYINPUT113), .A4(KEYINPUT52), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1062), .B1(new_n1070), .B2(new_n1061), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1021), .B1(new_n998), .B2(new_n1003), .ZN(new_n1072));
  OAI22_X1  g647(.A1(new_n1064), .A2(new_n1071), .B1(new_n1072), .B2(new_n1007), .ZN(new_n1073));
  NOR2_X1   g648(.A1(G286), .A2(new_n1021), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n977), .A2(KEYINPUT63), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1008), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1073), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1004), .A2(G8), .ZN(new_n1079));
  OAI21_X1  g654(.A(KEYINPUT116), .B1(new_n1024), .B2(new_n1037), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n1079), .A2(new_n1006), .B1(new_n1080), .B2(new_n1063), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n977), .A2(KEYINPUT63), .A3(new_n1074), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1082), .B1(new_n1007), .B2(new_n1072), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT119), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1078), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT63), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n977), .A2(new_n1074), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1086), .B1(new_n1043), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT118), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g665(.A(KEYINPUT118), .B(new_n1086), .C1(new_n1043), .C2(new_n1087), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1085), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1008), .B1(new_n1080), .B2(new_n1063), .ZN(new_n1093));
  OR3_X1    g668(.A1(new_n1024), .A2(G1976), .A3(G288), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1023), .B1(new_n1094), .B2(new_n1018), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  OR2_X1    g671(.A1(new_n1048), .A2(KEYINPUT53), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1097), .A2(KEYINPUT124), .A3(G301), .A4(new_n1047), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT124), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1049), .B2(G171), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT54), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n1103));
  OAI21_X1  g678(.A(KEYINPUT53), .B1(new_n1103), .B2(G2078), .ZN(new_n1104));
  AOI211_X1 g679(.A(new_n1104), .B(new_n946), .C1(new_n1103), .C2(G2078), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1105), .A2(new_n992), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1097), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1102), .B1(new_n1107), .B2(G171), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT125), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1101), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1109), .B1(new_n1101), .B2(new_n1108), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(G1956), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1040), .B2(new_n960), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n581), .B(KEYINPUT57), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT56), .B(G2072), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n992), .B(new_n1116), .C1(new_n963), .C2(new_n945), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1114), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1115), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1119));
  INV_X1    g694(.A(G1348), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1032), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1046), .A2(new_n1120), .B1(new_n799), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n610), .A2(new_n617), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1118), .B1(new_n1119), .B2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1122), .A2(KEYINPUT60), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1121), .A2(new_n799), .ZN(new_n1128));
  OAI211_X1 g703(.A(KEYINPUT60), .B(new_n1128), .C1(new_n1002), .C2(G1348), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1127), .B1(new_n1129), .B2(new_n618), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1122), .A2(KEYINPUT120), .A3(KEYINPUT60), .A4(new_n1123), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1129), .A2(KEYINPUT121), .A3(new_n618), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT121), .B1(new_n1129), .B2(new_n618), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1126), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(KEYINPUT58), .B(G1341), .ZN(new_n1137));
  OAI22_X1  g712(.A1(new_n993), .A2(G1996), .B1(new_n1121), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n564), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT59), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT61), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1118), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1141), .B1(new_n1142), .B2(new_n1119), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1115), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1146), .A2(KEYINPUT61), .A3(new_n1118), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1140), .A2(new_n1143), .A3(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1125), .B1(new_n1136), .B2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(G301), .B(new_n1106), .C1(new_n1048), .C2(KEYINPUT53), .ZN(new_n1150));
  AOI21_X1  g725(.A(KEYINPUT54), .B1(new_n1050), .B2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1151), .A2(new_n1043), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1149), .A2(new_n990), .A3(new_n989), .A4(new_n1152), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1092), .B(new_n1096), .C1(new_n1112), .C2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n957), .B1(new_n1056), .B2(new_n1154), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n949), .A2(G1986), .A3(G290), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1156), .B(KEYINPUT48), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1157), .B1(new_n955), .B2(new_n950), .ZN(new_n1158));
  INV_X1    g733(.A(G1996), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT127), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1159), .B1(new_n1160), .B2(KEYINPUT46), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(KEYINPUT46), .ZN(new_n1162));
  OR3_X1    g737(.A1(new_n949), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1162), .B1(new_n949), .B2(new_n1161), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n951), .A2(new_n779), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1163), .B(new_n1164), .C1(new_n1165), .C2(new_n949), .ZN(new_n1166));
  XOR2_X1   g741(.A(new_n1166), .B(KEYINPUT47), .Z(new_n1167));
  NAND2_X1  g742(.A1(new_n951), .A2(new_n952), .ZN(new_n1168));
  OAI22_X1  g743(.A1(new_n1168), .A2(new_n954), .B1(G2067), .B2(new_n797), .ZN(new_n1169));
  AOI211_X1 g744(.A(new_n1158), .B(new_n1167), .C1(new_n950), .C2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1155), .A2(new_n1170), .ZN(G329));
  assign    G231 = 1'b0;
  OR4_X1    g746(.A1(new_n461), .A2(G229), .A3(G401), .A4(G227), .ZN(new_n1173));
  AOI21_X1  g747(.A(new_n1173), .B1(new_n860), .B2(new_n862), .ZN(new_n1174));
  AND2_X1   g748(.A1(new_n1174), .A2(new_n925), .ZN(G308));
  NAND2_X1  g749(.A1(new_n1174), .A2(new_n925), .ZN(G225));
endmodule


