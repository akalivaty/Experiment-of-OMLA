//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 1 1 0 1 0 0 0 0 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n540, new_n541, new_n542, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n559, new_n560, new_n561, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n598, new_n601, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1155, new_n1156;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT66), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n452), .A2(new_n457), .B1(new_n458), .B2(new_n453), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT67), .Z(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  AOI22_X1  g036(.A1(new_n461), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n461), .A2(new_n463), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n464), .A2(new_n470), .ZN(G160));
  AND2_X1   g046(.A1(new_n461), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G124), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n463), .A2(G112), .ZN(new_n474));
  OAI21_X1  g049(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n468), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(G136), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT68), .ZN(G162));
  OAI21_X1  g054(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n482));
  OAI21_X1  g057(.A(G2105), .B1(new_n482), .B2(G114), .ZN(new_n483));
  INV_X1    g058(.A(G114), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(KEYINPUT69), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n481), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  AND2_X1   g061(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n487));
  NOR2_X1   g062(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n488));
  OAI211_X1 g063(.A(G126), .B(G2105), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g065(.A(G138), .B(new_n463), .C1(new_n487), .C2(new_n488), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n461), .A2(new_n493), .A3(G138), .A4(new_n463), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n490), .B1(new_n492), .B2(new_n494), .ZN(G164));
  INV_X1    g070(.A(G543), .ZN(new_n496));
  NAND2_X1  g071(.A1(KEYINPUT70), .A2(G651), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT6), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(KEYINPUT70), .A2(KEYINPUT6), .A3(G651), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n496), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G50), .ZN(new_n502));
  INV_X1    g077(.A(G88), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n499), .A2(new_n500), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(new_n496), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n502), .B1(new_n503), .B2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n510), .A2(new_n513), .ZN(G303));
  INV_X1    g089(.A(G303), .ZN(G166));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT7), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n504), .A2(G543), .ZN(new_n519));
  XOR2_X1   g094(.A(KEYINPUT71), .B(G51), .Z(new_n520));
  OAI211_X1 g095(.A(new_n517), .B(new_n518), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT72), .B(G89), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n509), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n521), .A2(new_n523), .ZN(G168));
  AOI22_X1  g099(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n504), .A2(new_n508), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n526), .A2(G651), .B1(new_n527), .B2(G90), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n501), .A2(G52), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(G301));
  INV_X1    g105(.A(G301), .ZN(G171));
  AOI22_X1  g106(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n532), .A2(new_n512), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n501), .A2(G43), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n527), .A2(G81), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G860), .ZN(G153));
  NAND4_X1  g113(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g114(.A1(G1), .A2(G3), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT8), .ZN(new_n541));
  NAND4_X1  g116(.A1(G319), .A2(G483), .A3(G661), .A4(new_n541), .ZN(new_n542));
  XOR2_X1   g117(.A(new_n542), .B(KEYINPUT73), .Z(G188));
  INV_X1    g118(.A(G65), .ZN(new_n544));
  INV_X1    g119(.A(new_n508), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT74), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n508), .A2(KEYINPUT74), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n544), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g124(.A1(G78), .A2(G543), .ZN(new_n550));
  OAI21_X1  g125(.A(G651), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(G53), .ZN(new_n552));
  OAI21_X1  g127(.A(KEYINPUT9), .B1(new_n519), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT9), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n501), .A2(new_n554), .A3(G53), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n553), .A2(new_n555), .B1(G91), .B2(new_n527), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n551), .A2(new_n556), .ZN(G299));
  INV_X1    g132(.A(G168), .ZN(G286));
  NAND2_X1  g133(.A1(new_n527), .A2(G87), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n501), .A2(G49), .ZN(new_n560));
  OAI21_X1  g135(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(G288));
  NAND2_X1  g137(.A1(G73), .A2(G543), .ZN(new_n563));
  OR2_X1    g138(.A1(new_n563), .A2(KEYINPUT75), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(KEYINPUT75), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(G61), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(new_n506), .B2(new_n507), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n501), .A2(G48), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(G86), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT76), .B1(new_n509), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n504), .A2(new_n508), .A3(new_n574), .A4(G86), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n571), .A2(new_n576), .ZN(G305));
  AOI22_X1  g152(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  OR3_X1    g153(.A1(new_n578), .A2(KEYINPUT77), .A3(new_n512), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT77), .B1(new_n578), .B2(new_n512), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n527), .A2(G85), .B1(G47), .B2(new_n501), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(G290));
  NAND2_X1  g157(.A1(G301), .A2(G868), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n527), .A2(G92), .ZN(new_n584));
  XOR2_X1   g159(.A(new_n584), .B(KEYINPUT10), .Z(new_n585));
  INV_X1    g160(.A(G79), .ZN(new_n586));
  OAI21_X1  g161(.A(KEYINPUT78), .B1(new_n586), .B2(new_n496), .ZN(new_n587));
  OR3_X1    g162(.A1(new_n586), .A2(new_n496), .A3(KEYINPUT78), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n508), .B(new_n546), .ZN(new_n589));
  INV_X1    g164(.A(G66), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n587), .B(new_n588), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(G54), .B2(new_n501), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n585), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n583), .B1(new_n594), .B2(G868), .ZN(G321));
  XNOR2_X1  g170(.A(G321), .B(KEYINPUT79), .ZN(G284));
  INV_X1    g171(.A(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(G299), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(new_n597), .B2(G168), .ZN(G297));
  OAI21_X1  g174(.A(new_n598), .B1(new_n597), .B2(G168), .ZN(G280));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n594), .B1(new_n601), .B2(G860), .ZN(G148));
  NAND2_X1  g177(.A1(new_n536), .A2(new_n597), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n593), .A2(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(new_n597), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g181(.A1(new_n461), .A2(new_n466), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT12), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT13), .ZN(new_n609));
  INV_X1    g184(.A(G2100), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI22_X1  g186(.A1(G135), .A2(new_n477), .B1(new_n472), .B2(G123), .ZN(new_n612));
  OAI21_X1  g187(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n613));
  INV_X1    g188(.A(G111), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n613), .A2(KEYINPUT80), .B1(new_n614), .B2(G2105), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(KEYINPUT80), .B2(new_n613), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(G2096), .Z(new_n618));
  NAND2_X1  g193(.A1(new_n609), .A2(new_n610), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n611), .A2(new_n618), .A3(new_n619), .ZN(G156));
  XOR2_X1   g195(.A(G2443), .B(G2446), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT82), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2451), .ZN(new_n623));
  XNOR2_X1  g198(.A(G1341), .B(G1348), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2427), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT15), .B(G2435), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n629), .A2(new_n630), .A3(KEYINPUT14), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n625), .B(new_n631), .Z(new_n632));
  XOR2_X1   g207(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2454), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n632), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(new_n636), .A3(G14), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(G401));
  XOR2_X1   g213(.A(G2072), .B(G2078), .Z(new_n639));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  XNOR2_X1  g215(.A(G2067), .B(G2678), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n639), .B1(new_n642), .B2(KEYINPUT18), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT83), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2100), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT18), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n642), .A2(KEYINPUT17), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n640), .A2(new_n641), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2096), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n645), .B(new_n650), .ZN(G227));
  XOR2_X1   g226(.A(KEYINPUT84), .B(KEYINPUT19), .Z(new_n652));
  XNOR2_X1  g227(.A(G1971), .B(G1976), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1956), .B(G2474), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1961), .B(G1966), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT20), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n655), .A2(new_n656), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n654), .A2(new_n661), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n657), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n659), .B(new_n662), .C1(new_n654), .C2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1991), .B(G1996), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1981), .B(G1986), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G229));
  MUX2_X1   g245(.A(G6), .B(G305), .S(G16), .Z(new_n671));
  XOR2_X1   g246(.A(KEYINPUT32), .B(G1981), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(G16), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(G22), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(G166), .B2(new_n674), .ZN(new_n676));
  INV_X1    g251(.A(G1971), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n674), .A2(G23), .ZN(new_n679));
  INV_X1    g254(.A(G288), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n679), .B1(new_n680), .B2(new_n674), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT33), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n673), .A2(new_n678), .A3(new_n683), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n684), .A2(KEYINPUT34), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(KEYINPUT34), .ZN(new_n686));
  INV_X1    g261(.A(G29), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G25), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT85), .Z(new_n689));
  OAI21_X1  g264(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(G107), .B2(new_n463), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT86), .ZN(new_n693));
  AOI22_X1  g268(.A1(G131), .A2(new_n477), .B1(new_n472), .B2(G119), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n689), .B1(new_n695), .B2(G29), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT87), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT35), .B(G1991), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(G16), .A2(G24), .ZN(new_n700));
  INV_X1    g275(.A(G290), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(G16), .ZN(new_n702));
  INV_X1    g277(.A(G1986), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND4_X1  g279(.A1(new_n685), .A2(new_n686), .A3(new_n699), .A4(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT36), .Z(new_n706));
  NOR2_X1   g281(.A1(G29), .A2(G35), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G162), .B2(G29), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT29), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n709), .A2(G2090), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(G2090), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT90), .B(KEYINPUT23), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n674), .A2(G20), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G299), .B2(G16), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G1956), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n710), .A2(new_n711), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n674), .A2(G4), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(new_n594), .B2(new_n674), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(G1348), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(G1348), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n674), .A2(G21), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G168), .B2(new_n674), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n723), .A2(G1966), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT89), .Z(new_n725));
  NAND3_X1  g300(.A1(new_n720), .A2(new_n721), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n687), .A2(G33), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n461), .A2(G127), .ZN(new_n728));
  NAND2_X1  g303(.A1(G115), .A2(G2104), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n463), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT25), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI211_X1 g310(.A(new_n730), .B(new_n735), .C1(G139), .C2(new_n477), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n727), .B1(new_n736), .B2(new_n687), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G2072), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n477), .A2(G140), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n472), .A2(G128), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n463), .A2(G116), .ZN(new_n741));
  OAI21_X1  g316(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n739), .B(new_n740), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G29), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n687), .A2(G26), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT28), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G2067), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n472), .A2(G129), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT88), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n477), .A2(G141), .ZN(new_n752));
  NAND3_X1  g327(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT26), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n466), .A2(G105), .ZN(new_n755));
  AND4_X1   g330(.A1(new_n751), .A2(new_n752), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n756), .A2(new_n687), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n687), .B2(G32), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT27), .B(G1996), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n749), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AOI211_X1 g335(.A(new_n738), .B(new_n760), .C1(G1966), .C2(new_n723), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT24), .ZN(new_n762));
  INV_X1    g337(.A(G34), .ZN(new_n763));
  AOI21_X1  g338(.A(G29), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n762), .B2(new_n763), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G160), .B2(new_n687), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n766), .A2(G2084), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n766), .A2(G2084), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT30), .B(G28), .ZN(new_n769));
  OR2_X1    g344(.A1(KEYINPUT31), .A2(G11), .ZN(new_n770));
  NAND2_X1  g345(.A1(KEYINPUT31), .A2(G11), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n769), .A2(new_n687), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n617), .B2(new_n687), .ZN(new_n773));
  NOR3_X1   g348(.A1(new_n767), .A2(new_n768), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G16), .A2(G19), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n537), .B2(G16), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G1341), .ZN(new_n777));
  NOR2_X1   g352(.A1(G171), .A2(new_n674), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G5), .B2(new_n674), .ZN(new_n779));
  INV_X1    g354(.A(G1961), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI211_X1 g356(.A(new_n777), .B(new_n781), .C1(new_n758), .C2(new_n759), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n687), .A2(G27), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G164), .B2(new_n687), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G2078), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n779), .B2(new_n780), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n761), .A2(new_n774), .A3(new_n782), .A4(new_n786), .ZN(new_n787));
  NOR4_X1   g362(.A1(new_n706), .A2(new_n717), .A3(new_n726), .A4(new_n787), .ZN(G311));
  INV_X1    g363(.A(G311), .ZN(G150));
  AOI22_X1  g364(.A1(new_n527), .A2(G93), .B1(G55), .B2(new_n501), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT92), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n792), .B1(new_n512), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n794), .A2(G860), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT93), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT37), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n593), .A2(new_n601), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT91), .B(KEYINPUT38), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n794), .A2(new_n536), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n794), .A2(new_n536), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n800), .B(new_n803), .Z(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n805), .A2(KEYINPUT39), .ZN(new_n806));
  INV_X1    g381(.A(G860), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n805), .B2(KEYINPUT39), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n797), .B1(new_n806), .B2(new_n808), .ZN(G145));
  NAND2_X1  g384(.A1(new_n477), .A2(G142), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n472), .A2(G130), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n463), .A2(G118), .ZN(new_n812));
  OAI21_X1  g387(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n810), .B(new_n811), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT97), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(new_n695), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n608), .B(KEYINPUT96), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(KEYINPUT98), .ZN(new_n819));
  INV_X1    g394(.A(new_n489), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n463), .B1(KEYINPUT69), .B2(new_n484), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n482), .A2(G114), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n480), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(KEYINPUT95), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n492), .A2(new_n494), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT95), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n486), .A2(new_n826), .A3(new_n489), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n824), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n743), .B(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n756), .B(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(new_n736), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n819), .B(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(G160), .B(KEYINPUT94), .ZN(new_n833));
  XNOR2_X1  g408(.A(G162), .B(new_n833), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(new_n617), .Z(new_n835));
  NOR2_X1   g410(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(G37), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n831), .A2(new_n818), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n831), .A2(new_n818), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n837), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n836), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(G395));
  NAND2_X1  g419(.A1(new_n794), .A2(new_n597), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n594), .A2(G299), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n593), .B1(new_n551), .B2(new_n556), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT41), .ZN(new_n849));
  NOR3_X1   g424(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n846), .A2(KEYINPUT100), .ZN(new_n851));
  INV_X1    g426(.A(new_n847), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT100), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(new_n594), .B2(G299), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n851), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n850), .B1(new_n855), .B2(new_n849), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n803), .B(new_n604), .ZN(new_n857));
  MUX2_X1   g432(.A(new_n848), .B(new_n856), .S(new_n857), .Z(new_n858));
  XOR2_X1   g433(.A(G290), .B(G305), .Z(new_n859));
  XNOR2_X1  g434(.A(G303), .B(G288), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT42), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n858), .B(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n845), .B1(new_n863), .B2(new_n597), .ZN(G295));
  OAI21_X1  g439(.A(new_n845), .B1(new_n863), .B2(new_n597), .ZN(G331));
  INV_X1    g440(.A(KEYINPUT43), .ZN(new_n866));
  AOI21_X1  g441(.A(G301), .B1(new_n801), .B2(new_n802), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n801), .A2(G301), .A3(new_n802), .ZN(new_n869));
  AOI21_X1  g444(.A(G168), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n869), .ZN(new_n871));
  NOR3_X1   g446(.A1(new_n871), .A2(G286), .A3(new_n867), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n848), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n861), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n874), .A2(KEYINPUT101), .ZN(new_n875));
  OAI21_X1  g450(.A(G286), .B1(new_n871), .B2(new_n867), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n868), .A2(G168), .A3(new_n869), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n856), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n873), .A2(new_n875), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(new_n837), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n875), .B1(new_n873), .B2(new_n878), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n866), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n873), .A2(new_n878), .ZN(new_n883));
  AOI21_X1  g458(.A(G37), .B1(new_n883), .B2(new_n874), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n876), .A2(new_n877), .A3(KEYINPUT41), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n874), .B1(new_n885), .B2(new_n848), .ZN(new_n886));
  INV_X1    g461(.A(new_n855), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n886), .B1(new_n887), .B2(new_n885), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n882), .B1(new_n889), .B2(new_n866), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(KEYINPUT44), .ZN(new_n891));
  OAI21_X1  g466(.A(KEYINPUT43), .B1(new_n880), .B2(new_n881), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(new_n889), .B2(KEYINPUT43), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n891), .A2(new_n895), .ZN(G397));
  INV_X1    g471(.A(KEYINPUT61), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT57), .B1(G299), .B2(KEYINPUT114), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT114), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT57), .ZN(new_n900));
  AOI211_X1 g475(.A(new_n899), .B(new_n900), .C1(new_n551), .C2(new_n556), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT106), .ZN(new_n903));
  INV_X1    g478(.A(G1384), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n828), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n903), .B1(new_n828), .B2(new_n904), .ZN(new_n906));
  OAI21_X1  g481(.A(KEYINPUT50), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(G40), .ZN(new_n908));
  NOR3_X1   g483(.A1(new_n464), .A2(new_n470), .A3(new_n908), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n492), .A2(new_n494), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n904), .B1(new_n910), .B2(new_n490), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n909), .B1(new_n911), .B2(KEYINPUT50), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(G1956), .B1(new_n907), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(KEYINPUT102), .B(KEYINPUT45), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n828), .A2(KEYINPUT45), .A3(new_n904), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(new_n918), .A3(new_n909), .ZN(new_n919));
  XNOR2_X1  g494(.A(KEYINPUT56), .B(G2072), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n902), .B1(new_n915), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n825), .A2(new_n827), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n826), .B1(new_n486), .B2(new_n489), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n904), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT106), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n828), .A2(new_n903), .A3(new_n904), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n912), .B1(new_n929), .B2(KEYINPUT50), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n922), .B(new_n902), .C1(new_n930), .C2(G1956), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n897), .B1(new_n923), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n919), .A2(new_n921), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT115), .B1(new_n914), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT115), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n922), .B(new_n936), .C1(new_n930), .C2(G1956), .ZN(new_n937));
  OR2_X1    g512(.A1(new_n898), .A2(new_n901), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n935), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n914), .A2(new_n934), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n897), .B1(new_n940), .B2(new_n902), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  XOR2_X1   g517(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n943));
  XOR2_X1   g518(.A(KEYINPUT117), .B(G1996), .Z(new_n944));
  NOR2_X1   g519(.A1(new_n919), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n927), .A2(new_n909), .A3(new_n928), .ZN(new_n946));
  XOR2_X1   g521(.A(KEYINPUT58), .B(G1341), .Z(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n945), .B1(new_n948), .B2(KEYINPUT118), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT118), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n946), .A2(new_n950), .A3(new_n947), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n943), .B1(new_n952), .B2(new_n537), .ZN(new_n953));
  INV_X1    g528(.A(new_n943), .ZN(new_n954));
  AOI211_X1 g529(.A(new_n536), .B(new_n954), .C1(new_n949), .C2(new_n951), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n933), .B(new_n942), .C1(new_n953), .C2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n909), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT50), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n927), .A2(new_n958), .A3(new_n928), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT107), .B1(new_n911), .B2(KEYINPUT50), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n957), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT107), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n927), .A2(new_n963), .A3(new_n958), .A4(new_n928), .ZN(new_n964));
  AOI21_X1  g539(.A(G1348), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n946), .A2(G2067), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT60), .B1(new_n593), .B2(KEYINPUT120), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n593), .A2(KEYINPUT120), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  NOR4_X1   g544(.A1(new_n965), .A2(new_n966), .A3(new_n967), .A4(new_n969), .ZN(new_n970));
  OR3_X1    g545(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n905), .A2(new_n906), .A3(KEYINPUT50), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n909), .B(new_n964), .C1(new_n972), .C2(new_n960), .ZN(new_n973));
  INV_X1    g548(.A(G1348), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n966), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n968), .B1(new_n975), .B2(KEYINPUT60), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n970), .B1(new_n971), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT116), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n931), .B(new_n594), .C1(new_n965), .C2(new_n966), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n978), .B1(new_n979), .B2(new_n939), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n979), .A2(new_n978), .A3(new_n939), .ZN(new_n981));
  OAI22_X1  g556(.A1(new_n956), .A2(new_n977), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT121), .ZN(new_n983));
  INV_X1    g558(.A(G8), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n959), .A2(new_n961), .ZN(new_n985));
  XNOR2_X1  g560(.A(KEYINPUT113), .B(G2084), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n985), .A2(new_n909), .A3(new_n964), .A4(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1966), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT45), .B1(new_n927), .B2(new_n928), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n909), .B1(new_n911), .B2(new_n916), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n984), .B1(new_n987), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT51), .B1(new_n992), .B2(KEYINPUT122), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n987), .A2(G168), .A3(new_n991), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n994), .A2(G8), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(G8), .ZN(new_n997));
  AOI21_X1  g572(.A(G168), .B1(new_n987), .B2(new_n991), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n996), .B1(new_n993), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n680), .A2(G1976), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n946), .A2(G8), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT52), .ZN(new_n1003));
  XNOR2_X1  g578(.A(KEYINPUT109), .B(G1976), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT52), .B1(G288), .B2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n946), .A2(G8), .A3(new_n1001), .A4(new_n1005), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1981), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n571), .A2(new_n576), .A3(new_n1008), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n569), .B(new_n570), .C1(new_n572), .C2(new_n509), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(G1981), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT49), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1009), .A2(new_n1011), .A3(KEYINPUT49), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1014), .A2(new_n946), .A3(G8), .A4(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT110), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n1009), .A2(new_n1011), .A3(KEYINPUT49), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT49), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT110), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1020), .A2(new_n1021), .A3(G8), .A4(new_n946), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1017), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G2090), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n930), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n919), .A2(KEYINPUT105), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT105), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n917), .A2(new_n918), .A3(new_n1027), .A4(new_n909), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1026), .A2(new_n677), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n984), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(G303), .A2(G8), .ZN(new_n1031));
  XOR2_X1   g606(.A(new_n1031), .B(KEYINPUT55), .Z(new_n1032));
  OAI211_X1 g607(.A(new_n1007), .B(new_n1023), .C1(new_n1030), .C2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n962), .A2(KEYINPUT108), .A3(new_n1024), .A4(new_n964), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n1029), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n962), .A2(new_n1024), .A3(new_n964), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT108), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n984), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1033), .B1(new_n1040), .B2(new_n1032), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1042));
  INV_X1    g617(.A(G2078), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n973), .A2(new_n780), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n989), .A2(new_n990), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1048), .A2(KEYINPUT53), .A3(new_n1043), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1047), .A2(KEYINPUT124), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT124), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1051));
  OAI211_X1 g626(.A(G301), .B(new_n1046), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1043), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1054));
  INV_X1    g629(.A(new_n462), .ZN(new_n1055));
  OR2_X1    g630(.A1(new_n1055), .A2(KEYINPUT125), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n463), .B1(new_n1055), .B2(KEYINPUT125), .ZN(new_n1057));
  AOI211_X1 g632(.A(new_n470), .B(new_n1054), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n926), .A2(new_n916), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1058), .A2(new_n918), .A3(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1046), .A2(new_n1047), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1053), .B1(new_n1061), .B2(G171), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1052), .A2(new_n1062), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1000), .A2(new_n1041), .A3(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT123), .B(KEYINPUT54), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1046), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n1066), .A2(G171), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1061), .A2(G171), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1065), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n1070));
  OAI221_X1 g645(.A(new_n1070), .B1(new_n981), .B2(new_n980), .C1(new_n956), .C2(new_n977), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n983), .A2(new_n1064), .A3(new_n1069), .A4(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1033), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1074));
  OAI211_X1 g649(.A(G8), .B(new_n1032), .C1(new_n1074), .C2(new_n1035), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1066), .A2(new_n1073), .A3(G171), .A4(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n999), .A2(new_n993), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n987), .A2(new_n991), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(G8), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT122), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n997), .B1(new_n1081), .B2(KEYINPUT51), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1077), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT62), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1076), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT62), .B1(new_n1077), .B2(new_n1082), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(KEYINPUT126), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT126), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1000), .A2(new_n1088), .A3(KEYINPUT62), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1085), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT112), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1007), .A2(new_n1023), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT111), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1007), .A2(new_n1023), .A3(KEYINPUT111), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1075), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(G1976), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1023), .A2(new_n1097), .A3(new_n680), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n1009), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n946), .A2(G8), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1091), .B1(new_n1096), .B2(new_n1102), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1104));
  OAI211_X1 g679(.A(KEYINPUT112), .B(new_n1101), .C1(new_n1104), .C2(new_n1075), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT63), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1106), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1079), .A2(G286), .ZN(new_n1108));
  OAI21_X1  g683(.A(G8), .B1(new_n1074), .B2(new_n1035), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1032), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1107), .A2(new_n1075), .A3(new_n1108), .A4(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1108), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1106), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1103), .A2(new_n1105), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1072), .A2(new_n1090), .A3(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1059), .A2(new_n957), .ZN(new_n1118));
  INV_X1    g693(.A(G1996), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  XOR2_X1   g695(.A(new_n1120), .B(KEYINPUT104), .Z(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n743), .B(new_n748), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n756), .B2(new_n1119), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1122), .A2(new_n756), .B1(new_n1118), .B2(new_n1124), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n695), .A2(new_n698), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n695), .A2(new_n698), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1118), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1118), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n701), .A2(new_n703), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1132), .B(KEYINPUT103), .ZN(new_n1133));
  NAND2_X1  g708(.A1(G290), .A2(G1986), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1131), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1130), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1117), .A2(new_n1136), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1121), .A2(KEYINPUT46), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1121), .A2(KEYINPUT46), .ZN(new_n1139));
  AND2_X1   g714(.A1(new_n756), .A2(new_n1123), .ZN(new_n1140));
  OAI22_X1  g715(.A1(new_n1138), .A2(new_n1139), .B1(new_n1131), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT47), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1143), .A2(KEYINPUT127), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT127), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1133), .A2(new_n1131), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(KEYINPUT48), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n743), .A2(G2067), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1149), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1150));
  OAI22_X1  g725(.A1(new_n1130), .A2(new_n1148), .B1(new_n1131), .B2(new_n1150), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n1145), .A2(new_n1146), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1137), .A2(new_n1152), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g728(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1155));
  NOR3_X1   g729(.A1(new_n842), .A2(G229), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g730(.A1(new_n1156), .A2(new_n893), .ZN(G225));
  INV_X1    g731(.A(G225), .ZN(G308));
endmodule


