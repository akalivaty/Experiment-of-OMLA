//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n543, new_n544, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n591, new_n592, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT65), .Z(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n466), .A2(new_n469), .B1(G101), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n473), .B1(new_n464), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT66), .B(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  NOR2_X1   g054(.A1(new_n464), .A2(new_n469), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n464), .A2(G2105), .ZN(new_n481));
  AOI22_X1  g056(.A1(G124), .A2(new_n480), .B1(new_n481), .B2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT67), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(new_n469), .B2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n490));
  AND2_X1   g065(.A1(G126), .A2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(new_n462), .B2(new_n463), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G138), .B1(new_n462), .B2(new_n463), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT4), .B1(new_n494), .B2(new_n476), .ZN(new_n495));
  XNOR2_X1  g070(.A(KEYINPUT3), .B(G2104), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n469), .A2(new_n496), .A3(new_n497), .A4(G138), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n493), .B1(new_n495), .B2(new_n498), .ZN(G164));
  NAND2_X1  g074(.A1(G75), .A2(G543), .ZN(new_n500));
  XOR2_X1   g075(.A(KEYINPUT5), .B(G543), .Z(new_n501));
  INV_X1    g076(.A(G62), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT68), .B(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(new_n505), .B(KEYINPUT69), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n507), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G50), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n501), .B1(new_n508), .B2(new_n510), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n506), .A2(new_n516), .ZN(G166));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT70), .ZN(new_n519));
  XOR2_X1   g094(.A(new_n519), .B(KEYINPUT7), .Z(new_n520));
  AOI21_X1  g095(.A(new_n520), .B1(G51), .B2(new_n511), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT5), .B(G543), .ZN(new_n522));
  AND2_X1   g097(.A1(G63), .A2(G651), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n513), .A2(G89), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n521), .A2(new_n524), .ZN(G286));
  INV_X1    g100(.A(G286), .ZN(G168));
  XNOR2_X1  g101(.A(KEYINPUT71), .B(G90), .ZN(new_n527));
  AOI22_X1  g102(.A1(G52), .A2(new_n511), .B1(new_n513), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT72), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  XOR2_X1   g105(.A(KEYINPUT68), .B(G651), .Z(new_n531));
  OR2_X1    g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n529), .A2(new_n532), .ZN(G301));
  INV_X1    g108(.A(G301), .ZN(G171));
  NAND2_X1  g109(.A1(new_n513), .A2(G81), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n511), .A2(G43), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n522), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(new_n531), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n535), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  NAND4_X1  g116(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND4_X1  g119(.A1(G319), .A2(G483), .A3(G661), .A4(new_n544), .ZN(G188));
  NAND2_X1  g120(.A1(new_n511), .A2(G53), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT9), .ZN(new_n547));
  NAND2_X1  g122(.A1(G78), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G65), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n501), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n513), .A2(G91), .B1(new_n550), .B2(G651), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n547), .A2(new_n551), .ZN(G299));
  INV_X1    g127(.A(G166), .ZN(G303));
  INV_X1    g128(.A(G651), .ZN(new_n554));
  INV_X1    g129(.A(G74), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n554), .B1(new_n501), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n556), .B1(new_n513), .B2(G87), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n511), .A2(G49), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(G288));
  AOI21_X1  g134(.A(KEYINPUT73), .B1(new_n522), .B2(G61), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n560), .B1(G73), .B2(G543), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n522), .A2(KEYINPUT73), .A3(G61), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(new_n504), .ZN(new_n564));
  AOI22_X1  g139(.A1(G48), .A2(new_n511), .B1(new_n513), .B2(G86), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n564), .A2(new_n565), .A3(KEYINPUT74), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT74), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n511), .A2(G48), .ZN(new_n568));
  INV_X1    g143(.A(G86), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n514), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n531), .B1(new_n561), .B2(new_n562), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n567), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AND2_X1   g147(.A1(new_n566), .A2(new_n572), .ZN(G305));
  AOI22_X1  g148(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n574), .A2(new_n531), .ZN(new_n575));
  XOR2_X1   g150(.A(new_n575), .B(KEYINPUT75), .Z(new_n576));
  AOI22_X1  g151(.A1(G47), .A2(new_n511), .B1(new_n513), .B2(G85), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(G290));
  NAND2_X1  g153(.A1(new_n513), .A2(G92), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT10), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n579), .B(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(G79), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G66), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n501), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n511), .A2(G54), .B1(new_n584), .B2(G651), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(G868), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n588), .B1(G171), .B2(new_n587), .ZN(G284));
  OAI21_X1  g164(.A(new_n588), .B1(G171), .B2(new_n587), .ZN(G321));
  NAND2_X1  g165(.A1(G286), .A2(G868), .ZN(new_n591));
  INV_X1    g166(.A(G299), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n592), .B2(G868), .ZN(G297));
  OAI21_X1  g168(.A(new_n591), .B1(new_n592), .B2(G868), .ZN(G280));
  INV_X1    g169(.A(new_n586), .ZN(new_n595));
  INV_X1    g170(.A(G559), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(G860), .ZN(G148));
  OAI21_X1  g172(.A(KEYINPUT76), .B1(new_n540), .B2(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n595), .A2(new_n596), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(G868), .ZN(new_n600));
  MUX2_X1   g175(.A(KEYINPUT76), .B(new_n598), .S(new_n600), .Z(G323));
  XNOR2_X1  g176(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g177(.A1(new_n496), .A2(new_n471), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT12), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT13), .ZN(new_n605));
  INV_X1    g180(.A(G2100), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n605), .A2(new_n606), .ZN(new_n608));
  AOI22_X1  g183(.A1(G123), .A2(new_n480), .B1(new_n481), .B2(G135), .ZN(new_n609));
  OAI221_X1 g184(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n469), .C2(G111), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(G2096), .Z(new_n612));
  NAND3_X1  g187(.A1(new_n607), .A2(new_n608), .A3(new_n612), .ZN(G156));
  XNOR2_X1  g188(.A(G2427), .B(G2430), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT78), .ZN(new_n615));
  XNOR2_X1  g190(.A(KEYINPUT77), .B(G2438), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n615), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT15), .B(G2435), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n615), .B(new_n616), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(new_n619), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n621), .A2(new_n623), .A3(KEYINPUT14), .ZN(new_n624));
  XOR2_X1   g199(.A(G2451), .B(G2454), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT16), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n624), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G2443), .B(G2446), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G1341), .B(G1348), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT79), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(G14), .B1(new_n629), .B2(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(KEYINPUT80), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n634), .B1(new_n629), .B2(new_n632), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n629), .A2(new_n634), .A3(new_n632), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n633), .B1(new_n636), .B2(new_n637), .ZN(G401));
  XNOR2_X1  g213(.A(G2072), .B(G2078), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT17), .Z(new_n640));
  XNOR2_X1  g215(.A(G2067), .B(G2678), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n641), .B2(new_n639), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT81), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n644), .A2(new_n641), .A3(new_n639), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT18), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n645), .A2(new_n641), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n650), .B1(new_n640), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2096), .B(G2100), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(G227));
  XOR2_X1   g230(.A(KEYINPUT82), .B(KEYINPUT19), .Z(new_n656));
  XNOR2_X1  g231(.A(G1971), .B(G1976), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1956), .B(G2474), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1961), .B(G1966), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT83), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OR3_X1    g238(.A1(new_n659), .A2(new_n660), .A3(new_n662), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n658), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT20), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n659), .A2(new_n660), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n661), .A2(new_n667), .ZN(new_n668));
  MUX2_X1   g243(.A(new_n668), .B(new_n667), .S(new_n658), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G1981), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT84), .ZN(new_n673));
  XOR2_X1   g248(.A(G1991), .B(G1996), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n671), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT85), .B(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(G229));
  NAND3_X1  g254(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT93), .B(KEYINPUT25), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n481), .A2(G139), .ZN(new_n683));
  AOI22_X1  g258(.A1(new_n496), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n682), .B(new_n683), .C1(new_n469), .C2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT94), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G29), .ZN(new_n687));
  INV_X1    g262(.A(G29), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G33), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n690), .A2(G2072), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT95), .Z(new_n692));
  AND2_X1   g267(.A1(new_n688), .A2(G32), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n480), .A2(G129), .ZN(new_n694));
  NAND3_X1  g269(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT26), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n481), .A2(G141), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n471), .A2(G105), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n693), .B1(new_n701), .B2(G29), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT27), .B(G1996), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT96), .ZN(new_n705));
  INV_X1    g280(.A(G2084), .ZN(new_n706));
  INV_X1    g281(.A(G34), .ZN(new_n707));
  AOI21_X1  g282(.A(G29), .B1(new_n707), .B2(KEYINPUT24), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(KEYINPUT24), .B2(new_n707), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(new_n478), .B2(new_n688), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n705), .B1(new_n706), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G2072), .B2(new_n690), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n692), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT97), .Z(new_n714));
  NAND2_X1  g289(.A1(new_n688), .A2(G35), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G162), .B2(new_n688), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT29), .Z(new_n717));
  INV_X1    g292(.A(G2090), .ZN(new_n718));
  NOR2_X1   g293(.A1(G16), .A2(G19), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n540), .B2(G16), .ZN(new_n720));
  AOI22_X1  g295(.A1(new_n717), .A2(new_n718), .B1(G1341), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT31), .B(G11), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT30), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n723), .A2(G28), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n688), .B1(new_n723), .B2(G28), .ZN(new_n725));
  OAI221_X1 g300(.A(new_n722), .B1(new_n724), .B2(new_n725), .C1(new_n611), .C2(new_n688), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n702), .A2(new_n703), .ZN(new_n727));
  AOI211_X1 g302(.A(new_n726), .B(new_n727), .C1(new_n706), .C2(new_n710), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n721), .B(new_n728), .C1(new_n718), .C2(new_n717), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n720), .A2(G1341), .ZN(new_n730));
  INV_X1    g305(.A(G16), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G21), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G168), .B2(new_n731), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G1966), .ZN(new_n734));
  NOR3_X1   g309(.A1(new_n729), .A2(new_n730), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n731), .A2(G20), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT98), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT23), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n592), .B2(new_n731), .ZN(new_n739));
  INV_X1    g314(.A(G1956), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n731), .A2(G5), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G171), .B2(new_n731), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(G1961), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n595), .A2(G16), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G4), .B2(G16), .ZN(new_n746));
  INV_X1    g321(.A(G1348), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n746), .A2(new_n747), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT92), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n688), .A2(G26), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n751), .B(new_n752), .Z(new_n753));
  AOI22_X1  g328(.A1(G128), .A2(new_n480), .B1(new_n481), .B2(G140), .ZN(new_n754));
  OAI221_X1 g329(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n469), .C2(G116), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G29), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2067), .ZN(new_n759));
  NOR2_X1   g334(.A1(G27), .A2(G29), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G164), .B2(G29), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G2078), .ZN(new_n762));
  NOR4_X1   g337(.A1(new_n748), .A2(new_n749), .A3(new_n759), .A4(new_n762), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n735), .A2(new_n741), .A3(new_n744), .A4(new_n763), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n714), .A2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT36), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n731), .B1(new_n566), .B2(new_n572), .ZN(new_n767));
  NOR2_X1   g342(.A1(G6), .A2(G16), .ZN(new_n768));
  OR3_X1    g343(.A1(new_n767), .A2(KEYINPUT88), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(KEYINPUT88), .B1(new_n767), .B2(new_n768), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT32), .B(G1981), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n769), .A2(new_n772), .A3(new_n770), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n731), .A2(G23), .ZN(new_n776));
  INV_X1    g351(.A(G288), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(new_n731), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT33), .B(G1976), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(G166), .A2(new_n731), .ZN(new_n781));
  INV_X1    g356(.A(G1971), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n731), .A2(G22), .ZN(new_n783));
  OR3_X1    g358(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n782), .B1(new_n781), .B2(new_n783), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n780), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n774), .A2(new_n775), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(KEYINPUT89), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT89), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n774), .A2(new_n789), .A3(new_n786), .A4(new_n775), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n788), .A2(KEYINPUT34), .A3(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT90), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(KEYINPUT34), .B1(new_n788), .B2(new_n790), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n688), .A2(G25), .ZN(new_n795));
  OAI221_X1 g370(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n469), .C2(G107), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT86), .ZN(new_n797));
  AOI22_X1  g372(.A1(G119), .A2(new_n480), .B1(new_n481), .B2(G131), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n795), .B1(new_n800), .B2(new_n688), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT35), .B(G1991), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n803), .A2(KEYINPUT87), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n803), .A2(KEYINPUT87), .ZN(new_n805));
  MUX2_X1   g380(.A(G24), .B(G290), .S(G16), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G1986), .ZN(new_n807));
  NOR4_X1   g382(.A1(new_n794), .A2(new_n804), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n766), .B1(new_n793), .B2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n793), .A2(new_n808), .A3(new_n766), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n765), .B1(new_n810), .B2(new_n811), .ZN(G311));
  NOR2_X1   g387(.A1(new_n714), .A2(new_n764), .ZN(new_n813));
  INV_X1    g388(.A(new_n811), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(new_n809), .ZN(G150));
  NAND2_X1  g390(.A1(new_n595), .A2(G559), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT38), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n513), .A2(G93), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n511), .A2(G55), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n522), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n818), .B(new_n819), .C1(new_n531), .C2(new_n820), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(new_n539), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n539), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n817), .B(new_n824), .ZN(new_n825));
  AND2_X1   g400(.A1(new_n825), .A2(KEYINPUT39), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n825), .A2(KEYINPUT39), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n826), .A2(new_n827), .A3(G860), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n821), .A2(G860), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT99), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT37), .Z(new_n831));
  OR2_X1    g406(.A1(new_n828), .A2(new_n831), .ZN(G145));
  INV_X1    g407(.A(G37), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n611), .B(new_n478), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(G162), .ZN(new_n835));
  INV_X1    g410(.A(new_n701), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n686), .B(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n493), .ZN(new_n838));
  INV_X1    g413(.A(G138), .ZN(new_n839));
  OR2_X1    g414(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n840));
  NAND2_X1  g415(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n497), .B1(new_n842), .B2(new_n469), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n494), .A2(new_n476), .A3(KEYINPUT4), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n838), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n756), .B(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n837), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n799), .B(new_n604), .ZN(new_n848));
  AOI22_X1  g423(.A1(G130), .A2(new_n480), .B1(new_n481), .B2(G142), .ZN(new_n849));
  OAI221_X1 g424(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n469), .C2(G118), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n848), .B(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT100), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n837), .A2(new_n846), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n847), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n847), .A2(new_n855), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n852), .B(new_n853), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT101), .ZN(new_n860));
  AND3_X1   g435(.A1(new_n859), .A2(new_n860), .A3(new_n835), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n860), .B1(new_n859), .B2(new_n835), .ZN(new_n862));
  OAI221_X1 g437(.A(new_n833), .B1(new_n835), .B2(new_n859), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g439(.A(G305), .B(KEYINPUT104), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n865), .A2(G303), .ZN(new_n866));
  XNOR2_X1  g441(.A(G290), .B(G288), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(G303), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n867), .B1(new_n866), .B2(new_n868), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT42), .ZN(new_n872));
  NOR3_X1   g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n871), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n869), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(new_n872), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n599), .B(new_n824), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n595), .A2(G299), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n592), .A2(new_n586), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT41), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT103), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n881), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n879), .B(new_n883), .C1(new_n886), .C2(KEYINPUT41), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n878), .A2(new_n882), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n888), .A2(KEYINPUT102), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(KEYINPUT102), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n887), .A2(new_n889), .A3(KEYINPUT105), .A4(new_n890), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n874), .A2(new_n877), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(KEYINPUT42), .B1(new_n875), .B2(new_n869), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n892), .B(new_n891), .C1(new_n896), .C2(new_n873), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n897), .A3(G868), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n899), .B1(new_n821), .B2(new_n587), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n898), .A2(KEYINPUT106), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(G295));
  NOR2_X1   g478(.A1(new_n901), .A2(new_n902), .ZN(G331));
  NAND2_X1  g479(.A1(G171), .A2(G168), .ZN(new_n905));
  NAND2_X1  g480(.A1(G301), .A2(G286), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n907), .A2(new_n824), .ZN(new_n908));
  INV_X1    g483(.A(new_n824), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n909), .B1(new_n905), .B2(new_n906), .ZN(new_n910));
  OAI221_X1 g485(.A(new_n883), .B1(new_n908), .B2(new_n910), .C1(new_n886), .C2(KEYINPUT41), .ZN(new_n911));
  INV_X1    g486(.A(new_n882), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n910), .A2(KEYINPUT107), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n910), .A2(KEYINPUT107), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n911), .A2(KEYINPUT108), .A3(new_n916), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(new_n876), .A3(new_n920), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n911), .A2(new_n916), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n870), .A2(new_n871), .ZN(new_n923));
  AOI21_X1  g498(.A(G37), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT43), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n914), .B(new_n915), .C1(new_n824), .C2(new_n907), .ZN(new_n926));
  XOR2_X1   g501(.A(new_n885), .B(new_n881), .Z(new_n927));
  INV_X1    g502(.A(KEYINPUT109), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(new_n928), .A3(KEYINPUT41), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n927), .A2(KEYINPUT41), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT109), .B1(new_n912), .B2(KEYINPUT41), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n926), .B(new_n929), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  OR3_X1    g507(.A1(new_n908), .A2(new_n912), .A3(new_n910), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n923), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n833), .B1(new_n917), .B2(new_n876), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT44), .B1(new_n925), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n936), .B1(new_n921), .B2(new_n924), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n934), .A2(new_n935), .A3(KEYINPUT43), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n938), .A2(new_n942), .ZN(G397));
  INV_X1    g518(.A(KEYINPUT125), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT45), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(G164), .B2(G1384), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n472), .A2(G40), .A3(new_n477), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n800), .A2(new_n802), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n800), .A2(new_n802), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n948), .A2(G1996), .A3(new_n701), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  OR2_X1    g528(.A1(new_n953), .A2(KEYINPUT111), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(KEYINPUT111), .ZN(new_n955));
  INV_X1    g530(.A(G2067), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n756), .B(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(G1996), .B2(new_n701), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n954), .A2(new_n955), .B1(new_n948), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(G290), .A2(G1986), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(KEYINPUT110), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n961), .B1(G1986), .B2(G290), .ZN(new_n962));
  INV_X1    g537(.A(new_n948), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n951), .B(new_n959), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(G286), .A2(G8), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT122), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n967));
  INV_X1    g542(.A(G1384), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n845), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n969), .A2(new_n970), .A3(KEYINPUT113), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n845), .A2(new_n968), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT113), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(new_n973), .A3(KEYINPUT50), .ZN(new_n974));
  AOI211_X1 g549(.A(G2084), .B(new_n947), .C1(new_n971), .C2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n947), .B1(new_n972), .B2(new_n945), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n845), .A2(KEYINPUT45), .A3(new_n968), .ZN(new_n977));
  AOI21_X1  g552(.A(G1966), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n966), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n947), .B1(new_n971), .B2(new_n974), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n706), .ZN(new_n981));
  INV_X1    g556(.A(new_n978), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n981), .A2(new_n982), .A3(KEYINPUT122), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n965), .B1(new_n979), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n979), .A2(new_n983), .A3(G168), .ZN(new_n985));
  AND2_X1   g560(.A1(KEYINPUT51), .A2(G8), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n981), .A2(new_n982), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(G8), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT51), .B1(G286), .B2(G8), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n984), .B1(new_n987), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT54), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n977), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G2078), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n845), .A2(KEYINPUT112), .A3(KEYINPUT45), .A4(new_n968), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n976), .A2(new_n995), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n947), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n997), .A2(new_n1001), .A3(new_n946), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n1002), .A2(KEYINPUT53), .A3(new_n996), .A4(new_n995), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n1000), .B(new_n1003), .C1(G1961), .C2(new_n980), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n993), .B1(new_n1004), .B2(G171), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n976), .A2(KEYINPUT53), .A3(new_n996), .A4(new_n977), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1006), .B1(new_n980), .B2(G1961), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT123), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g584(.A(KEYINPUT123), .B(new_n1006), .C1(new_n980), .C2(G1961), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1009), .A2(G301), .A3(new_n1000), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1005), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n971), .A2(new_n974), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n947), .A2(G2090), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n976), .A2(new_n995), .A3(new_n997), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n782), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1015), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1013), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1021), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1023), .A2(KEYINPUT115), .A3(new_n1019), .A4(new_n1017), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n1025));
  INV_X1    g600(.A(G8), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1025), .B1(G166), .B2(new_n1026), .ZN(new_n1027));
  OAI211_X1 g602(.A(KEYINPUT55), .B(G8), .C1(new_n506), .C2(new_n516), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1022), .A2(new_n1024), .A3(G8), .A4(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1981), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n564), .A2(new_n565), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(G1981), .B1(new_n570), .B2(new_n571), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT49), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1034), .A2(KEYINPUT118), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n495), .A2(new_n498), .ZN(new_n1037));
  AOI21_X1  g612(.A(G1384), .B1(new_n1037), .B2(new_n838), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1026), .B1(new_n1001), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT118), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1032), .B(new_n1033), .C1(new_n1040), .C2(KEYINPUT49), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1036), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n557), .A2(G1976), .A3(new_n558), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT116), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n557), .A2(new_n1046), .A3(G1976), .A4(new_n558), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1039), .A2(new_n1044), .A3(new_n1045), .A4(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G1976), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1039), .A2(new_n1046), .A3(new_n1049), .A4(G288), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n1048), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1048), .B1(new_n1051), .B2(new_n1050), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1042), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n969), .A2(new_n1001), .A3(new_n970), .ZN(new_n1055));
  OR2_X1    g630(.A1(new_n1055), .A2(G2090), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1019), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1029), .B1(new_n1057), .B2(G8), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1054), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1012), .A2(new_n1030), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT124), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n997), .A2(new_n1001), .A3(new_n946), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT112), .B1(new_n1038), .B2(KEYINPUT45), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n1062), .A2(G2078), .A3(new_n1063), .ZN(new_n1064));
  OAI22_X1  g639(.A1(new_n1064), .A2(KEYINPUT53), .B1(new_n980), .B2(G1961), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1003), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1065), .A2(new_n1066), .A3(G171), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1009), .A2(new_n1000), .A3(new_n1010), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1067), .B1(G171), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1061), .B1(new_n1069), .B2(KEYINPUT54), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n1010), .A2(new_n1000), .ZN(new_n1071));
  AOI21_X1  g646(.A(G301), .B1(new_n1071), .B2(new_n1009), .ZN(new_n1072));
  OAI211_X1 g647(.A(KEYINPUT124), .B(new_n993), .C1(new_n1072), .C2(new_n1067), .ZN(new_n1073));
  AOI211_X1 g648(.A(new_n992), .B(new_n1060), .C1(new_n1070), .C2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1018), .A2(G1996), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n972), .A2(new_n947), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT58), .B(G1341), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n540), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g654(.A(new_n1079), .B(KEYINPUT59), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT56), .B(G2072), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1002), .A2(new_n995), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1055), .A2(new_n740), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n547), .A2(new_n1087), .A3(new_n551), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1085), .A2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1083), .A2(new_n1086), .A3(new_n1088), .A4(new_n1084), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1081), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1092), .A2(KEYINPUT61), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1092), .A2(KEYINPUT61), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1080), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1076), .A2(new_n956), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n980), .B2(G1348), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT119), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g674(.A(KEYINPUT119), .B(new_n1096), .C1(new_n980), .C2(G1348), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT60), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n586), .B1(new_n1102), .B2(KEYINPUT121), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT60), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1104), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT121), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1105), .A2(new_n1106), .A3(new_n595), .ZN(new_n1107));
  OAI22_X1  g682(.A1(new_n1103), .A2(new_n1107), .B1(KEYINPUT121), .B2(new_n1102), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1099), .A2(new_n1104), .A3(new_n1100), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1095), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1099), .A2(new_n595), .A3(new_n1100), .A4(new_n1091), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n1090), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1074), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT63), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1030), .A2(new_n1059), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n988), .A2(G8), .A3(G168), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1114), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1022), .A2(new_n1024), .A3(G8), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1118), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1054), .A2(new_n1116), .A3(new_n1114), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1119), .A2(new_n1030), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n992), .A2(new_n1123), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1030), .A2(new_n1059), .A3(new_n1072), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n985), .A2(new_n986), .B1(new_n989), .B2(new_n990), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT62), .B1(new_n1126), .B2(new_n984), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1124), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1030), .A2(new_n1054), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1042), .A2(new_n1049), .A3(new_n777), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n1032), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1129), .B1(new_n1039), .B2(new_n1131), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1122), .A2(new_n1128), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n964), .B1(new_n1113), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n963), .A2(G1996), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1135), .B(KEYINPUT46), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n963), .B1(new_n836), .B2(new_n957), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  XOR2_X1   g713(.A(new_n1138), .B(KEYINPUT47), .Z(new_n1139));
  NAND2_X1  g714(.A1(new_n961), .A2(new_n948), .ZN(new_n1140));
  XOR2_X1   g715(.A(new_n1140), .B(KEYINPUT48), .Z(new_n1141));
  NAND2_X1  g716(.A1(new_n959), .A2(new_n951), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1139), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n756), .A2(G2067), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1144), .B1(new_n959), .B2(new_n949), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1145), .A2(new_n963), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n944), .B1(new_n1134), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1122), .A2(new_n1128), .A3(new_n1132), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1112), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1102), .A2(KEYINPUT121), .A3(new_n586), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n595), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n1152), .A2(new_n1153), .B1(new_n1106), .B2(new_n1105), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1109), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1151), .B1(new_n1156), .B2(new_n1095), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1150), .B1(new_n1157), .B2(new_n1074), .ZN(new_n1158));
  OAI211_X1 g733(.A(KEYINPUT125), .B(new_n1147), .C1(new_n1158), .C2(new_n964), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1149), .A2(new_n1159), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g735(.A1(new_n940), .A2(new_n941), .ZN(new_n1162));
  NOR2_X1   g736(.A1(G227), .A2(new_n460), .ZN(new_n1163));
  NAND2_X1  g737(.A1(new_n678), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g738(.A1(new_n1164), .A2(G401), .ZN(new_n1165));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n1166));
  NOR2_X1   g740(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NOR3_X1   g741(.A1(new_n1164), .A2(G401), .A3(KEYINPUT126), .ZN(new_n1168));
  OAI21_X1  g742(.A(new_n863), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g743(.A1(new_n1162), .A2(new_n1169), .ZN(G308));
  OAI221_X1 g744(.A(new_n863), .B1(new_n1167), .B2(new_n1168), .C1(new_n940), .C2(new_n941), .ZN(G225));
endmodule


