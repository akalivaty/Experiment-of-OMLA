//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 0 1 1 1 0 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1265, new_n1266, new_n1267, new_n1268;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  NOR2_X1   g0006(.A1(G97), .A2(G107), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G107), .ZN(new_n210));
  INV_X1    g0010(.A(G264), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G116), .A2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G87), .ZN(new_n215));
  INV_X1    g0015(.A(G250), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n213), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n212), .B(new_n217), .C1(G50), .C2(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G58), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G20), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT1), .Z(new_n226));
  NOR2_X1   g0026(.A1(new_n224), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(G257), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n216), .B(new_n228), .C1(new_n229), .C2(new_n211), .ZN(new_n230));
  OR2_X1    g0030(.A1(new_n230), .A2(KEYINPUT0), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n230), .A2(KEYINPUT0), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n234), .A2(G20), .ZN(new_n235));
  INV_X1    g0035(.A(new_n201), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n236), .A2(G50), .ZN(new_n237));
  OAI211_X1 g0037(.A(new_n231), .B(new_n232), .C1(new_n235), .C2(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT65), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n226), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT66), .ZN(G361));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G232), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT2), .B(G226), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G250), .B(G257), .Z(new_n246));
  XNOR2_X1  g0046(.A(G264), .B(G270), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G358));
  XOR2_X1   g0049(.A(G68), .B(G77), .Z(new_n250));
  XOR2_X1   g0050(.A(G50), .B(G58), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(G87), .B(G97), .Z(new_n253));
  XNOR2_X1  g0053(.A(G107), .B(G116), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XOR2_X1   g0055(.A(new_n252), .B(new_n255), .Z(G351));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  OAI21_X1  g0057(.A(KEYINPUT68), .B1(new_n224), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT68), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n259), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n258), .A2(new_n233), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G20), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n204), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT8), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n219), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT69), .B(G58), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n265), .B1(new_n266), .B2(new_n264), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n262), .A2(G33), .ZN(new_n268));
  INV_X1    g0068(.A(G150), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n262), .A2(new_n257), .ZN(new_n270));
  OAI22_X1  g0070(.A1(new_n267), .A2(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n261), .B1(new_n263), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G1), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G20), .ZN(new_n274));
  INV_X1    g0074(.A(G13), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n202), .ZN(new_n277));
  AND3_X1   g0077(.A1(new_n258), .A2(new_n233), .A3(new_n260), .ZN(new_n278));
  INV_X1    g0078(.A(new_n276), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n278), .A2(KEYINPUT70), .A3(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT70), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n281), .B1(new_n261), .B2(new_n276), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n280), .A2(new_n274), .A3(new_n282), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n272), .B(new_n277), .C1(new_n283), .C2(new_n202), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT9), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n284), .B1(KEYINPUT72), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(KEYINPUT72), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n286), .B(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT3), .B(G33), .ZN(new_n290));
  INV_X1    g0090(.A(G1698), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(G222), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT67), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT3), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G77), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n290), .A2(G223), .A3(G1698), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT67), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n290), .A2(new_n300), .A3(G222), .A4(new_n291), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n293), .A2(new_n298), .A3(new_n299), .A4(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G41), .ZN(new_n305));
  OAI211_X1 g0105(.A(G1), .B(G13), .C1(new_n257), .C2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n273), .B1(G41), .B2(G45), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G226), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n273), .B(G274), .C1(G41), .C2(G45), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n304), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(KEYINPUT73), .B1(new_n313), .B2(G190), .ZN(new_n314));
  INV_X1    g0114(.A(G200), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT73), .ZN(new_n317));
  INV_X1    g0117(.A(G190), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n312), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n314), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n289), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT10), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT10), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n289), .A2(new_n323), .A3(new_n320), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G179), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n313), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n327), .B(new_n284), .C1(G169), .C2(new_n313), .ZN(new_n328));
  NOR2_X1   g0128(.A1(G226), .A2(G1698), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(new_n220), .B2(G1698), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n330), .A2(new_n290), .B1(G33), .B2(G97), .ZN(new_n331));
  OAI221_X1 g0131(.A(new_n311), .B1(new_n222), .B2(new_n308), .C1(new_n331), .C2(new_n306), .ZN(new_n332));
  OR2_X1    g0132(.A1(new_n332), .A2(KEYINPUT13), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT74), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(KEYINPUT13), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n332), .A2(KEYINPUT74), .A3(KEYINPUT13), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(G169), .A3(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(KEYINPUT75), .B2(KEYINPUT14), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n333), .A2(new_n335), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n340), .A2(G179), .B1(KEYINPUT75), .B2(KEYINPUT14), .ZN(new_n341));
  NOR2_X1   g0141(.A1(KEYINPUT75), .A2(KEYINPUT14), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n336), .A2(G169), .A3(new_n342), .A4(new_n337), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n339), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n270), .A2(new_n202), .B1(new_n262), .B2(G68), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n268), .A2(new_n205), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n261), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n347), .B(KEYINPUT11), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n276), .A2(new_n221), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n349), .B(KEYINPUT12), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n278), .A2(new_n274), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n348), .B(new_n350), .C1(new_n221), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n344), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n340), .A2(G190), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n336), .A2(G200), .A3(new_n337), .ZN(new_n355));
  INV_X1    g0155(.A(new_n352), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n325), .A2(new_n328), .A3(new_n353), .A4(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n294), .A2(KEYINPUT76), .A3(G33), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT76), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(KEYINPUT3), .B2(new_n257), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n359), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT77), .B(KEYINPUT7), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n262), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT7), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT76), .B1(new_n294), .B2(G33), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n295), .ZN(new_n369));
  AOI21_X1  g0169(.A(G20), .B1(new_n369), .B2(new_n359), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n366), .B(G68), .C1(new_n367), .C2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G159), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n270), .A2(new_n372), .ZN(new_n373));
  XOR2_X1   g0173(.A(KEYINPUT69), .B(G58), .Z(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G68), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n236), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n373), .B1(new_n376), .B2(G20), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n371), .A2(new_n377), .A3(KEYINPUT16), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT16), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n201), .B1(new_n374), .B2(G68), .ZN(new_n380));
  OAI22_X1  g0180(.A1(new_n380), .A2(new_n262), .B1(new_n372), .B2(new_n270), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n365), .B1(G20), .B2(new_n290), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n297), .A2(KEYINPUT7), .A3(new_n262), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n221), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n379), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n378), .A2(new_n385), .A3(new_n261), .ZN(new_n386));
  MUX2_X1   g0186(.A(new_n283), .B(new_n279), .S(new_n267), .Z(new_n387));
  OR2_X1    g0187(.A1(G223), .A2(G1698), .ZN(new_n388));
  OR2_X1    g0188(.A1(new_n291), .A2(G226), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n369), .A2(new_n359), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G33), .A2(G87), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n303), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n309), .A2(G232), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n393), .A2(new_n318), .A3(new_n311), .A4(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n311), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n306), .B1(new_n390), .B2(new_n391), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n315), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n386), .A2(new_n387), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT78), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT78), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n386), .A2(new_n387), .A3(new_n399), .A4(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT79), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n405), .A3(KEYINPUT17), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n386), .A2(new_n387), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n396), .A2(new_n397), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(G179), .ZN(new_n409));
  INV_X1    g0209(.A(G169), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n409), .B1(new_n410), .B2(new_n408), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT18), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n407), .A2(KEYINPUT18), .A3(new_n411), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT17), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(new_n401), .B2(new_n403), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT79), .B1(new_n400), .B2(KEYINPUT17), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n406), .B(new_n416), .C1(new_n418), .C2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n290), .A2(G232), .A3(new_n291), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n290), .A2(G238), .A3(G1698), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n421), .B(new_n422), .C1(new_n210), .C2(new_n290), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n303), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n309), .A2(G244), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n424), .A2(new_n311), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(G190), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G20), .A2(G77), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT15), .B(G87), .ZN(new_n429));
  XNOR2_X1  g0229(.A(KEYINPUT8), .B(G58), .ZN(new_n430));
  OAI221_X1 g0230(.A(new_n428), .B1(new_n429), .B2(new_n268), .C1(new_n270), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n261), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n276), .A2(new_n205), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n278), .A2(G77), .A3(new_n274), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n427), .B(new_n436), .C1(new_n315), .C2(new_n426), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n426), .A2(new_n326), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n438), .B(new_n435), .C1(G169), .C2(new_n426), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n440), .B(KEYINPUT71), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n358), .A2(new_n420), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT22), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n443), .A2(new_n215), .A3(G20), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n444), .B(new_n359), .C1(new_n361), .C2(new_n362), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n215), .A2(G20), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n446), .A2(new_n295), .A3(new_n296), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n443), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G33), .A2(G116), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n262), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT23), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n262), .B2(G107), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n210), .A2(KEYINPUT23), .A3(G20), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n445), .A2(new_n448), .A3(new_n451), .A4(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT24), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n447), .A2(new_n443), .B1(new_n453), .B2(new_n454), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n459), .A2(KEYINPUT24), .A3(new_n445), .A4(new_n451), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n458), .A2(new_n261), .A3(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n257), .A2(G1), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n261), .A2(new_n276), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G107), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n216), .A2(new_n291), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n229), .A2(G1698), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n369), .A2(new_n359), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G294), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n303), .ZN(new_n471));
  INV_X1    g0271(.A(G45), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(G1), .ZN(new_n473));
  AND2_X1   g0273(.A1(KEYINPUT5), .A2(G41), .ZN(new_n474));
  NOR2_X1   g0274(.A1(KEYINPUT5), .A2(G41), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n476), .A2(G264), .A3(new_n306), .ZN(new_n477));
  XNOR2_X1  g0277(.A(KEYINPUT5), .B(G41), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n478), .A2(G274), .A3(new_n473), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n471), .A2(new_n318), .A3(new_n477), .A4(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n306), .B1(new_n468), .B2(new_n469), .ZN(new_n481));
  INV_X1    g0281(.A(new_n477), .ZN(new_n482));
  INV_X1    g0282(.A(new_n479), .ZN(new_n483));
  NOR3_X1   g0283(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n480), .B1(new_n484), .B2(G200), .ZN(new_n485));
  OAI211_X1 g0285(.A(KEYINPUT86), .B(KEYINPUT25), .C1(new_n279), .C2(G107), .ZN(new_n486));
  NAND2_X1  g0286(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n487));
  OR2_X1    g0287(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n276), .A2(new_n210), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n465), .A2(new_n485), .A3(new_n486), .A4(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n364), .B1(new_n262), .B2(new_n297), .ZN(new_n491));
  NOR3_X1   g0291(.A1(new_n290), .A2(new_n367), .A3(G20), .ZN(new_n492));
  OAI21_X1  g0292(.A(G107), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n210), .A2(KEYINPUT6), .A3(G97), .ZN(new_n494));
  INV_X1    g0294(.A(G97), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(new_n210), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(new_n207), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n494), .B1(new_n497), .B2(KEYINPUT6), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G20), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT80), .B1(new_n270), .B2(new_n205), .ZN(new_n500));
  OR3_X1    g0300(.A1(new_n270), .A2(KEYINPUT80), .A3(new_n205), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n493), .A2(new_n499), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n261), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n279), .A2(G97), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n504), .B1(new_n463), .B2(G97), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n291), .A2(G244), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n359), .B(new_n508), .C1(new_n361), .C2(new_n362), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT4), .ZN(new_n510));
  OAI22_X1  g0310(.A1(new_n507), .A2(new_n510), .B1(new_n216), .B2(new_n291), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n509), .A2(new_n510), .B1(new_n290), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G283), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n306), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n476), .A2(G257), .A3(new_n306), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n479), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n410), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n509), .A2(new_n510), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n511), .A2(new_n290), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(new_n513), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n303), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT81), .B1(new_n515), .B2(new_n479), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n515), .A2(KEYINPUT81), .A3(new_n479), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n521), .B(new_n326), .C1(new_n522), .C2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n506), .A2(new_n517), .A3(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n524), .A2(new_n522), .ZN(new_n527));
  OAI21_X1  g0327(.A(G200), .B1(new_n527), .B2(new_n514), .ZN(new_n528));
  INV_X1    g0328(.A(new_n516), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n521), .A2(G190), .A3(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n528), .A2(new_n503), .A3(new_n530), .A4(new_n505), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n476), .A2(G270), .A3(new_n306), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT85), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n476), .A2(KEYINPUT85), .A3(G270), .A4(new_n306), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n483), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n229), .A2(new_n291), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n211), .A2(G1698), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n369), .A2(new_n359), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n297), .A2(G303), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n303), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G200), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n279), .A2(G116), .ZN(new_n545));
  INV_X1    g0345(.A(G116), .ZN(new_n546));
  NOR4_X1   g0346(.A1(new_n261), .A2(new_n546), .A3(new_n276), .A4(new_n462), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(G20), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n513), .B(new_n262), .C1(G33), .C2(new_n495), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n261), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT20), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n261), .A2(KEYINPUT20), .A3(new_n548), .A4(new_n549), .ZN(new_n553));
  AOI211_X1 g0353(.A(new_n545), .B(new_n547), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n544), .B(new_n554), .C1(new_n318), .C2(new_n543), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n490), .A2(new_n526), .A3(new_n531), .A4(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n461), .A2(new_n486), .A3(new_n464), .A4(new_n489), .ZN(new_n557));
  INV_X1    g0357(.A(new_n484), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n410), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n484), .A2(new_n326), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n557), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT21), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n543), .A2(G169), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n562), .B1(new_n563), .B2(new_n554), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n547), .B1(new_n552), .B2(new_n553), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(G116), .B2(new_n279), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n566), .A2(KEYINPUT21), .A3(G169), .A4(new_n543), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n534), .A2(new_n535), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n542), .A2(new_n568), .A3(G179), .A4(new_n479), .ZN(new_n569));
  OR2_X1    g0369(.A1(new_n554), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n561), .A2(new_n564), .A3(new_n567), .A4(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n556), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT84), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT82), .ZN(new_n574));
  NOR2_X1   g0374(.A1(G238), .A2(G1698), .ZN(new_n575));
  INV_X1    g0375(.A(G244), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n575), .B1(new_n576), .B2(G1698), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n369), .A2(new_n577), .A3(new_n359), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n306), .B1(new_n578), .B2(new_n449), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n473), .A2(G274), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n306), .B1(G1), .B2(new_n472), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n580), .B1(new_n581), .B2(new_n216), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n574), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n303), .A2(new_n473), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n584), .A2(G250), .B1(G274), .B2(new_n473), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n294), .A2(KEYINPUT76), .A3(G33), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n586), .B1(new_n295), .B2(new_n368), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n450), .B1(new_n587), .B2(new_n577), .ZN(new_n588));
  OAI211_X1 g0388(.A(KEYINPUT82), .B(new_n585), .C1(new_n588), .C2(new_n306), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n583), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G200), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n583), .A2(new_n589), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G190), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n369), .A2(new_n262), .A3(G68), .A4(new_n359), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT19), .ZN(new_n595));
  NOR3_X1   g0395(.A1(new_n595), .A2(new_n257), .A3(new_n495), .ZN(new_n596));
  OAI22_X1  g0396(.A1(new_n596), .A2(G20), .B1(G87), .B2(new_n208), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n595), .B1(new_n268), .B2(new_n495), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n594), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n599), .A2(new_n261), .B1(new_n276), .B2(new_n429), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n463), .A2(G87), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n591), .A2(new_n593), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT83), .B1(new_n592), .B2(new_n326), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n592), .A2(KEYINPUT83), .A3(new_n326), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n583), .A2(new_n589), .A3(new_n410), .ZN(new_n608));
  INV_X1    g0408(.A(new_n429), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n463), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n600), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n573), .B(new_n603), .C1(new_n607), .C2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT83), .ZN(new_n614));
  AOI211_X1 g0414(.A(new_n614), .B(G179), .C1(new_n583), .C2(new_n589), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n604), .A2(new_n615), .A3(new_n612), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n591), .A2(new_n593), .A3(new_n602), .ZN(new_n617));
  OAI21_X1  g0417(.A(KEYINPUT84), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n572), .A2(new_n613), .A3(new_n618), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n442), .A2(new_n619), .ZN(G372));
  AND3_X1   g0420(.A1(new_n506), .A2(new_n517), .A3(new_n525), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n618), .A2(new_n613), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT26), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n579), .A2(new_n582), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n593), .B(new_n602), .C1(new_n315), .C2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n592), .A2(new_n326), .ZN(new_n628));
  INV_X1    g0428(.A(new_n626), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n410), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n628), .A2(new_n611), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n621), .A2(new_n627), .A3(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n632), .A2(KEYINPUT26), .ZN(new_n633));
  INV_X1    g0433(.A(new_n631), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT87), .ZN(new_n636));
  XNOR2_X1  g0436(.A(new_n571), .B(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n627), .A2(new_n631), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n526), .A2(new_n531), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(new_n490), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n635), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n625), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n442), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n328), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n419), .B1(new_n404), .B2(KEYINPUT17), .ZN(new_n646));
  AOI211_X1 g0446(.A(KEYINPUT79), .B(new_n417), .C1(new_n401), .C2(new_n403), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n439), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n344), .A2(new_n352), .B1(new_n357), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n416), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n645), .B1(new_n652), .B2(new_n325), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n644), .A2(new_n653), .ZN(G369));
  NOR2_X1   g0454(.A1(new_n275), .A2(G20), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n273), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n657), .A2(G213), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G343), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT88), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n566), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT89), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n564), .A2(new_n567), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n570), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n664), .A2(new_n570), .A3(new_n555), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n666), .B1(new_n667), .B2(new_n663), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(G330), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n561), .A2(new_n661), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n661), .A2(new_n557), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n490), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n671), .B1(new_n561), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n661), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n674), .A2(new_n665), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n671), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n675), .A2(new_n680), .ZN(G399));
  NOR2_X1   g0481(.A1(new_n228), .A2(G41), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G1), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n207), .A2(new_n215), .A3(new_n546), .ZN(new_n685));
  OAI22_X1  g0485(.A1(new_n684), .A2(new_n685), .B1(new_n237), .B2(new_n683), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT28), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n622), .A2(new_n623), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n632), .A2(KEYINPUT26), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n631), .ZN(new_n690));
  INV_X1    g0490(.A(new_n640), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n690), .B1(new_n691), .B2(new_n571), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n661), .B1(new_n688), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT29), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n661), .B1(new_n625), .B2(new_n642), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n694), .B1(new_n695), .B2(KEYINPUT29), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT90), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n527), .A2(new_n514), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n697), .B1(new_n698), .B2(new_n484), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n629), .A2(new_n543), .A3(new_n326), .ZN(new_n700));
  OAI211_X1 g0500(.A(new_n558), .B(KEYINPUT90), .C1(new_n514), .C2(new_n527), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n569), .B1(new_n583), .B2(new_n589), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n482), .B1(new_n470), .B2(new_n303), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n521), .A2(new_n705), .A3(new_n529), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n703), .B1(new_n704), .B2(new_n707), .ZN(new_n708));
  NOR4_X1   g0508(.A1(new_n590), .A2(new_n706), .A3(KEYINPUT30), .A4(new_n569), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n702), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(KEYINPUT91), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT91), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n702), .B(new_n712), .C1(new_n708), .C2(new_n709), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n711), .A2(new_n661), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT31), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n572), .A2(new_n618), .A3(new_n613), .A4(new_n676), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n710), .A2(KEYINPUT31), .A3(new_n661), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G330), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n696), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n687), .B1(new_n721), .B2(G1), .ZN(G364));
  AOI21_X1  g0522(.A(new_n684), .B1(G45), .B2(new_n655), .ZN(new_n723));
  XOR2_X1   g0523(.A(new_n723), .B(KEYINPUT92), .Z(new_n724));
  AOI21_X1  g0524(.A(new_n233), .B1(G20), .B2(new_n410), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(G303), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n262), .A2(new_n318), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n315), .A2(G179), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n728), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n731), .A2(new_n326), .A3(G200), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(G322), .ZN(new_n734));
  OAI221_X1 g0534(.A(new_n297), .B1(new_n727), .B2(new_n730), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n326), .A2(new_n315), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n262), .A2(G190), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  XNOR2_X1  g0539(.A(KEYINPUT33), .B(G317), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n735), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n736), .A2(new_n728), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G326), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n737), .A2(new_n729), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G179), .A2(G200), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n737), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI22_X1  g0549(.A1(G283), .A2(new_n746), .B1(new_n749), .B2(G329), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT96), .ZN(new_n751));
  INV_X1    g0551(.A(new_n737), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n752), .A2(new_n326), .A3(G200), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n262), .B1(new_n747), .B2(G190), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n753), .A2(G311), .B1(G294), .B2(new_n755), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n741), .A2(new_n744), .A3(new_n751), .A4(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n754), .A2(new_n495), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(G107), .B2(new_n746), .ZN(new_n759));
  INV_X1    g0559(.A(new_n730), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G87), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n753), .A2(G77), .ZN(new_n762));
  AND3_X1   g0562(.A1(new_n759), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n732), .A2(new_n374), .B1(new_n743), .B2(G50), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n297), .B1(new_n739), .B2(G68), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n748), .A2(new_n372), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT32), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n763), .A2(new_n764), .A3(new_n765), .A4(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n726), .B1(new_n757), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(G355), .A2(new_n290), .A3(new_n227), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(G116), .B2(new_n227), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT93), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n252), .A2(G45), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT94), .Z(new_n774));
  NOR2_X1   g0574(.A1(new_n587), .A2(new_n228), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(G45), .B2(new_n237), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n772), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G13), .A2(G33), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(G20), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n725), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT95), .Z(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n724), .B(new_n769), .C1(new_n777), .C2(new_n783), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT97), .Z(new_n785));
  INV_X1    g0585(.A(new_n780), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n785), .B1(new_n668), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n723), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n669), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n668), .A2(G330), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n787), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n791), .B(KEYINPUT98), .Z(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(G396));
  OAI211_X1 g0593(.A(new_n439), .B(new_n437), .C1(new_n436), .C2(new_n676), .ZN(new_n794));
  INV_X1    g0594(.A(KEYINPUT99), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n794), .B(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n797), .B(new_n676), .C1(new_n624), .C2(new_n641), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n650), .A2(new_n661), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n798), .B1(new_n695), .B2(new_n800), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n801), .A2(new_n720), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n720), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n802), .A2(new_n788), .A3(new_n803), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n796), .A2(new_n799), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n724), .B1(new_n805), .B2(new_n778), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n725), .A2(new_n778), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n205), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n730), .A2(new_n210), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n758), .B(new_n809), .C1(G116), .C2(new_n753), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n739), .A2(G283), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n290), .B1(new_n732), .B2(G294), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n742), .A2(new_n727), .B1(new_n745), .B2(new_n215), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(G311), .B2(new_n749), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n810), .A2(new_n811), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  AOI22_X1  g0615(.A1(G143), .A2(new_n732), .B1(new_n753), .B2(G159), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n743), .A2(G137), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n816), .B(new_n817), .C1(new_n269), .C2(new_n738), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT34), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n745), .A2(new_n221), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(G50), .B2(new_n760), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n363), .B1(G132), .B2(new_n749), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n819), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n754), .A2(new_n266), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n815), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n725), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n806), .A2(new_n808), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n804), .A2(new_n827), .ZN(G384));
  NAND4_X1  g0628(.A1(new_n711), .A2(KEYINPUT31), .A3(new_n661), .A4(new_n713), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n716), .A2(new_n717), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n442), .A2(new_n830), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n659), .B(KEYINPUT100), .Z(new_n832));
  NAND2_X1  g0632(.A1(new_n407), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n420), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(KEYINPUT37), .B1(new_n407), .B2(new_n832), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n404), .A2(new_n412), .A3(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n412), .A2(new_n833), .A3(new_n400), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(KEYINPUT37), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(KEYINPUT38), .B1(new_n835), .B2(new_n840), .ZN(new_n841));
  AND3_X1   g0641(.A1(new_n404), .A2(new_n412), .A3(new_n836), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT37), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n378), .A2(new_n261), .ZN(new_n844));
  AOI21_X1  g0644(.A(KEYINPUT16), .B1(new_n371), .B2(new_n377), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n387), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n411), .B2(new_n659), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n843), .B1(new_n404), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(KEYINPUT101), .B1(new_n842), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n404), .A2(new_n847), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(KEYINPUT37), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT101), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n851), .A2(new_n852), .A3(new_n837), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n846), .A2(new_n659), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n849), .A2(new_n853), .B1(new_n420), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n841), .B1(KEYINPUT38), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n661), .A2(new_n352), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n353), .A2(new_n357), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n344), .A2(new_n352), .A3(new_n661), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n830), .A2(new_n800), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT40), .B1(new_n856), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n849), .A2(new_n853), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n420), .A2(new_n854), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT38), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n863), .A2(KEYINPUT38), .A3(new_n864), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT40), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n830), .A2(new_n870), .A3(new_n800), .A4(new_n860), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n831), .B1(new_n862), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n861), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n833), .B1(new_n648), .B2(new_n416), .ZN(new_n876));
  INV_X1    g0676(.A(new_n840), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n866), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n868), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n870), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n871), .B1(new_n868), .B2(new_n867), .ZN(new_n881));
  OAI21_X1  g0681(.A(G330), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n442), .A2(G330), .A3(new_n830), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n874), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n884), .B(KEYINPUT102), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n442), .B(new_n694), .C1(new_n695), .C2(KEYINPUT29), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n653), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n885), .B(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n353), .A2(new_n661), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT39), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(new_n867), .B2(new_n868), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n878), .A2(new_n868), .A3(new_n890), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n416), .A2(new_n832), .ZN(new_n894));
  INV_X1    g0694(.A(new_n860), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n439), .A2(new_n661), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n895), .B1(new_n798), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n894), .B1(new_n869), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n893), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n888), .B(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n273), .B2(new_n655), .ZN(new_n902));
  OAI211_X1 g0702(.A(G20), .B(new_n234), .C1(new_n498), .C2(KEYINPUT35), .ZN(new_n903));
  AOI211_X1 g0703(.A(new_n546), .B(new_n903), .C1(KEYINPUT35), .C2(new_n498), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n904), .B(KEYINPUT36), .Z(new_n905));
  NAND4_X1  g0705(.A1(new_n375), .A2(G50), .A3(G77), .A4(new_n236), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(G50), .B2(new_n221), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n907), .A2(G1), .A3(new_n275), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n902), .A2(new_n905), .A3(new_n908), .ZN(G367));
  NOR2_X1   g0709(.A1(new_n730), .A2(new_n266), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n739), .A2(G159), .B1(new_n749), .B2(G137), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n743), .A2(G143), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n911), .B(new_n912), .C1(new_n205), .C2(new_n745), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n910), .B(new_n913), .C1(G50), .C2(new_n753), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n297), .B1(new_n755), .B2(G68), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n914), .B(new_n915), .C1(new_n269), .C2(new_n733), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n916), .B(KEYINPUT108), .Z(new_n917));
  AOI22_X1  g0717(.A1(new_n753), .A2(G283), .B1(G107), .B2(new_n755), .ZN(new_n918));
  XNOR2_X1  g0718(.A(KEYINPUT107), .B(G311), .ZN(new_n919));
  OAI221_X1 g0719(.A(new_n918), .B1(new_n495), .B2(new_n745), .C1(new_n742), .C2(new_n919), .ZN(new_n920));
  AOI211_X1 g0720(.A(new_n587), .B(new_n920), .C1(G294), .C2(new_n739), .ZN(new_n921));
  INV_X1    g0721(.A(G317), .ZN(new_n922));
  OAI221_X1 g0722(.A(new_n921), .B1(new_n727), .B2(new_n733), .C1(new_n922), .C2(new_n748), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n730), .A2(new_n546), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT46), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n917), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT47), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n725), .ZN(new_n928));
  INV_X1    g0728(.A(new_n724), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n676), .A2(new_n602), .ZN(new_n930));
  MUX2_X1   g0730(.A(new_n638), .B(new_n634), .S(new_n930), .Z(new_n931));
  OR2_X1    g0731(.A1(new_n931), .A2(new_n786), .ZN(new_n932));
  INV_X1    g0732(.A(new_n775), .ZN(new_n933));
  OAI221_X1 g0733(.A(new_n783), .B1(new_n227), .B2(new_n429), .C1(new_n248), .C2(new_n933), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n928), .A2(new_n929), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n273), .B1(new_n655), .B2(G45), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n661), .A2(new_n506), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n639), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n621), .A2(new_n661), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n680), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n942), .B(new_n943), .Z(new_n944));
  INV_X1    g0744(.A(KEYINPUT105), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n945), .B(KEYINPUT44), .C1(new_n680), .C2(new_n941), .ZN(new_n946));
  INV_X1    g0746(.A(new_n941), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(KEYINPUT44), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n945), .A2(KEYINPUT44), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n679), .A2(new_n947), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n944), .A2(new_n946), .A3(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n675), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n951), .B(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n665), .A2(new_n676), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(new_n674), .Z(new_n955));
  INV_X1    g0755(.A(KEYINPUT106), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n669), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n956), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n957), .B(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n721), .B1(new_n953), .B2(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n682), .B(KEYINPUT41), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n937), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(KEYINPUT42), .B1(new_n677), .B2(new_n939), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT42), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n679), .B1(new_n964), .B2(new_n671), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n963), .B1(new_n526), .B2(new_n661), .C1(new_n965), .C2(new_n939), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n931), .A2(KEYINPUT43), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n931), .A2(KEYINPUT43), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n966), .A2(new_n968), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n971), .A2(KEYINPUT103), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(KEYINPUT103), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n952), .A2(new_n941), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n935), .B1(new_n962), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT109), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OAI211_X1 g0779(.A(KEYINPUT109), .B(new_n935), .C1(new_n962), .C2(new_n976), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(G387));
  INV_X1    g0781(.A(new_n959), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n982), .A2(new_n721), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n721), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n983), .A2(new_n682), .A3(new_n984), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n742), .A2(new_n734), .B1(new_n738), .B2(new_n919), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT111), .Z(new_n987));
  INV_X1    g0787(.A(new_n753), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n987), .B1(new_n727), .B2(new_n988), .C1(new_n922), .C2(new_n733), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT48), .ZN(new_n990));
  INV_X1    g0790(.A(G283), .ZN(new_n991));
  INV_X1    g0791(.A(G294), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n990), .B1(new_n991), .B2(new_n754), .C1(new_n992), .C2(new_n730), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT49), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n587), .B1(new_n993), .B2(new_n994), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n746), .A2(G116), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n749), .A2(G326), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n995), .A2(new_n996), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n988), .A2(new_n221), .B1(new_n267), .B2(new_n738), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT110), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n205), .B2(new_n730), .C1(new_n372), .C2(new_n742), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n754), .A2(new_n429), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n495), .B2(new_n745), .C1(new_n733), .C2(new_n202), .ZN(new_n1005));
  NOR3_X1   g0805(.A1(new_n1002), .A2(new_n363), .A3(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n269), .B2(new_n748), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n726), .B1(new_n999), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n775), .B1(new_n245), .B2(new_n472), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n290), .A2(new_n685), .A3(new_n227), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AOI211_X1 g0811(.A(G45), .B(new_n685), .C1(G68), .C2(G77), .ZN(new_n1012));
  OAI21_X1  g0812(.A(KEYINPUT50), .B1(new_n430), .B2(G50), .ZN(new_n1013));
  OR3_X1    g0813(.A1(new_n430), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1011), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n228), .A2(new_n210), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n782), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n1008), .A2(new_n724), .A3(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n674), .B2(new_n786), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n985), .B(new_n1020), .C1(new_n936), .C2(new_n959), .ZN(G393));
  AOI21_X1  g0821(.A(new_n683), .B1(new_n953), .B2(new_n984), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n953), .B2(new_n984), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n953), .A2(new_n936), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n724), .B1(new_n947), .B2(new_n780), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n783), .B1(new_n495), .B2(new_n227), .C1(new_n255), .C2(new_n933), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n290), .B1(new_n749), .B2(G322), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n210), .B2(new_n745), .C1(new_n991), .C2(new_n730), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT112), .Z(new_n1029));
  AOI22_X1  g0829(.A1(new_n732), .A2(G311), .B1(new_n743), .B2(G317), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT52), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G294), .B2(new_n753), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n739), .A2(G303), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n755), .A2(G116), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1029), .A2(new_n1032), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n988), .A2(new_n430), .B1(new_n215), .B2(new_n745), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n363), .B(new_n1036), .C1(G143), .C2(new_n749), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n732), .A2(G159), .B1(new_n743), .B2(G150), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT51), .Z(new_n1039));
  NAND2_X1  g0839(.A1(new_n739), .A2(G50), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n760), .A2(G68), .B1(new_n755), .B2(G77), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1037), .A2(new_n1039), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n1035), .A2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1025), .B(new_n1026), .C1(new_n726), .C2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1023), .A2(new_n1024), .A3(new_n1044), .ZN(G390));
  NAND3_X1  g0845(.A1(new_n886), .A2(new_n653), .A3(new_n883), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n619), .A2(new_n676), .B1(new_n714), .B2(new_n715), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n805), .B1(new_n1047), .B2(new_n829), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT113), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1048), .A2(new_n1049), .A3(G330), .A4(new_n860), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n830), .A2(G330), .A3(new_n800), .A4(new_n860), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(KEYINPUT113), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n719), .A2(G330), .A3(new_n800), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n895), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1050), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n798), .A2(new_n897), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n830), .A2(new_n800), .ZN(new_n1058));
  INV_X1    g0858(.A(G330), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n895), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n896), .B1(new_n693), .B2(new_n797), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(new_n895), .C2(new_n1053), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1046), .B1(new_n1057), .B2(new_n1062), .ZN(new_n1063));
  AND3_X1   g0863(.A1(new_n863), .A2(KEYINPUT38), .A3(new_n864), .ZN(new_n1064));
  AOI21_X1  g0864(.A(KEYINPUT38), .B1(new_n863), .B2(new_n864), .ZN(new_n1065));
  OAI21_X1  g0865(.A(KEYINPUT39), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n878), .A2(new_n868), .A3(new_n890), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1066), .B(new_n1067), .C1(new_n889), .C2(new_n898), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n889), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1069), .B(new_n879), .C1(new_n1061), .C2(new_n895), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1053), .A2(new_n895), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1063), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n682), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(KEYINPUT114), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1063), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1078), .A2(KEYINPUT115), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT115), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT114), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1075), .A2(new_n1084), .A3(new_n682), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1077), .A2(new_n1080), .A3(new_n1083), .A4(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1066), .A2(new_n778), .A3(new_n1067), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n267), .A2(new_n807), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n732), .A2(G132), .B1(new_n743), .B2(G128), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT117), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n760), .A2(G150), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1090), .B1(KEYINPUT53), .B2(new_n1091), .C1(new_n372), .C2(new_n754), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n297), .B(new_n1092), .C1(KEYINPUT53), .C2(new_n1091), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n746), .A2(G50), .ZN(new_n1094));
  XOR2_X1   g0894(.A(KEYINPUT54), .B(G143), .Z(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT116), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n753), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n739), .A2(G137), .B1(new_n749), .B2(G125), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1093), .A2(new_n1094), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n988), .A2(new_n495), .B1(new_n210), .B2(new_n738), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT118), .ZN(new_n1101));
  OR2_X1    g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1102), .B(new_n1103), .C1(new_n991), .C2(new_n742), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT119), .Z(new_n1105));
  NOR2_X1   g0905(.A1(new_n1105), .A2(new_n290), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n749), .A2(G294), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n732), .A2(G116), .B1(G77), .B2(new_n755), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT120), .Z(new_n1109));
  NAND4_X1  g0909(.A1(new_n1106), .A2(new_n761), .A3(new_n1107), .A4(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1099), .B1(new_n1110), .B2(new_n820), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n725), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1087), .A2(new_n929), .A3(new_n1088), .A4(new_n1112), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1086), .B(new_n1113), .C1(new_n936), .C2(new_n1078), .ZN(G378));
  INV_X1    g0914(.A(new_n1046), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1075), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1059), .B1(new_n862), .B2(new_n873), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n900), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n882), .A2(new_n893), .A3(new_n899), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n325), .A2(new_n328), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n284), .A2(new_n659), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1120), .B(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1122), .B(new_n1123), .Z(new_n1124));
  NAND3_X1  g0924(.A1(new_n1118), .A2(new_n1119), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1124), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1116), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT57), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n683), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1116), .B(KEYINPUT57), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT123), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1124), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1136), .A2(new_n1125), .B1(new_n1115), .B2(new_n1075), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1137), .A2(KEYINPUT123), .A3(KEYINPUT57), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1130), .A2(new_n1133), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1124), .A2(new_n778), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n363), .A2(new_n305), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1141), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n742), .A2(new_n546), .B1(new_n754), .B2(new_n221), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT121), .Z(new_n1144));
  NOR2_X1   g0944(.A1(new_n730), .A2(new_n205), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n746), .A2(new_n374), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n988), .B2(new_n429), .ZN(new_n1147));
  NOR4_X1   g0947(.A1(new_n1144), .A2(new_n1145), .A3(new_n1141), .A4(new_n1147), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n1148), .B1(new_n495), .B2(new_n738), .C1(new_n991), .C2(new_n748), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G107), .B2(new_n732), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1142), .B1(new_n1150), .B2(KEYINPUT58), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT122), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n257), .B(new_n305), .C1(new_n745), .C2(new_n372), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(G124), .B2(new_n749), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1096), .A2(new_n760), .B1(G125), .B2(new_n743), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(G128), .A2(new_n732), .B1(new_n753), .B2(G137), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1155), .B(new_n1156), .C1(new_n269), .C2(new_n754), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(G132), .B2(new_n739), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT59), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1150), .A2(KEYINPUT58), .B1(new_n1154), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1152), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n725), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n807), .A2(new_n202), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1140), .A2(new_n723), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1136), .A2(new_n1125), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1165), .B1(new_n1166), .B2(new_n937), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1139), .A2(new_n1167), .ZN(G375));
  AND2_X1   g0968(.A1(new_n1057), .A2(new_n1062), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1169), .A2(new_n936), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1004), .B1(new_n495), .B2(new_n730), .C1(new_n727), .C2(new_n748), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n733), .A2(new_n991), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n988), .A2(new_n210), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n742), .A2(new_n992), .ZN(new_n1174));
  NOR4_X1   g0974(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n290), .B1(new_n746), .B2(G77), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1175), .B(new_n1176), .C1(new_n546), .C2(new_n738), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT124), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n749), .A2(G128), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1146), .B(new_n1179), .C1(new_n372), .C2(new_n730), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n363), .B(new_n1180), .C1(G150), .C2(new_n753), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n743), .A2(KEYINPUT125), .A3(G132), .ZN(new_n1182));
  AOI21_X1  g0982(.A(KEYINPUT125), .B1(new_n743), .B2(G132), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G50), .B2(new_n755), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1096), .A2(new_n739), .B1(G137), .B2(new_n732), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1181), .A2(new_n1182), .A3(new_n1184), .A4(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n726), .B1(new_n1178), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n929), .B1(new_n860), .B2(new_n779), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1187), .B(new_n1188), .C1(new_n221), .C2(new_n807), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1170), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1169), .A2(new_n1046), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1191), .A2(new_n961), .A3(new_n1079), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1190), .A2(new_n1192), .ZN(G381));
  OAI21_X1  g0993(.A(new_n1113), .B1(new_n1078), .B2(new_n936), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1085), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1084), .B1(new_n1075), .B2(new_n682), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1083), .A2(new_n1080), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1194), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1139), .A2(new_n1199), .A3(new_n1167), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1200), .A2(G384), .A3(G381), .ZN(new_n1201));
  INV_X1    g1001(.A(G390), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n979), .A2(new_n980), .A3(new_n1202), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(new_n1203), .A2(G396), .A3(G393), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1201), .A2(new_n1204), .ZN(G407));
  OAI211_X1 g1005(.A(G407), .B(G213), .C1(G343), .C2(new_n1200), .ZN(G409));
  XNOR2_X1  g1006(.A(new_n977), .B(G390), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(G393), .B(G396), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n977), .A2(G390), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1203), .A2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1209), .B1(new_n1208), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT61), .ZN(new_n1213));
  INV_X1    g1013(.A(G213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1214), .A2(G343), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  AND4_X1   g1016(.A1(KEYINPUT126), .A2(new_n1166), .A3(new_n961), .A4(new_n1116), .ZN(new_n1217));
  AOI21_X1  g1017(.A(KEYINPUT126), .B1(new_n1137), .B2(new_n961), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1167), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1216), .B1(new_n1219), .B2(G378), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1199), .B1(new_n1139), .B2(new_n1167), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1169), .A2(KEYINPUT60), .A3(new_n1046), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1222), .A2(new_n682), .A3(new_n1079), .ZN(new_n1223));
  AOI21_X1  g1023(.A(KEYINPUT60), .B1(new_n1169), .B2(new_n1046), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1190), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(G384), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  OAI211_X1 g1027(.A(G384), .B(new_n1190), .C1(new_n1223), .C2(new_n1224), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1220), .A2(new_n1221), .A3(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT127), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(KEYINPUT62), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1213), .B1(new_n1230), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1215), .A2(G2897), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1227), .A2(new_n1228), .A3(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1234), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(G375), .A2(G378), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1166), .A2(new_n937), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1164), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT126), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n961), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1243), .B1(new_n1128), .B2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1137), .A2(KEYINPUT126), .A3(new_n961), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1242), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1215), .B1(new_n1247), .B2(new_n1199), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1229), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1240), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  XOR2_X1   g1050(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1251));
  OAI21_X1  g1051(.A(new_n1239), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1212), .B1(new_n1233), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1234), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1229), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1235), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(new_n1240), .B2(new_n1248), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT63), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1250), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1211), .A2(new_n1208), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n1208), .B2(new_n1207), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1230), .A2(KEYINPUT63), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1259), .A2(new_n1213), .A3(new_n1261), .A4(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1253), .A2(new_n1263), .ZN(G405));
  NAND2_X1  g1064(.A1(new_n1240), .A2(new_n1200), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1249), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1240), .A2(new_n1200), .A3(new_n1229), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(new_n1268), .B(new_n1261), .ZN(G402));
endmodule


