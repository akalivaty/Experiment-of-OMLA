

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589;

  XNOR2_X1 U325 ( .A(n380), .B(n322), .ZN(n323) );
  XNOR2_X1 U326 ( .A(n408), .B(KEYINPUT64), .ZN(n409) );
  XNOR2_X1 U327 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U328 ( .A(n410), .B(n409), .ZN(n534) );
  XNOR2_X1 U329 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U330 ( .A(KEYINPUT123), .B(KEYINPUT55), .ZN(n457) );
  XNOR2_X1 U331 ( .A(n331), .B(n330), .ZN(n335) );
  XNOR2_X1 U332 ( .A(n458), .B(n457), .ZN(n459) );
  INV_X1 U333 ( .A(G190GAT), .ZN(n461) );
  XNOR2_X1 U334 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U335 ( .A(n464), .B(n463), .ZN(G1351GAT) );
  XOR2_X1 U336 ( .A(G183GAT), .B(KEYINPUT88), .Z(n294) );
  XNOR2_X1 U337 ( .A(G169GAT), .B(KEYINPUT89), .ZN(n293) );
  XNOR2_X1 U338 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U339 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n296) );
  XNOR2_X1 U340 ( .A(G190GAT), .B(KEYINPUT18), .ZN(n295) );
  XNOR2_X1 U341 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U342 ( .A(n298), .B(n297), .Z(n321) );
  XOR2_X1 U343 ( .A(G43GAT), .B(G134GAT), .Z(n381) );
  XNOR2_X1 U344 ( .A(G99GAT), .B(G71GAT), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n299), .B(G120GAT), .ZN(n333) );
  XOR2_X1 U346 ( .A(n381), .B(n333), .Z(n301) );
  NAND2_X1 U347 ( .A1(G227GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U348 ( .A(n301), .B(n300), .ZN(n303) );
  XNOR2_X1 U349 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n302) );
  XNOR2_X1 U350 ( .A(n302), .B(KEYINPUT86), .ZN(n425) );
  XOR2_X1 U351 ( .A(n303), .B(n425), .Z(n305) );
  XNOR2_X1 U352 ( .A(KEYINPUT20), .B(G176GAT), .ZN(n304) );
  XNOR2_X1 U353 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U354 ( .A(G15GAT), .B(G127GAT), .Z(n367) );
  XOR2_X1 U355 ( .A(n306), .B(n367), .Z(n308) );
  XNOR2_X1 U356 ( .A(KEYINPUT90), .B(KEYINPUT87), .ZN(n307) );
  XOR2_X1 U357 ( .A(n308), .B(n307), .Z(n309) );
  XNOR2_X1 U358 ( .A(n321), .B(n309), .ZN(n467) );
  INV_X1 U359 ( .A(n467), .ZN(n536) );
  XOR2_X1 U360 ( .A(KEYINPUT54), .B(KEYINPUT122), .Z(n412) );
  XOR2_X1 U361 ( .A(G36GAT), .B(G8GAT), .Z(n345) );
  XOR2_X1 U362 ( .A(G64GAT), .B(KEYINPUT75), .Z(n311) );
  XNOR2_X1 U363 ( .A(G176GAT), .B(G204GAT), .ZN(n310) );
  XNOR2_X1 U364 ( .A(n311), .B(n310), .ZN(n324) );
  XOR2_X1 U365 ( .A(KEYINPUT102), .B(n324), .Z(n316) );
  XOR2_X1 U366 ( .A(KEYINPUT93), .B(G218GAT), .Z(n313) );
  XNOR2_X1 U367 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n312) );
  XNOR2_X1 U368 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U369 ( .A(G197GAT), .B(n314), .Z(n444) );
  XNOR2_X1 U370 ( .A(n444), .B(G92GAT), .ZN(n315) );
  XNOR2_X1 U371 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U372 ( .A(n345), .B(n317), .Z(n319) );
  NAND2_X1 U373 ( .A1(G226GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U375 ( .A(n321), .B(n320), .ZN(n484) );
  XOR2_X1 U376 ( .A(G85GAT), .B(G92GAT), .Z(n380) );
  AND2_X1 U377 ( .A1(G230GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U378 ( .A(n325), .B(KEYINPUT73), .ZN(n331) );
  XOR2_X1 U379 ( .A(G57GAT), .B(KEYINPUT13), .Z(n374) );
  XOR2_X1 U380 ( .A(n374), .B(KEYINPUT32), .Z(n329) );
  XOR2_X1 U381 ( .A(KEYINPUT31), .B(KEYINPUT72), .Z(n327) );
  XNOR2_X1 U382 ( .A(KEYINPUT33), .B(KEYINPUT74), .ZN(n326) );
  XOR2_X1 U383 ( .A(n327), .B(n326), .Z(n328) );
  XNOR2_X1 U384 ( .A(G106GAT), .B(G78GAT), .ZN(n332) );
  XNOR2_X1 U385 ( .A(n332), .B(G148GAT), .ZN(n440) );
  XNOR2_X1 U386 ( .A(n333), .B(n440), .ZN(n334) );
  XNOR2_X1 U387 ( .A(n335), .B(n334), .ZN(n578) );
  INV_X1 U388 ( .A(KEYINPUT41), .ZN(n336) );
  XNOR2_X1 U389 ( .A(n578), .B(n336), .ZN(n553) );
  XOR2_X1 U390 ( .A(G113GAT), .B(G15GAT), .Z(n338) );
  XNOR2_X1 U391 ( .A(G169GAT), .B(G197GAT), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U393 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n340) );
  XNOR2_X1 U394 ( .A(KEYINPUT29), .B(KEYINPUT67), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U396 ( .A(n342), .B(n341), .ZN(n355) );
  XOR2_X1 U397 ( .A(G22GAT), .B(G141GAT), .Z(n344) );
  XNOR2_X1 U398 ( .A(G50GAT), .B(G43GAT), .ZN(n343) );
  XNOR2_X1 U399 ( .A(n344), .B(n343), .ZN(n346) );
  XOR2_X1 U400 ( .A(n346), .B(n345), .Z(n353) );
  XOR2_X1 U401 ( .A(G29GAT), .B(KEYINPUT7), .Z(n348) );
  XNOR2_X1 U402 ( .A(KEYINPUT70), .B(KEYINPUT8), .ZN(n347) );
  XNOR2_X1 U403 ( .A(n348), .B(n347), .ZN(n391) );
  XOR2_X1 U404 ( .A(n391), .B(KEYINPUT69), .Z(n350) );
  NAND2_X1 U405 ( .A1(G229GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U407 ( .A(G1GAT), .B(KEYINPUT71), .Z(n375) );
  XNOR2_X1 U408 ( .A(n351), .B(n375), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U410 ( .A(n355), .B(n354), .ZN(n563) );
  INV_X1 U411 ( .A(n563), .ZN(n574) );
  NOR2_X1 U412 ( .A1(n553), .A2(n574), .ZN(n357) );
  INV_X1 U413 ( .A(KEYINPUT46), .ZN(n356) );
  XNOR2_X1 U414 ( .A(n357), .B(n356), .ZN(n401) );
  XOR2_X1 U415 ( .A(G22GAT), .B(G155GAT), .Z(n439) );
  XOR2_X1 U416 ( .A(n439), .B(KEYINPUT84), .Z(n359) );
  NAND2_X1 U417 ( .A1(G231GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U418 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U419 ( .A(KEYINPUT85), .B(KEYINPUT12), .Z(n361) );
  XNOR2_X1 U420 ( .A(KEYINPUT15), .B(KEYINPUT83), .ZN(n360) );
  XNOR2_X1 U421 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U422 ( .A(n363), .B(n362), .Z(n369) );
  XOR2_X1 U423 ( .A(KEYINPUT82), .B(KEYINPUT14), .Z(n365) );
  XNOR2_X1 U424 ( .A(G8GAT), .B(G64GAT), .ZN(n364) );
  XNOR2_X1 U425 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U426 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U427 ( .A(n369), .B(n368), .ZN(n373) );
  XOR2_X1 U428 ( .A(G78GAT), .B(G211GAT), .Z(n371) );
  XNOR2_X1 U429 ( .A(G183GAT), .B(G71GAT), .ZN(n370) );
  XNOR2_X1 U430 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U431 ( .A(n373), .B(n372), .Z(n377) );
  XNOR2_X1 U432 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U433 ( .A(n377), .B(n376), .ZN(n569) );
  INV_X1 U434 ( .A(n569), .ZN(n583) );
  XOR2_X1 U435 ( .A(KEYINPUT77), .B(KEYINPUT79), .Z(n379) );
  XNOR2_X1 U436 ( .A(G190GAT), .B(G99GAT), .ZN(n378) );
  XNOR2_X1 U437 ( .A(n379), .B(n378), .ZN(n399) );
  XOR2_X1 U438 ( .A(n380), .B(G218GAT), .Z(n383) );
  XNOR2_X1 U439 ( .A(G36GAT), .B(n381), .ZN(n382) );
  XNOR2_X1 U440 ( .A(n383), .B(n382), .ZN(n395) );
  XOR2_X1 U441 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n385) );
  XNOR2_X1 U442 ( .A(KEYINPUT78), .B(KEYINPUT81), .ZN(n384) );
  XNOR2_X1 U443 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U444 ( .A(KEYINPUT66), .B(KEYINPUT80), .Z(n387) );
  XNOR2_X1 U445 ( .A(G106GAT), .B(KEYINPUT9), .ZN(n386) );
  XNOR2_X1 U446 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U447 ( .A(n389), .B(n388), .Z(n393) );
  XNOR2_X1 U448 ( .A(G50GAT), .B(KEYINPUT76), .ZN(n390) );
  XNOR2_X1 U449 ( .A(n390), .B(G162GAT), .ZN(n452) );
  XNOR2_X1 U450 ( .A(n391), .B(n452), .ZN(n392) );
  XNOR2_X1 U451 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U452 ( .A(n395), .B(n394), .Z(n397) );
  NAND2_X1 U453 ( .A1(G232GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U455 ( .A(n399), .B(n398), .Z(n460) );
  AND2_X1 U456 ( .A1(n583), .A2(n460), .ZN(n400) );
  NAND2_X1 U457 ( .A1(n401), .A2(n400), .ZN(n402) );
  XNOR2_X1 U458 ( .A(n402), .B(KEYINPUT47), .ZN(n407) );
  XNOR2_X1 U459 ( .A(KEYINPUT36), .B(n460), .ZN(n586) );
  NOR2_X1 U460 ( .A1(n586), .A2(n583), .ZN(n403) );
  XNOR2_X1 U461 ( .A(KEYINPUT45), .B(n403), .ZN(n404) );
  NAND2_X1 U462 ( .A1(n404), .A2(n578), .ZN(n405) );
  NOR2_X1 U463 ( .A1(n405), .A2(n563), .ZN(n406) );
  NOR2_X1 U464 ( .A1(n407), .A2(n406), .ZN(n410) );
  INV_X1 U465 ( .A(KEYINPUT48), .ZN(n408) );
  NAND2_X1 U466 ( .A1(n484), .A2(n534), .ZN(n411) );
  XNOR2_X1 U467 ( .A(n412), .B(n411), .ZN(n437) );
  XOR2_X1 U468 ( .A(KEYINPUT101), .B(G148GAT), .Z(n414) );
  XNOR2_X1 U469 ( .A(G127GAT), .B(G120GAT), .ZN(n413) );
  XNOR2_X1 U470 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U471 ( .A(G85GAT), .B(KEYINPUT79), .Z(n416) );
  XNOR2_X1 U472 ( .A(G134GAT), .B(G155GAT), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U474 ( .A(n418), .B(n417), .ZN(n436) );
  XOR2_X1 U475 ( .A(G57GAT), .B(KEYINPUT99), .Z(n420) );
  XNOR2_X1 U476 ( .A(KEYINPUT100), .B(KEYINPUT4), .ZN(n419) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n424) );
  XOR2_X1 U478 ( .A(KEYINPUT5), .B(KEYINPUT97), .Z(n422) );
  XNOR2_X1 U479 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n421) );
  XNOR2_X1 U480 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U481 ( .A(n424), .B(n423), .Z(n430) );
  XOR2_X1 U482 ( .A(G162GAT), .B(n425), .Z(n427) );
  NAND2_X1 U483 ( .A1(G225GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U485 ( .A(G29GAT), .B(n428), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U487 ( .A(n431), .B(KEYINPUT98), .Z(n434) );
  XNOR2_X1 U488 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n432), .B(KEYINPUT2), .ZN(n451) );
  XNOR2_X1 U490 ( .A(G1GAT), .B(n451), .ZN(n433) );
  XNOR2_X1 U491 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n523) );
  NAND2_X1 U493 ( .A1(n437), .A2(n523), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n438), .B(KEYINPUT65), .ZN(n572) );
  XOR2_X1 U495 ( .A(n440), .B(n439), .Z(n442) );
  NAND2_X1 U496 ( .A1(G228GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n456) );
  XOR2_X1 U499 ( .A(G204GAT), .B(KEYINPUT95), .Z(n446) );
  XNOR2_X1 U500 ( .A(KEYINPUT23), .B(KEYINPUT96), .ZN(n445) );
  XNOR2_X1 U501 ( .A(n446), .B(n445), .ZN(n450) );
  XOR2_X1 U502 ( .A(KEYINPUT94), .B(KEYINPUT22), .Z(n448) );
  XNOR2_X1 U503 ( .A(KEYINPUT92), .B(KEYINPUT24), .ZN(n447) );
  XNOR2_X1 U504 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U505 ( .A(n450), .B(n449), .Z(n454) );
  XNOR2_X1 U506 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U507 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U508 ( .A(n456), .B(n455), .ZN(n475) );
  NAND2_X1 U509 ( .A1(n572), .A2(n475), .ZN(n458) );
  NOR2_X1 U510 ( .A1(n536), .A2(n459), .ZN(n570) );
  INV_X1 U511 ( .A(n460), .ZN(n559) );
  NAND2_X1 U512 ( .A1(n570), .A2(n559), .ZN(n464) );
  XOR2_X1 U513 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n462) );
  NAND2_X1 U514 ( .A1(n563), .A2(n578), .ZN(n495) );
  INV_X1 U515 ( .A(n495), .ZN(n481) );
  NOR2_X1 U516 ( .A1(n467), .A2(n475), .ZN(n465) );
  XNOR2_X1 U517 ( .A(KEYINPUT26), .B(n465), .ZN(n573) );
  XOR2_X1 U518 ( .A(KEYINPUT27), .B(n484), .Z(n474) );
  INV_X1 U519 ( .A(n474), .ZN(n466) );
  NAND2_X1 U520 ( .A1(n573), .A2(n466), .ZN(n471) );
  NAND2_X1 U521 ( .A1(n467), .A2(n484), .ZN(n468) );
  NAND2_X1 U522 ( .A1(n475), .A2(n468), .ZN(n469) );
  XOR2_X1 U523 ( .A(KEYINPUT25), .B(n469), .Z(n470) );
  NAND2_X1 U524 ( .A1(n471), .A2(n470), .ZN(n472) );
  NAND2_X1 U525 ( .A1(n472), .A2(n523), .ZN(n473) );
  XNOR2_X1 U526 ( .A(n473), .B(KEYINPUT103), .ZN(n478) );
  NOR2_X1 U527 ( .A1(n523), .A2(n474), .ZN(n549) );
  XNOR2_X1 U528 ( .A(n475), .B(KEYINPUT28), .ZN(n530) );
  NAND2_X1 U529 ( .A1(n549), .A2(n530), .ZN(n535) );
  XNOR2_X1 U530 ( .A(KEYINPUT91), .B(n536), .ZN(n476) );
  NOR2_X1 U531 ( .A1(n535), .A2(n476), .ZN(n477) );
  NOR2_X1 U532 ( .A1(n478), .A2(n477), .ZN(n492) );
  NOR2_X1 U533 ( .A1(n559), .A2(n583), .ZN(n479) );
  XOR2_X1 U534 ( .A(KEYINPUT16), .B(n479), .Z(n480) );
  NOR2_X1 U535 ( .A1(n492), .A2(n480), .ZN(n509) );
  NAND2_X1 U536 ( .A1(n481), .A2(n509), .ZN(n490) );
  NOR2_X1 U537 ( .A1(n523), .A2(n490), .ZN(n482) );
  XOR2_X1 U538 ( .A(KEYINPUT34), .B(n482), .Z(n483) );
  XNOR2_X1 U539 ( .A(G1GAT), .B(n483), .ZN(G1324GAT) );
  INV_X1 U540 ( .A(n484), .ZN(n526) );
  NOR2_X1 U541 ( .A1(n526), .A2(n490), .ZN(n485) );
  XOR2_X1 U542 ( .A(KEYINPUT104), .B(n485), .Z(n486) );
  XNOR2_X1 U543 ( .A(G8GAT), .B(n486), .ZN(G1325GAT) );
  NOR2_X1 U544 ( .A1(n536), .A2(n490), .ZN(n488) );
  XNOR2_X1 U545 ( .A(KEYINPUT105), .B(KEYINPUT35), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U547 ( .A(G15GAT), .B(n489), .Z(G1326GAT) );
  NOR2_X1 U548 ( .A1(n530), .A2(n490), .ZN(n491) );
  XOR2_X1 U549 ( .A(G22GAT), .B(n491), .Z(G1327GAT) );
  XNOR2_X1 U550 ( .A(KEYINPUT39), .B(KEYINPUT106), .ZN(n498) );
  NOR2_X1 U551 ( .A1(n492), .A2(n586), .ZN(n493) );
  NAND2_X1 U552 ( .A1(n583), .A2(n493), .ZN(n494) );
  XOR2_X1 U553 ( .A(KEYINPUT37), .B(n494), .Z(n522) );
  NOR2_X1 U554 ( .A1(n522), .A2(n495), .ZN(n496) );
  XOR2_X1 U555 ( .A(KEYINPUT38), .B(n496), .Z(n507) );
  NOR2_X1 U556 ( .A1(n523), .A2(n507), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U558 ( .A(G29GAT), .B(n499), .ZN(G1328GAT) );
  XNOR2_X1 U559 ( .A(G36GAT), .B(KEYINPUT107), .ZN(n501) );
  NOR2_X1 U560 ( .A1(n526), .A2(n507), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n501), .B(n500), .ZN(G1329GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT40), .B(KEYINPUT110), .Z(n503) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(KEYINPUT109), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n503), .B(n502), .ZN(n505) );
  NOR2_X1 U565 ( .A1(n507), .A2(n536), .ZN(n504) );
  XOR2_X1 U566 ( .A(n505), .B(n504), .Z(n506) );
  XNOR2_X1 U567 ( .A(KEYINPUT108), .B(n506), .ZN(G1330GAT) );
  NOR2_X1 U568 ( .A1(n507), .A2(n530), .ZN(n508) );
  XOR2_X1 U569 ( .A(G50GAT), .B(n508), .Z(G1331GAT) );
  XNOR2_X1 U570 ( .A(n553), .B(KEYINPUT111), .ZN(n565) );
  NAND2_X1 U571 ( .A1(n574), .A2(n565), .ZN(n521) );
  INV_X1 U572 ( .A(n521), .ZN(n510) );
  NAND2_X1 U573 ( .A1(n510), .A2(n509), .ZN(n517) );
  NOR2_X1 U574 ( .A1(n523), .A2(n517), .ZN(n512) );
  XNOR2_X1 U575 ( .A(KEYINPUT42), .B(KEYINPUT112), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U577 ( .A(G57GAT), .B(n513), .Z(G1332GAT) );
  NOR2_X1 U578 ( .A1(n526), .A2(n517), .ZN(n515) );
  XNOR2_X1 U579 ( .A(G64GAT), .B(KEYINPUT113), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(G1333GAT) );
  NOR2_X1 U581 ( .A1(n536), .A2(n517), .ZN(n516) );
  XOR2_X1 U582 ( .A(G71GAT), .B(n516), .Z(G1334GAT) );
  NOR2_X1 U583 ( .A1(n530), .A2(n517), .ZN(n519) );
  XNOR2_X1 U584 ( .A(KEYINPUT43), .B(KEYINPUT114), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U586 ( .A(G78GAT), .B(n520), .ZN(G1335GAT) );
  OR2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n529) );
  NOR2_X1 U588 ( .A1(n523), .A2(n529), .ZN(n525) );
  XNOR2_X1 U589 ( .A(G85GAT), .B(KEYINPUT115), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(G1336GAT) );
  NOR2_X1 U591 ( .A1(n526), .A2(n529), .ZN(n527) );
  XOR2_X1 U592 ( .A(G92GAT), .B(n527), .Z(G1337GAT) );
  NOR2_X1 U593 ( .A1(n536), .A2(n529), .ZN(n528) );
  XOR2_X1 U594 ( .A(G99GAT), .B(n528), .Z(G1338GAT) );
  NOR2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n532) );
  XNOR2_X1 U596 ( .A(KEYINPUT116), .B(KEYINPUT44), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U598 ( .A(G106GAT), .B(n533), .Z(G1339GAT) );
  NOR2_X1 U599 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U600 ( .A1(n534), .A2(n537), .ZN(n538) );
  XNOR2_X1 U601 ( .A(n538), .B(KEYINPUT117), .ZN(n546) );
  NAND2_X1 U602 ( .A1(n546), .A2(n563), .ZN(n539) );
  XNOR2_X1 U603 ( .A(n539), .B(KEYINPUT118), .ZN(n540) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(n540), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .Z(n542) );
  NAND2_X1 U606 ( .A1(n546), .A2(n565), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(G1341GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n544) );
  NAND2_X1 U609 ( .A1(n546), .A2(n569), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n545), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U613 ( .A1(n546), .A2(n559), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  AND2_X1 U615 ( .A1(n549), .A2(n573), .ZN(n550) );
  NAND2_X1 U616 ( .A1(n534), .A2(n550), .ZN(n552) );
  INV_X1 U617 ( .A(n552), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n563), .A2(n560), .ZN(n551) );
  XNOR2_X1 U619 ( .A(G141GAT), .B(n551), .ZN(G1344GAT) );
  NOR2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n555) );
  XNOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(n556), .ZN(G1345GAT) );
  NAND2_X1 U624 ( .A1(n560), .A2(n569), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n557), .B(KEYINPUT120), .ZN(n558) );
  XNOR2_X1 U626 ( .A(G155GAT), .B(n558), .ZN(G1346GAT) );
  XOR2_X1 U627 ( .A(G162GAT), .B(KEYINPUT121), .Z(n562) );
  NAND2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1347GAT) );
  NAND2_X1 U630 ( .A1(n570), .A2(n563), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n567) );
  NAND2_X1 U633 ( .A1(n570), .A2(n565), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(G176GAT), .B(n568), .ZN(G1349GAT) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U638 ( .A1(n572), .A2(n573), .ZN(n585) );
  NOR2_X1 U639 ( .A1(n574), .A2(n585), .ZN(n576) );
  XNOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(n577), .ZN(G1352GAT) );
  NOR2_X1 U643 ( .A1(n585), .A2(n578), .ZN(n582) );
  XOR2_X1 U644 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n580) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NOR2_X1 U648 ( .A1(n583), .A2(n585), .ZN(n584) );
  XOR2_X1 U649 ( .A(G211GAT), .B(n584), .Z(G1354GAT) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n588) );
  XNOR2_X1 U651 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

