

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588;

  XNOR2_X1 U324 ( .A(G211GAT), .B(KEYINPUT85), .ZN(n336) );
  XOR2_X1 U325 ( .A(G8GAT), .B(G183GAT), .Z(n438) );
  XNOR2_X1 U326 ( .A(n333), .B(n332), .ZN(n334) );
  NOR2_X1 U327 ( .A1(n534), .A2(n478), .ZN(n567) );
  XNOR2_X1 U328 ( .A(n456), .B(KEYINPUT38), .ZN(n502) );
  XNOR2_X1 U329 ( .A(n348), .B(n347), .ZN(n522) );
  AND2_X1 U330 ( .A1(G231GAT), .A2(G233GAT), .ZN(n292) );
  XOR2_X1 U331 ( .A(n337), .B(KEYINPUT21), .Z(n293) );
  XNOR2_X1 U332 ( .A(n335), .B(n334), .ZN(n459) );
  XNOR2_X1 U333 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U334 ( .A(n448), .B(n316), .ZN(n321) );
  XNOR2_X1 U335 ( .A(KEYINPUT114), .B(KEYINPUT46), .ZN(n460) );
  XNOR2_X1 U336 ( .A(n461), .B(n460), .ZN(n463) );
  NOR2_X1 U337 ( .A1(n413), .A2(n412), .ZN(n414) );
  XNOR2_X1 U338 ( .A(n444), .B(n292), .ZN(n445) );
  INV_X1 U339 ( .A(n586), .ZN(n453) );
  XNOR2_X1 U340 ( .A(n339), .B(KEYINPUT94), .ZN(n340) );
  XNOR2_X1 U341 ( .A(n471), .B(KEYINPUT54), .ZN(n472) );
  XNOR2_X1 U342 ( .A(n446), .B(n445), .ZN(n447) );
  NAND2_X1 U343 ( .A1(n453), .A2(n583), .ZN(n454) );
  XNOR2_X1 U344 ( .A(n384), .B(n340), .ZN(n341) );
  XNOR2_X1 U345 ( .A(KEYINPUT121), .B(KEYINPUT55), .ZN(n476) );
  XNOR2_X1 U346 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U347 ( .A(n452), .B(n451), .Z(n563) );
  XOR2_X1 U348 ( .A(n404), .B(n403), .Z(n525) );
  XOR2_X1 U349 ( .A(n371), .B(n370), .Z(n519) );
  XNOR2_X1 U350 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U351 ( .A(G36GAT), .B(KEYINPUT104), .ZN(n457) );
  XNOR2_X1 U352 ( .A(n482), .B(n481), .ZN(G1349GAT) );
  XNOR2_X1 U353 ( .A(n458), .B(n457), .ZN(G1329GAT) );
  XOR2_X1 U354 ( .A(G36GAT), .B(G50GAT), .Z(n295) );
  XOR2_X1 U355 ( .A(G141GAT), .B(G22GAT), .Z(n374) );
  XOR2_X1 U356 ( .A(G113GAT), .B(G1GAT), .Z(n361) );
  XNOR2_X1 U357 ( .A(n374), .B(n361), .ZN(n294) );
  XNOR2_X1 U358 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U359 ( .A(n296), .B(G15GAT), .Z(n303) );
  XOR2_X1 U360 ( .A(G29GAT), .B(G43GAT), .Z(n298) );
  XNOR2_X1 U361 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n297) );
  XNOR2_X1 U362 ( .A(n298), .B(n297), .ZN(n424) );
  XOR2_X1 U363 ( .A(n424), .B(KEYINPUT68), .Z(n300) );
  NAND2_X1 U364 ( .A1(G229GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U365 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U366 ( .A(G169GAT), .B(n301), .ZN(n302) );
  XNOR2_X1 U367 ( .A(n303), .B(n302), .ZN(n311) );
  XOR2_X1 U368 ( .A(KEYINPUT67), .B(KEYINPUT29), .Z(n305) );
  XNOR2_X1 U369 ( .A(G197GAT), .B(G8GAT), .ZN(n304) );
  XNOR2_X1 U370 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U371 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n307) );
  XNOR2_X1 U372 ( .A(KEYINPUT70), .B(KEYINPUT69), .ZN(n306) );
  XNOR2_X1 U373 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U374 ( .A(n309), .B(n308), .Z(n310) );
  XOR2_X1 U375 ( .A(n311), .B(n310), .Z(n574) );
  INV_X1 U376 ( .A(n574), .ZN(n561) );
  XOR2_X1 U377 ( .A(KEYINPUT71), .B(KEYINPUT13), .Z(n313) );
  XNOR2_X1 U378 ( .A(G71GAT), .B(G57GAT), .ZN(n312) );
  XNOR2_X1 U379 ( .A(n313), .B(n312), .ZN(n448) );
  NAND2_X1 U380 ( .A1(G230GAT), .A2(G233GAT), .ZN(n315) );
  INV_X1 U381 ( .A(KEYINPUT31), .ZN(n314) );
  INV_X1 U382 ( .A(n321), .ZN(n320) );
  XOR2_X1 U383 ( .A(G64GAT), .B(G92GAT), .Z(n318) );
  XNOR2_X1 U384 ( .A(G176GAT), .B(G204GAT), .ZN(n317) );
  XNOR2_X1 U385 ( .A(n318), .B(n317), .ZN(n346) );
  INV_X1 U386 ( .A(n346), .ZN(n319) );
  NAND2_X1 U387 ( .A1(n320), .A2(n319), .ZN(n323) );
  NAND2_X1 U388 ( .A1(n321), .A2(n346), .ZN(n322) );
  NAND2_X1 U389 ( .A1(n323), .A2(n322), .ZN(n326) );
  XNOR2_X1 U390 ( .A(G106GAT), .B(G78GAT), .ZN(n324) );
  XNOR2_X1 U391 ( .A(n324), .B(G148GAT), .ZN(n383) );
  XOR2_X1 U392 ( .A(G120GAT), .B(n383), .Z(n325) );
  XNOR2_X1 U393 ( .A(n326), .B(n325), .ZN(n328) );
  INV_X1 U394 ( .A(KEYINPUT72), .ZN(n327) );
  XNOR2_X1 U395 ( .A(n328), .B(n327), .ZN(n335) );
  XNOR2_X1 U396 ( .A(G99GAT), .B(G85GAT), .ZN(n329) );
  XNOR2_X1 U397 ( .A(n329), .B(KEYINPUT73), .ZN(n418) );
  XNOR2_X1 U398 ( .A(n418), .B(KEYINPUT33), .ZN(n333) );
  XOR2_X1 U399 ( .A(KEYINPUT74), .B(KEYINPUT32), .Z(n331) );
  XNOR2_X1 U400 ( .A(KEYINPUT76), .B(KEYINPUT75), .ZN(n330) );
  XOR2_X1 U401 ( .A(n331), .B(n330), .Z(n332) );
  INV_X1 U402 ( .A(n459), .ZN(n580) );
  NAND2_X1 U403 ( .A1(n561), .A2(n580), .ZN(n487) );
  XOR2_X1 U404 ( .A(G36GAT), .B(G190GAT), .Z(n421) );
  XNOR2_X1 U405 ( .A(n336), .B(KEYINPUT86), .ZN(n337) );
  XNOR2_X1 U406 ( .A(G197GAT), .B(G218GAT), .ZN(n338) );
  XNOR2_X1 U407 ( .A(n293), .B(n338), .ZN(n384) );
  XOR2_X1 U408 ( .A(n438), .B(KEYINPUT93), .Z(n339) );
  XOR2_X1 U409 ( .A(n421), .B(n341), .Z(n343) );
  NAND2_X1 U410 ( .A1(G226GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U411 ( .A(n343), .B(n342), .ZN(n348) );
  XOR2_X1 U412 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n345) );
  XNOR2_X1 U413 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n344) );
  XNOR2_X1 U414 ( .A(n345), .B(n344), .ZN(n399) );
  XOR2_X1 U415 ( .A(n399), .B(n346), .Z(n347) );
  XOR2_X1 U416 ( .A(KEYINPUT27), .B(n522), .Z(n410) );
  XNOR2_X1 U417 ( .A(G134GAT), .B(G120GAT), .ZN(n349) );
  XNOR2_X1 U418 ( .A(n349), .B(KEYINPUT0), .ZN(n400) );
  XOR2_X1 U419 ( .A(KEYINPUT92), .B(KEYINPUT4), .Z(n351) );
  XNOR2_X1 U420 ( .A(G141GAT), .B(G148GAT), .ZN(n350) );
  XNOR2_X1 U421 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U422 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n353) );
  XNOR2_X1 U423 ( .A(KEYINPUT91), .B(G57GAT), .ZN(n352) );
  XNOR2_X1 U424 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U425 ( .A(n355), .B(n354), .Z(n367) );
  XOR2_X1 U426 ( .A(KEYINPUT5), .B(KEYINPUT88), .Z(n357) );
  XNOR2_X1 U427 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n356) );
  XNOR2_X1 U428 ( .A(n357), .B(n356), .ZN(n365) );
  XOR2_X1 U429 ( .A(G85GAT), .B(G162GAT), .Z(n359) );
  XNOR2_X1 U430 ( .A(G29GAT), .B(G127GAT), .ZN(n358) );
  XNOR2_X1 U431 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U432 ( .A(n361), .B(n360), .Z(n363) );
  NAND2_X1 U433 ( .A1(G225GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U434 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U435 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U436 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U437 ( .A(n400), .B(n368), .ZN(n371) );
  XNOR2_X1 U438 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n369) );
  XOR2_X1 U439 ( .A(n369), .B(KEYINPUT2), .Z(n381) );
  INV_X1 U440 ( .A(n381), .ZN(n370) );
  INV_X1 U441 ( .A(n519), .ZN(n549) );
  XOR2_X1 U442 ( .A(KEYINPUT23), .B(KEYINPUT87), .Z(n373) );
  XNOR2_X1 U443 ( .A(KEYINPUT84), .B(KEYINPUT22), .ZN(n372) );
  XNOR2_X1 U444 ( .A(n373), .B(n372), .ZN(n378) );
  XOR2_X1 U445 ( .A(KEYINPUT24), .B(G204GAT), .Z(n376) );
  XOR2_X1 U446 ( .A(G50GAT), .B(G162GAT), .Z(n423) );
  XNOR2_X1 U447 ( .A(n374), .B(n423), .ZN(n375) );
  XNOR2_X1 U448 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U449 ( .A(n378), .B(n377), .Z(n380) );
  NAND2_X1 U450 ( .A1(G228GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U451 ( .A(n380), .B(n379), .ZN(n382) );
  XNOR2_X1 U452 ( .A(n382), .B(n381), .ZN(n386) );
  XNOR2_X1 U453 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U454 ( .A(n386), .B(n385), .ZN(n475) );
  XOR2_X1 U455 ( .A(n475), .B(KEYINPUT28), .Z(n527) );
  OR2_X1 U456 ( .A1(n549), .A2(n527), .ZN(n387) );
  NOR2_X1 U457 ( .A1(n410), .A2(n387), .ZN(n532) );
  XOR2_X1 U458 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n389) );
  XNOR2_X1 U459 ( .A(KEYINPUT65), .B(G71GAT), .ZN(n388) );
  XNOR2_X1 U460 ( .A(n389), .B(n388), .ZN(n404) );
  XOR2_X1 U461 ( .A(G15GAT), .B(G127GAT), .Z(n439) );
  XOR2_X1 U462 ( .A(KEYINPUT83), .B(G190GAT), .Z(n391) );
  XNOR2_X1 U463 ( .A(G43GAT), .B(G99GAT), .ZN(n390) );
  XNOR2_X1 U464 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U465 ( .A(n439), .B(n392), .Z(n394) );
  NAND2_X1 U466 ( .A1(G227GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U467 ( .A(n394), .B(n393), .ZN(n398) );
  XOR2_X1 U468 ( .A(G183GAT), .B(G176GAT), .Z(n396) );
  XNOR2_X1 U469 ( .A(G113GAT), .B(KEYINPUT20), .ZN(n395) );
  XNOR2_X1 U470 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U471 ( .A(n398), .B(n397), .Z(n402) );
  XNOR2_X1 U472 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U473 ( .A(n402), .B(n401), .ZN(n403) );
  INV_X1 U474 ( .A(n525), .ZN(n534) );
  NAND2_X1 U475 ( .A1(n532), .A2(n534), .ZN(n405) );
  XNOR2_X1 U476 ( .A(n405), .B(KEYINPUT95), .ZN(n417) );
  NAND2_X1 U477 ( .A1(n525), .A2(n522), .ZN(n406) );
  XOR2_X1 U478 ( .A(KEYINPUT97), .B(n406), .Z(n407) );
  NAND2_X1 U479 ( .A1(n475), .A2(n407), .ZN(n408) );
  XNOR2_X1 U480 ( .A(KEYINPUT25), .B(n408), .ZN(n413) );
  NOR2_X1 U481 ( .A1(n525), .A2(n475), .ZN(n409) );
  XNOR2_X1 U482 ( .A(KEYINPUT26), .B(n409), .ZN(n572) );
  INV_X1 U483 ( .A(n572), .ZN(n411) );
  NOR2_X1 U484 ( .A1(n411), .A2(n410), .ZN(n546) );
  XNOR2_X1 U485 ( .A(KEYINPUT96), .B(n546), .ZN(n412) );
  XNOR2_X1 U486 ( .A(KEYINPUT98), .B(n414), .ZN(n415) );
  NOR2_X1 U487 ( .A1(n519), .A2(n415), .ZN(n416) );
  NOR2_X1 U488 ( .A1(n417), .A2(n416), .ZN(n485) );
  XNOR2_X1 U489 ( .A(KEYINPUT103), .B(KEYINPUT36), .ZN(n435) );
  XOR2_X1 U490 ( .A(n418), .B(G92GAT), .Z(n420) );
  NAND2_X1 U491 ( .A1(G232GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U492 ( .A(n420), .B(n419), .ZN(n422) );
  XOR2_X1 U493 ( .A(n422), .B(n421), .Z(n426) );
  XNOR2_X1 U494 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U495 ( .A(n426), .B(n425), .ZN(n434) );
  XOR2_X1 U496 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n428) );
  XNOR2_X1 U497 ( .A(G218GAT), .B(KEYINPUT77), .ZN(n427) );
  XNOR2_X1 U498 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U499 ( .A(KEYINPUT9), .B(KEYINPUT64), .Z(n430) );
  XNOR2_X1 U500 ( .A(G134GAT), .B(G106GAT), .ZN(n429) );
  XNOR2_X1 U501 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U502 ( .A(n432), .B(n431), .Z(n433) );
  XNOR2_X1 U503 ( .A(n434), .B(n433), .ZN(n566) );
  XNOR2_X1 U504 ( .A(n435), .B(n566), .ZN(n586) );
  XOR2_X1 U505 ( .A(G64GAT), .B(G211GAT), .Z(n437) );
  XNOR2_X1 U506 ( .A(G22GAT), .B(G1GAT), .ZN(n436) );
  XNOR2_X1 U507 ( .A(n437), .B(n436), .ZN(n452) );
  XOR2_X1 U508 ( .A(n438), .B(G155GAT), .Z(n441) );
  XNOR2_X1 U509 ( .A(n439), .B(G78GAT), .ZN(n440) );
  XNOR2_X1 U510 ( .A(n441), .B(n440), .ZN(n446) );
  XOR2_X1 U511 ( .A(KEYINPUT15), .B(KEYINPUT78), .Z(n443) );
  XNOR2_X1 U512 ( .A(KEYINPUT80), .B(KEYINPUT79), .ZN(n442) );
  XNOR2_X1 U513 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U514 ( .A(n447), .B(KEYINPUT14), .Z(n450) );
  XNOR2_X1 U515 ( .A(n448), .B(KEYINPUT12), .ZN(n449) );
  XNOR2_X1 U516 ( .A(n450), .B(n449), .ZN(n451) );
  INV_X1 U517 ( .A(n563), .ZN(n583) );
  OR2_X1 U518 ( .A1(n485), .A2(n454), .ZN(n455) );
  XOR2_X1 U519 ( .A(KEYINPUT37), .B(n455), .Z(n518) );
  NOR2_X1 U520 ( .A1(n487), .A2(n518), .ZN(n456) );
  NAND2_X1 U521 ( .A1(n502), .A2(n522), .ZN(n458) );
  XOR2_X1 U522 ( .A(KEYINPUT41), .B(n459), .Z(n552) );
  XOR2_X1 U523 ( .A(n552), .B(KEYINPUT107), .Z(n536) );
  NAND2_X1 U524 ( .A1(n561), .A2(n552), .ZN(n461) );
  NOR2_X1 U525 ( .A1(n566), .A2(n563), .ZN(n462) );
  AND2_X1 U526 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U527 ( .A(n464), .B(KEYINPUT47), .ZN(n469) );
  NOR2_X1 U528 ( .A1(n586), .A2(n583), .ZN(n465) );
  XOR2_X1 U529 ( .A(KEYINPUT45), .B(n465), .Z(n466) );
  NOR2_X1 U530 ( .A1(n459), .A2(n466), .ZN(n467) );
  NAND2_X1 U531 ( .A1(n467), .A2(n574), .ZN(n468) );
  NAND2_X1 U532 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U533 ( .A(n470), .B(KEYINPUT48), .ZN(n547) );
  AND2_X1 U534 ( .A1(n522), .A2(n547), .ZN(n473) );
  INV_X1 U535 ( .A(KEYINPUT120), .ZN(n471) );
  XNOR2_X1 U536 ( .A(n473), .B(n472), .ZN(n474) );
  NOR2_X1 U537 ( .A1(n519), .A2(n474), .ZN(n573) );
  NAND2_X1 U538 ( .A1(n573), .A2(n475), .ZN(n477) );
  NAND2_X1 U539 ( .A1(n536), .A2(n567), .ZN(n482) );
  XOR2_X1 U540 ( .A(G176GAT), .B(KEYINPUT122), .Z(n480) );
  XNOR2_X1 U541 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n479) );
  XOR2_X1 U542 ( .A(KEYINPUT34), .B(KEYINPUT100), .Z(n489) );
  NOR2_X1 U543 ( .A1(n566), .A2(n583), .ZN(n483) );
  XOR2_X1 U544 ( .A(KEYINPUT16), .B(n483), .Z(n484) );
  NOR2_X1 U545 ( .A1(n485), .A2(n484), .ZN(n486) );
  XNOR2_X1 U546 ( .A(KEYINPUT99), .B(n486), .ZN(n505) );
  NOR2_X1 U547 ( .A1(n487), .A2(n505), .ZN(n495) );
  NAND2_X1 U548 ( .A1(n495), .A2(n519), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U550 ( .A(G1GAT), .B(n490), .Z(G1324GAT) );
  NAND2_X1 U551 ( .A1(n522), .A2(n495), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n491), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT35), .B(KEYINPUT101), .Z(n493) );
  NAND2_X1 U554 ( .A1(n495), .A2(n525), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U556 ( .A(G15GAT), .B(n494), .Z(G1326GAT) );
  NAND2_X1 U557 ( .A1(n495), .A2(n527), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n496), .B(KEYINPUT102), .ZN(n497) );
  XNOR2_X1 U559 ( .A(G22GAT), .B(n497), .ZN(G1327GAT) );
  XOR2_X1 U560 ( .A(G29GAT), .B(KEYINPUT39), .Z(n499) );
  NAND2_X1 U561 ( .A1(n502), .A2(n519), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  NAND2_X1 U563 ( .A1(n502), .A2(n525), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n500), .B(KEYINPUT40), .ZN(n501) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(n501), .ZN(G1330GAT) );
  XOR2_X1 U566 ( .A(G50GAT), .B(KEYINPUT105), .Z(n504) );
  NAND2_X1 U567 ( .A1(n527), .A2(n502), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(G1331GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n507) );
  NAND2_X1 U570 ( .A1(n574), .A2(n536), .ZN(n517) );
  NOR2_X1 U571 ( .A1(n505), .A2(n517), .ZN(n513) );
  NAND2_X1 U572 ( .A1(n513), .A2(n519), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U574 ( .A(G57GAT), .B(n508), .Z(G1332GAT) );
  NAND2_X1 U575 ( .A1(n522), .A2(n513), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n509), .B(KEYINPUT108), .ZN(n510) );
  XNOR2_X1 U577 ( .A(G64GAT), .B(n510), .ZN(G1333GAT) );
  XOR2_X1 U578 ( .A(G71GAT), .B(KEYINPUT109), .Z(n512) );
  NAND2_X1 U579 ( .A1(n513), .A2(n525), .ZN(n511) );
  XNOR2_X1 U580 ( .A(n512), .B(n511), .ZN(G1334GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n515) );
  NAND2_X1 U582 ( .A1(n513), .A2(n527), .ZN(n514) );
  XNOR2_X1 U583 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(n516), .ZN(G1335GAT) );
  XOR2_X1 U585 ( .A(G85GAT), .B(KEYINPUT111), .Z(n521) );
  NOR2_X1 U586 ( .A1(n518), .A2(n517), .ZN(n528) );
  NAND2_X1 U587 ( .A1(n528), .A2(n519), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(G1336GAT) );
  NAND2_X1 U589 ( .A1(n522), .A2(n528), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n523), .B(KEYINPUT112), .ZN(n524) );
  XNOR2_X1 U591 ( .A(G92GAT), .B(n524), .ZN(G1337GAT) );
  NAND2_X1 U592 ( .A1(n528), .A2(n525), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n526), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT44), .B(KEYINPUT113), .Z(n530) );
  NAND2_X1 U595 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  NAND2_X1 U598 ( .A1(n547), .A2(n532), .ZN(n533) );
  NOR2_X1 U599 ( .A1(n534), .A2(n533), .ZN(n543) );
  NAND2_X1 U600 ( .A1(n561), .A2(n543), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n535), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n538) );
  NAND2_X1 U603 ( .A1(n543), .A2(n536), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U605 ( .A(G120GAT), .B(n539), .Z(G1341GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n541) );
  NAND2_X1 U607 ( .A1(n543), .A2(n563), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U609 ( .A(G127GAT), .B(n542), .Z(G1342GAT) );
  XOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U611 ( .A1(n543), .A2(n566), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(G1343GAT) );
  XOR2_X1 U613 ( .A(G141GAT), .B(KEYINPUT117), .Z(n551) );
  NAND2_X1 U614 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n559) );
  NAND2_X1 U616 ( .A1(n559), .A2(n561), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1344GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n554) );
  NAND2_X1 U619 ( .A1(n559), .A2(n552), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(n555), .ZN(G1345GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n557) );
  NAND2_X1 U623 ( .A1(n559), .A2(n563), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U625 ( .A(G155GAT), .B(n558), .ZN(G1346GAT) );
  NAND2_X1 U626 ( .A1(n566), .A2(n559), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n567), .A2(n561), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U630 ( .A(G183GAT), .B(KEYINPUT123), .Z(n565) );
  NAND2_X1 U631 ( .A1(n567), .A2(n563), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1350GAT) );
  XNOR2_X1 U633 ( .A(G190GAT), .B(KEYINPUT124), .ZN(n571) );
  XOR2_X1 U634 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n569) );
  NAND2_X1 U635 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1351GAT) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n585) );
  NOR2_X1 U639 ( .A1(n574), .A2(n585), .ZN(n579) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT127), .Z(n576) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(KEYINPUT126), .B(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n585), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NOR2_X1 U648 ( .A1(n583), .A2(n585), .ZN(n584) );
  XOR2_X1 U649 ( .A(G211GAT), .B(n584), .Z(G1354GAT) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(KEYINPUT62), .B(n587), .Z(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

