//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n619, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1175, new_n1176, new_n1177;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT64), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n451), .B(new_n452), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  XNOR2_X1  g030(.A(G325), .B(KEYINPUT66), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OR2_X1    g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n463), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n465), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n463), .A2(new_n465), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n466), .A2(new_n471), .ZN(G160));
  NOR2_X1   g047(.A1(new_n461), .A2(new_n462), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n473), .A2(new_n465), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  OR2_X1    g056(.A1(G102), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G114), .C2(new_n465), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT67), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n485), .B1(new_n469), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n476), .A2(G126), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n474), .A2(KEYINPUT4), .A3(G138), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n484), .A2(new_n487), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G164));
  INV_X1    g066(.A(G543), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT5), .ZN(new_n493));
  OAI211_X1 g068(.A(KEYINPUT69), .B(new_n492), .C1(new_n493), .C2(KEYINPUT68), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n495), .B1(new_n496), .B2(KEYINPUT5), .ZN(new_n497));
  OAI21_X1  g072(.A(G543), .B1(new_n493), .B2(KEYINPUT69), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n494), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n499), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OR2_X1    g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n492), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G50), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n503), .A2(new_n504), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n499), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n502), .A2(new_n510), .ZN(G166));
  NAND3_X1  g086(.A1(new_n499), .A2(G89), .A3(new_n507), .ZN(new_n512));
  AND2_X1   g087(.A1(G63), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n499), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT7), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT7), .ZN(new_n517));
  NAND4_X1  g092(.A1(new_n517), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n505), .A2(G51), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n512), .A2(new_n514), .A3(new_n519), .ZN(G286));
  INV_X1    g095(.A(G286), .ZN(G168));
  INV_X1    g096(.A(G64), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n492), .B1(new_n495), .B2(KEYINPUT5), .ZN(new_n523));
  OAI21_X1  g098(.A(KEYINPUT69), .B1(new_n493), .B2(KEYINPUT68), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n522), .B1(new_n525), .B2(new_n494), .ZN(new_n526));
  AND2_X1   g101(.A1(G77), .A2(G543), .ZN(new_n527));
  OAI21_X1  g102(.A(G651), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n504), .ZN(new_n529));
  NOR2_X1   g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  OAI211_X1 g105(.A(G52), .B(G543), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n529), .A2(new_n530), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n533), .B1(new_n525), .B2(new_n494), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n532), .B1(new_n534), .B2(G90), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n528), .A2(new_n535), .ZN(G171));
  NAND3_X1  g111(.A1(new_n499), .A2(G81), .A3(new_n507), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n505), .A2(G43), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n537), .A2(KEYINPUT71), .A3(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(KEYINPUT71), .B1(new_n537), .B2(new_n538), .ZN(new_n541));
  AND2_X1   g116(.A1(G68), .A2(G543), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n542), .B1(new_n499), .B2(G56), .ZN(new_n543));
  OAI21_X1  g118(.A(G651), .B1(new_n543), .B2(KEYINPUT70), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n545), .B1(new_n525), .B2(new_n494), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT70), .ZN(new_n547));
  NOR3_X1   g122(.A1(new_n546), .A2(new_n547), .A3(new_n542), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n540), .A2(new_n541), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  OAI211_X1 g130(.A(G53), .B(G543), .C1(new_n529), .C2(new_n530), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(KEYINPUT72), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n556), .B(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n499), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n560), .B2(new_n501), .ZN(new_n561));
  AND3_X1   g136(.A1(new_n499), .A2(KEYINPUT73), .A3(new_n507), .ZN(new_n562));
  AOI21_X1  g137(.A(KEYINPUT73), .B1(new_n499), .B2(new_n507), .ZN(new_n563));
  INV_X1    g138(.A(G91), .ZN(new_n564));
  NOR3_X1   g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  XOR2_X1   g143(.A(G166), .B(KEYINPUT74), .Z(G303));
  INV_X1    g144(.A(KEYINPUT73), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n508), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n499), .A2(KEYINPUT73), .A3(new_n507), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n571), .A2(G87), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n505), .A2(G49), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n505), .A2(KEYINPUT75), .A3(G49), .ZN(new_n577));
  INV_X1    g152(.A(G74), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n525), .A2(new_n578), .A3(new_n494), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n576), .A2(new_n577), .B1(G651), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n573), .A2(new_n580), .ZN(G288));
  AOI22_X1  g156(.A1(new_n499), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n582), .A2(new_n501), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n505), .A2(G48), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT76), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(G86), .ZN(new_n587));
  NOR3_X1   g162(.A1(new_n562), .A2(new_n563), .A3(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n586), .A2(new_n589), .ZN(G305));
  AND2_X1   g165(.A1(G72), .A2(G543), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n591), .B1(new_n499), .B2(G60), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(G60), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(new_n525), .B2(new_n494), .ZN(new_n596));
  OAI21_X1  g171(.A(KEYINPUT77), .B1(new_n596), .B2(new_n591), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n594), .A2(new_n597), .A3(G651), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n534), .A2(G85), .B1(G47), .B2(new_n505), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(G290));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NOR2_X1   g176(.A1(G171), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT78), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n499), .A2(G66), .ZN(new_n604));
  INV_X1    g179(.A(G79), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(new_n492), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n606), .A2(G651), .B1(G54), .B2(new_n505), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n562), .A2(new_n563), .ZN(new_n608));
  AOI21_X1  g183(.A(KEYINPUT10), .B1(new_n608), .B2(G92), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n571), .A2(KEYINPUT10), .A3(G92), .A4(new_n572), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n607), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n603), .B1(G868), .B2(new_n613), .ZN(G284));
  OAI21_X1  g189(.A(new_n603), .B1(G868), .B2(new_n613), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(new_n566), .B2(G868), .ZN(G297));
  OAI21_X1  g192(.A(new_n616), .B1(new_n566), .B2(G868), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n613), .B1(new_n619), .B2(G860), .ZN(G148));
  NOR2_X1   g195(.A1(new_n549), .A2(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n613), .A2(new_n619), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT79), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n621), .B1(new_n623), .B2(G868), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n463), .A2(new_n467), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  INV_X1    g203(.A(G2100), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n474), .A2(G135), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n476), .A2(G123), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n465), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(G2096), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n630), .A2(new_n631), .A3(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(G2451), .B(G2454), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT82), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT81), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n643), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT80), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2427), .B(G2430), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(KEYINPUT14), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n654), .B1(new_n653), .B2(new_n651), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n647), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n647), .A2(new_n655), .ZN(new_n657));
  AND3_X1   g232(.A1(new_n656), .A2(G14), .A3(new_n657), .ZN(G401));
  INV_X1    g233(.A(KEYINPUT18), .ZN(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(KEYINPUT17), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n660), .A2(new_n661), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n659), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(new_n629), .ZN(new_n666));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n662), .B2(KEYINPUT18), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(new_n637), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n666), .B(new_n669), .ZN(G227));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT19), .Z(new_n672));
  XNOR2_X1  g247(.A(G1956), .B(G2474), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1961), .B(G1966), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT83), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT20), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n672), .A2(KEYINPUT84), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n673), .A2(new_n674), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n671), .B(KEYINPUT19), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n681), .B1(new_n682), .B2(new_n675), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n680), .B(new_n683), .Z(new_n684));
  NAND2_X1  g259(.A1(new_n677), .A2(new_n678), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n679), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(G229));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n695), .A2(G6), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G305), .B2(G16), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT32), .B(G1981), .Z(new_n698));
  AND2_X1   g273(.A1(new_n695), .A2(G23), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G288), .B2(G16), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT33), .B(G1976), .ZN(new_n701));
  AOI22_X1  g276(.A1(new_n697), .A2(new_n698), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(new_n700), .B2(new_n701), .ZN(new_n703));
  INV_X1    g278(.A(G22), .ZN(new_n704));
  OR3_X1    g279(.A1(new_n704), .A2(KEYINPUT85), .A3(G16), .ZN(new_n705));
  OAI21_X1  g280(.A(KEYINPUT85), .B1(new_n704), .B2(G16), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n705), .B(new_n706), .C1(G166), .C2(new_n695), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(G1971), .Z(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(new_n698), .B2(new_n697), .ZN(new_n709));
  OR3_X1    g284(.A1(new_n703), .A2(new_n709), .A3(KEYINPUT34), .ZN(new_n710));
  OAI21_X1  g285(.A(KEYINPUT34), .B1(new_n703), .B2(new_n709), .ZN(new_n711));
  MUX2_X1   g286(.A(G24), .B(G290), .S(G16), .Z(new_n712));
  AND2_X1   g287(.A1(new_n712), .A2(G1986), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(G1986), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n474), .A2(G131), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n476), .A2(G119), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n465), .A2(G107), .ZN(new_n717));
  OAI21_X1  g292(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n715), .B(new_n716), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  MUX2_X1   g294(.A(G25), .B(new_n719), .S(G29), .Z(new_n720));
  XOR2_X1   g295(.A(KEYINPUT35), .B(G1991), .Z(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n720), .B(new_n722), .ZN(new_n723));
  NOR3_X1   g298(.A1(new_n713), .A2(new_n714), .A3(new_n723), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n710), .A2(new_n711), .A3(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT36), .Z(new_n726));
  NOR2_X1   g301(.A1(G16), .A2(G19), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n550), .B2(G16), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT86), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(G1341), .Z(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT30), .B(G28), .ZN(new_n731));
  INV_X1    g306(.A(G29), .ZN(new_n732));
  OR2_X1    g307(.A1(KEYINPUT31), .A2(G11), .ZN(new_n733));
  NAND2_X1  g308(.A1(KEYINPUT31), .A2(G11), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n731), .A2(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n732), .A2(G33), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT25), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n474), .A2(G139), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n463), .A2(G127), .ZN(new_n743));
  NAND2_X1  g318(.A1(G115), .A2(G2104), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n465), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n736), .B1(new_n746), .B2(new_n732), .ZN(new_n747));
  OAI221_X1 g322(.A(new_n735), .B1(new_n732), .B2(new_n636), .C1(new_n747), .C2(G2072), .ZN(new_n748));
  INV_X1    g323(.A(G2078), .ZN(new_n749));
  NAND2_X1  g324(.A1(G164), .A2(G29), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G27), .B2(G29), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n748), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n732), .A2(G32), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n467), .A2(G105), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT90), .Z(new_n755));
  INV_X1    g330(.A(G141), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n469), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT91), .B(KEYINPUT26), .Z(new_n758));
  NAND3_X1  g333(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n476), .A2(G129), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n753), .B1(new_n763), .B2(new_n732), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT27), .B(G1996), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(G160), .A2(G29), .ZN(new_n767));
  AND2_X1   g342(.A1(KEYINPUT24), .A2(G34), .ZN(new_n768));
  NOR2_X1   g343(.A1(KEYINPUT24), .A2(G34), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n732), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT88), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G2084), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n772), .A2(new_n773), .B1(new_n747), .B2(G2072), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n752), .A2(new_n766), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n772), .A2(new_n773), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT89), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n695), .A2(G21), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G168), .B2(new_n695), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(G1966), .Z(new_n780));
  NAND2_X1  g355(.A1(new_n732), .A2(G35), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G162), .B2(new_n732), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT29), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n780), .B1(new_n783), .B2(G2090), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n474), .A2(G140), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n476), .A2(G128), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n465), .A2(G116), .ZN(new_n787));
  OAI21_X1  g362(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n785), .B(new_n786), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G29), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n732), .A2(G26), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT87), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT28), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(G2067), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n749), .B2(new_n751), .ZN(new_n797));
  NOR4_X1   g372(.A1(new_n775), .A2(new_n777), .A3(new_n784), .A4(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(G171), .A2(new_n695), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G5), .B2(new_n695), .ZN(new_n800));
  INV_X1    g375(.A(G1961), .ZN(new_n801));
  AOI22_X1  g376(.A1(G2090), .A2(new_n783), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n801), .B2(new_n800), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT92), .B(KEYINPUT23), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT93), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n695), .A2(G20), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n805), .B(new_n806), .Z(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n566), .B2(new_n695), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT94), .B(G1956), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n803), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(G4), .A2(G16), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n613), .B2(G16), .ZN(new_n813));
  INV_X1    g388(.A(G1348), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n730), .A2(new_n798), .A3(new_n811), .A4(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n726), .A2(new_n816), .ZN(G311));
  INV_X1    g392(.A(G311), .ZN(G150));
  NAND2_X1  g393(.A1(new_n613), .A2(G559), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT38), .ZN(new_n820));
  INV_X1    g395(.A(G67), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n525), .B2(new_n494), .ZN(new_n822));
  AND2_X1   g397(.A1(G80), .A2(G543), .ZN(new_n823));
  OAI21_X1  g398(.A(G651), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT95), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g401(.A(KEYINPUT95), .B(G651), .C1(new_n822), .C2(new_n823), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n499), .A2(G93), .A3(new_n507), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n505), .A2(G55), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n826), .A2(new_n827), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n549), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n537), .A2(new_n538), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT71), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(new_n539), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n830), .B1(new_n824), .B2(new_n825), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n543), .A2(KEYINPUT70), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n547), .B1(new_n546), .B2(new_n542), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n839), .A2(new_n840), .A3(G651), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n837), .A2(new_n838), .A3(new_n841), .A4(new_n827), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n833), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n820), .B(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT39), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT96), .ZN(new_n847));
  AOI21_X1  g422(.A(G860), .B1(new_n844), .B2(new_n845), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n832), .A2(G860), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT37), .Z(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(G145));
  NAND2_X1  g427(.A1(new_n474), .A2(G142), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n476), .A2(G130), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n465), .A2(G118), .ZN(new_n855));
  OAI21_X1  g430(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n853), .B(new_n854), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n627), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n719), .ZN(new_n859));
  INV_X1    g434(.A(new_n763), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n490), .A2(new_n789), .ZN(new_n861));
  INV_X1    g436(.A(new_n746), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n490), .A2(new_n789), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n862), .B1(new_n861), .B2(new_n863), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n860), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n866), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n868), .A2(new_n763), .A3(new_n864), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n859), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n867), .A2(new_n869), .A3(new_n859), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n871), .A2(KEYINPUT97), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT97), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n867), .A2(new_n869), .A3(new_n874), .A4(new_n859), .ZN(new_n875));
  XNOR2_X1  g450(.A(G160), .B(new_n636), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(G162), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(G37), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT98), .ZN(new_n880));
  INV_X1    g455(.A(new_n877), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n872), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n880), .B1(new_n882), .B2(new_n870), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n871), .A2(KEYINPUT98), .A3(new_n881), .A4(new_n872), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n879), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT99), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT99), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n879), .A2(new_n885), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT40), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT40), .B1(new_n887), .B2(new_n889), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(G395));
  XNOR2_X1  g469(.A(new_n623), .B(new_n843), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n571), .A2(G92), .A3(new_n572), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT10), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n610), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n899), .A2(new_n566), .A3(new_n607), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n566), .B1(new_n899), .B2(new_n607), .ZN(new_n901));
  NOR3_X1   g476(.A1(new_n900), .A2(new_n901), .A3(KEYINPUT41), .ZN(new_n902));
  XOR2_X1   g477(.A(KEYINPUT100), .B(KEYINPUT41), .Z(new_n903));
  NAND2_X1  g478(.A1(new_n612), .A2(G299), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n899), .A2(new_n566), .A3(new_n607), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n895), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n900), .A2(new_n901), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n908), .B1(new_n909), .B2(new_n895), .ZN(new_n910));
  INV_X1    g485(.A(G166), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n586), .A2(new_n911), .A3(new_n589), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n583), .A2(new_n585), .ZN(new_n913));
  OAI21_X1  g488(.A(G166), .B1(new_n913), .B2(new_n588), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(G290), .A2(G288), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n598), .A2(new_n573), .A3(new_n580), .A4(new_n599), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n917), .B1(new_n916), .B2(new_n918), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n915), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n912), .A2(new_n914), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n916), .A2(new_n918), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n922), .B1(new_n923), .B2(new_n917), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT103), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n925), .A2(KEYINPUT42), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n926), .A2(new_n931), .A3(new_n927), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n929), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n910), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n910), .A2(new_n933), .ZN(new_n935));
  OAI21_X1  g510(.A(G868), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n832), .A2(new_n601), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(G295));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n937), .ZN(G331));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n940));
  AND3_X1   g515(.A1(G286), .A2(new_n528), .A3(new_n535), .ZN(new_n941));
  AOI21_X1  g516(.A(G286), .B1(new_n528), .B2(new_n535), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n833), .A2(new_n842), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n943), .B1(new_n833), .B2(new_n842), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n904), .A2(new_n905), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n940), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n946), .B1(new_n902), .B2(new_n906), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n909), .B(KEYINPUT105), .C1(new_n944), .C2(new_n945), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n948), .A2(new_n949), .A3(new_n925), .A4(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G37), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT41), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(new_n900), .B2(new_n901), .ZN(new_n955));
  INV_X1    g530(.A(new_n903), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n904), .A2(new_n905), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n945), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n833), .A2(new_n842), .A3(new_n943), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n955), .A2(new_n957), .A3(new_n958), .A4(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n909), .B1(new_n944), .B2(new_n945), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n946), .A2(KEYINPUT106), .A3(new_n957), .A4(new_n955), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n926), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n953), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT43), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n968), .B1(new_n969), .B2(new_n926), .ZN(new_n970));
  AOI22_X1  g545(.A1(new_n967), .A2(new_n968), .B1(new_n953), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n969), .A2(new_n926), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n974), .A2(new_n968), .A3(new_n952), .A4(new_n951), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT107), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT107), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n953), .A2(new_n977), .A3(new_n968), .A4(new_n974), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n980), .B1(new_n967), .B2(KEYINPUT43), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n979), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n982), .B1(new_n979), .B2(new_n981), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n973), .B1(new_n983), .B2(new_n984), .ZN(G397));
  INV_X1    g560(.A(G1384), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT45), .B1(new_n490), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G40), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n466), .A2(new_n471), .A3(new_n988), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G1996), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n992), .B(KEYINPUT109), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n990), .B(KEYINPUT110), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n763), .A2(new_n991), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n789), .B(G2067), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n993), .A2(new_n763), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n719), .A2(new_n722), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n719), .A2(new_n722), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n994), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  OR2_X1    g577(.A1(G290), .A2(G1986), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  AND2_X1   g579(.A1(G290), .A2(G1986), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n990), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n1007), .B(KEYINPUT111), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n471), .A2(new_n988), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(new_n465), .B2(new_n464), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n987), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n490), .A2(KEYINPUT45), .A3(new_n986), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(new_n749), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1012), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n1016), .A2(new_n1010), .A3(new_n987), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1014), .A2(G2078), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n490), .A2(new_n986), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT50), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n490), .A2(new_n1022), .A3(new_n986), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1021), .A2(new_n1023), .A3(new_n989), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n801), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1015), .A2(new_n1019), .A3(G301), .A4(new_n1025), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1026), .A2(KEYINPUT54), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT126), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1015), .A2(new_n1025), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1012), .A2(new_n1018), .ZN(new_n1030));
  INV_X1    g605(.A(new_n464), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n1031), .A2(KEYINPUT124), .ZN(new_n1032));
  OAI21_X1  g607(.A(G2105), .B1(new_n1031), .B2(KEYINPUT124), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1009), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n987), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT125), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT125), .B1(new_n987), .B2(new_n1034), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1030), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1028), .B1(new_n1029), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(G171), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1029), .A2(new_n1028), .A3(new_n1039), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1027), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(G303), .A2(G8), .ZN(new_n1044));
  XNOR2_X1  g619(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(G303), .A2(G8), .A3(new_n1045), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  OAI22_X1  g624(.A1(new_n1017), .A2(G1971), .B1(new_n1024), .B2(G2090), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(G8), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  OR3_X1    g627(.A1(new_n913), .A2(new_n588), .A3(G1981), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n508), .A2(new_n587), .ZN(new_n1054));
  OAI21_X1  g629(.A(G1981), .B1(new_n913), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1053), .A2(KEYINPUT49), .A3(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n989), .A2(new_n986), .A3(new_n490), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1057), .A2(G8), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT49), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1059), .A2(KEYINPUT115), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n1061));
  AOI211_X1 g636(.A(new_n1061), .B(KEYINPUT49), .C1(new_n1053), .C2(new_n1055), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1056), .B(new_n1058), .C1(new_n1060), .C2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1047), .A2(new_n1050), .A3(G8), .A4(new_n1048), .ZN(new_n1064));
  INV_X1    g639(.A(G1976), .ZN(new_n1065));
  NOR2_X1   g640(.A1(G288), .A2(new_n1065), .ZN(new_n1066));
  OR2_X1    g641(.A1(new_n1066), .A2(KEYINPUT113), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(KEYINPUT113), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(new_n1058), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT52), .B1(G288), .B2(new_n1065), .ZN(new_n1072));
  XOR2_X1   g647(.A(new_n1072), .B(KEYINPUT114), .Z(new_n1073));
  OAI21_X1  g648(.A(new_n1071), .B1(new_n1069), .B2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1052), .A2(new_n1063), .A3(new_n1064), .A4(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1029), .ZN(new_n1078));
  AOI21_X1  g653(.A(G301), .B1(new_n1078), .B2(new_n1019), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n1029), .A2(G171), .A3(new_n1039), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1077), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  OAI22_X1  g656(.A1(new_n1017), .A2(G1966), .B1(new_n1024), .B2(G2084), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(G8), .ZN(new_n1083));
  NAND2_X1  g658(.A1(G286), .A2(G8), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1083), .B(new_n1084), .C1(new_n1085), .C2(KEYINPUT51), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT51), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1087));
  OAI211_X1 g662(.A(G8), .B(new_n1087), .C1(new_n1082), .C2(G286), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1082), .A2(G8), .A3(G286), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1086), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1043), .A2(new_n1076), .A3(new_n1081), .A4(new_n1090), .ZN(new_n1091));
  OR2_X1    g666(.A1(new_n1057), .A2(KEYINPUT118), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1057), .A2(KEYINPUT118), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(new_n795), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1024), .A2(new_n814), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n1097), .A2(KEYINPUT60), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1095), .A2(KEYINPUT60), .A3(new_n1096), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(new_n613), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1095), .A2(KEYINPUT60), .A3(new_n612), .A4(new_n1096), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1017), .A2(new_n991), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n1104), .B(G1341), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1092), .A2(new_n1093), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT120), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1103), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1107), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1109));
  OAI211_X1 g684(.A(KEYINPUT121), .B(new_n550), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1098), .A2(new_n1102), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT56), .B(G2072), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1017), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(G1956), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1024), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT117), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT57), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(G299), .A2(new_n1118), .A3(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n566), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1117), .A2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1114), .A2(new_n1122), .A3(new_n1123), .A4(new_n1116), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(KEYINPUT122), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1127), .A2(new_n1128), .A3(KEYINPUT61), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT61), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1125), .B(new_n1126), .C1(KEYINPUT122), .C2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1112), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1125), .B1(new_n1097), .B2(new_n612), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n1126), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1091), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1090), .A2(KEYINPUT62), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT62), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1086), .A2(new_n1088), .A3(new_n1139), .A4(new_n1089), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1138), .A2(new_n1079), .A3(new_n1076), .A4(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT63), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1082), .A2(G8), .A3(G168), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1142), .B1(new_n1075), .B2(new_n1143), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1063), .A2(new_n1074), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT116), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1051), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1050), .A2(KEYINPUT116), .A3(G8), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1147), .A2(new_n1049), .A3(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1143), .A2(new_n1142), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1145), .A2(new_n1149), .A3(new_n1064), .A4(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1144), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1063), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n573), .A2(new_n1065), .A3(new_n580), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1053), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1064), .ZN(new_n1156));
  AOI22_X1  g731(.A1(new_n1155), .A2(new_n1058), .B1(new_n1156), .B2(new_n1145), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1141), .A2(new_n1152), .A3(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1008), .B1(new_n1137), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n994), .B1(new_n860), .B2(new_n996), .ZN(new_n1160));
  XOR2_X1   g735(.A(new_n992), .B(KEYINPUT109), .Z(new_n1161));
  AND2_X1   g736(.A1(new_n1161), .A2(KEYINPUT46), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1161), .A2(KEYINPUT46), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1160), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1164), .B(KEYINPUT47), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n998), .A2(new_n999), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n789), .A2(G2067), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n994), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1004), .A2(new_n990), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1169), .B(KEYINPUT48), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1002), .A2(new_n1170), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1165), .A2(new_n1168), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1159), .A2(new_n1172), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g748(.A(G229), .ZN(new_n1175));
  OR3_X1    g749(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1176));
  INV_X1    g750(.A(new_n1176), .ZN(new_n1177));
  NAND4_X1  g751(.A1(new_n1175), .A2(new_n890), .A3(new_n971), .A4(new_n1177), .ZN(G225));
  INV_X1    g752(.A(G225), .ZN(G308));
endmodule


