//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n565, new_n567, new_n568, new_n569, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n645, new_n646, new_n649, new_n651, new_n652, new_n653, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206, new_n1207;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT65), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n459), .A2(G101), .A3(G2104), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT69), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n460), .B(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT70), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(G137), .A3(new_n459), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n462), .A2(new_n463), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n463), .B1(new_n462), .B2(new_n469), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  INV_X1    g048(.A(new_n467), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(KEYINPUT66), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT66), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n466), .A2(new_n477), .A3(new_n467), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n476), .A2(G125), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT67), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n473), .B1(new_n482), .B2(G2105), .ZN(new_n483));
  AOI211_X1 g058(.A(KEYINPUT68), .B(new_n459), .C1(new_n479), .C2(new_n481), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n472), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G160));
  NAND2_X1  g061(.A1(new_n468), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT71), .B1(G100), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NOR3_X1   g066(.A1(KEYINPUT71), .A2(G100), .A3(G2105), .ZN(new_n492));
  OAI221_X1 g067(.A(G2104), .B1(G112), .B2(new_n459), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G136), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n468), .A2(new_n459), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n489), .B(new_n493), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G162));
  INV_X1    g072(.A(G126), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n459), .A2(G114), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  OAI22_X1  g075(.A1(new_n487), .A2(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G138), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT72), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n506));
  AOI211_X1 g081(.A(new_n502), .B(G2105), .C1(new_n504), .C2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(new_n476), .A3(new_n478), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT4), .B1(new_n495), .B2(new_n502), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n501), .B1(new_n508), .B2(new_n509), .ZN(G164));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  OAI21_X1  g099(.A(G543), .B1(new_n521), .B2(new_n522), .ZN(new_n525));
  INV_X1    g100(.A(G50), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n523), .A2(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n518), .A2(new_n527), .ZN(G166));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT73), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g106(.A(KEYINPUT73), .B(G543), .C1(new_n521), .C2(new_n522), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT7), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n536), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g113(.A(G63), .B(G651), .C1(new_n520), .C2(new_n519), .ZN(new_n539));
  INV_X1    g114(.A(G89), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n538), .B(new_n539), .C1(new_n523), .C2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n533), .A2(new_n541), .ZN(G168));
  AOI22_X1  g117(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G90), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n543), .A2(new_n517), .B1(new_n544), .B2(new_n523), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT74), .B(G52), .Z(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n547), .B1(new_n531), .B2(new_n532), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(G171));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n550), .B1(new_n531), .B2(new_n532), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n520), .A2(new_n519), .ZN(new_n554));
  INV_X1    g129(.A(G56), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OR2_X1    g131(.A1(KEYINPUT6), .A2(G651), .ZN(new_n557));
  NAND2_X1  g132(.A1(KEYINPUT6), .A2(G651), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n557), .A2(new_n558), .B1(new_n513), .B2(new_n514), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n556), .A2(G651), .B1(new_n559), .B2(G81), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n552), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(G860), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT75), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT76), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(new_n569));
  XOR2_X1   g144(.A(new_n569), .B(KEYINPUT77), .Z(G188));
  INV_X1    g145(.A(G53), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT9), .B1(new_n525), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n557), .A2(new_n558), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n573), .A2(new_n574), .A3(G53), .A4(G543), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n572), .A2(new_n575), .B1(G91), .B2(new_n559), .ZN(new_n576));
  INV_X1    g151(.A(G65), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT78), .B1(new_n520), .B2(new_n519), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n513), .A2(new_n579), .A3(new_n514), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n577), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  AND2_X1   g156(.A1(G78), .A2(G543), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n576), .A2(new_n583), .ZN(G299));
  NAND2_X1  g159(.A1(G77), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G64), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n554), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n587), .A2(G651), .B1(new_n559), .B2(G90), .ZN(new_n588));
  AOI21_X1  g163(.A(KEYINPUT73), .B1(new_n573), .B2(G543), .ZN(new_n589));
  INV_X1    g164(.A(new_n532), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n546), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n588), .A2(new_n591), .ZN(G301));
  INV_X1    g167(.A(KEYINPUT79), .ZN(new_n593));
  INV_X1    g168(.A(new_n541), .ZN(new_n594));
  OAI21_X1  g169(.A(G51), .B1(new_n589), .B2(new_n590), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NOR3_X1   g171(.A1(new_n533), .A2(new_n541), .A3(KEYINPUT79), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n596), .A2(new_n597), .ZN(G286));
  INV_X1    g173(.A(G166), .ZN(G303));
  INV_X1    g174(.A(new_n525), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G49), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n559), .A2(G87), .ZN(new_n602));
  OAI21_X1  g177(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(G288));
  NAND2_X1  g179(.A1(G73), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G61), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n554), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G651), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(KEYINPUT80), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n515), .A2(G61), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n517), .B1(new_n610), .B2(new_n605), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT80), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(G86), .ZN(new_n614));
  INV_X1    g189(.A(G48), .ZN(new_n615));
  OAI22_X1  g190(.A1(new_n523), .A2(new_n614), .B1(new_n525), .B2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n609), .A2(new_n613), .A3(new_n617), .ZN(G305));
  NAND2_X1  g193(.A1(new_n531), .A2(new_n532), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G47), .ZN(new_n620));
  NAND2_X1  g195(.A1(G72), .A2(G543), .ZN(new_n621));
  INV_X1    g196(.A(G60), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n554), .B2(new_n622), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n623), .A2(G651), .B1(new_n559), .B2(G85), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(KEYINPUT81), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT81), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n620), .A2(new_n624), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n628), .ZN(G290));
  NAND2_X1  g204(.A1(G301), .A2(G868), .ZN(new_n630));
  INV_X1    g205(.A(G66), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n631), .B1(new_n578), .B2(new_n580), .ZN(new_n632));
  AND2_X1   g207(.A1(G79), .A2(G543), .ZN(new_n633));
  OAI21_X1  g208(.A(G651), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT10), .ZN(new_n635));
  INV_X1    g210(.A(G92), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n523), .B2(new_n636), .ZN(new_n637));
  NAND4_X1  g212(.A1(new_n573), .A2(new_n515), .A3(KEYINPUT10), .A4(G92), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(G54), .B1(new_n589), .B2(new_n590), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n634), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n630), .B1(new_n642), .B2(G868), .ZN(G284));
  OAI21_X1  g218(.A(new_n630), .B1(new_n642), .B2(G868), .ZN(G321));
  NOR2_X1   g219(.A1(G299), .A2(G868), .ZN(new_n645));
  INV_X1    g220(.A(G286), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n645), .B1(new_n646), .B2(G868), .ZN(G280));
  XOR2_X1   g222(.A(G280), .B(KEYINPUT82), .Z(G297));
  INV_X1    g223(.A(G559), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n642), .B1(new_n649), .B2(G860), .ZN(G148));
  NAND2_X1  g225(.A1(new_n642), .A2(new_n649), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(G868), .ZN(new_n652));
  INV_X1    g227(.A(new_n561), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n652), .B1(G868), .B2(new_n653), .ZN(G323));
  XNOR2_X1  g229(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g230(.A1(new_n465), .A2(G2105), .ZN(new_n656));
  AND3_X1   g231(.A1(new_n476), .A2(new_n656), .A3(new_n478), .ZN(new_n657));
  INV_X1    g232(.A(KEYINPUT12), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT13), .ZN(new_n662));
  INV_X1    g237(.A(G2100), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  INV_X1    g240(.A(new_n495), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(G135), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n488), .A2(G123), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n459), .A2(G111), .ZN(new_n669));
  OAI21_X1  g244(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n667), .B(new_n668), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(G2096), .Z(new_n672));
  NAND3_X1  g247(.A1(new_n664), .A2(new_n665), .A3(new_n672), .ZN(G156));
  INV_X1    g248(.A(KEYINPUT14), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2427), .B(G2438), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2430), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT15), .B(G2435), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n674), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(new_n677), .B2(new_n676), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2451), .B(G2454), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT16), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1341), .B(G1348), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n679), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G2443), .B(G2446), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G14), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n684), .A2(new_n685), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(G401));
  XOR2_X1   g264(.A(G2072), .B(G2078), .Z(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT17), .Z(new_n691));
  XNOR2_X1  g266(.A(G2067), .B(G2678), .ZN(new_n692));
  XOR2_X1   g267(.A(G2084), .B(G2090), .Z(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  NOR3_X1   g269(.A1(new_n691), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT83), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n691), .A2(new_n692), .ZN(new_n697));
  INV_X1    g272(.A(new_n690), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n697), .B(new_n694), .C1(new_n698), .C2(new_n692), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n698), .A2(new_n692), .A3(new_n693), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT18), .Z(new_n701));
  NAND3_X1  g276(.A1(new_n696), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G2096), .B(G2100), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(G227));
  XOR2_X1   g280(.A(G1971), .B(G1976), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT19), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1956), .B(G2474), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1961), .B(G1966), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  NOR3_X1   g286(.A1(new_n707), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n707), .A2(new_n710), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT20), .Z(new_n714));
  AOI211_X1 g289(.A(new_n712), .B(new_n714), .C1(new_n707), .C2(new_n711), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(G1991), .B(G1996), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(G1981), .B(G1986), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(G229));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G25), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n666), .A2(G131), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n488), .A2(G119), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n459), .A2(G107), .ZN(new_n726));
  OAI21_X1  g301(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n724), .B(new_n725), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT84), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n723), .B1(new_n730), .B2(new_n722), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT35), .B(G1991), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G1986), .ZN(new_n734));
  INV_X1    g309(.A(G16), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n735), .A2(G24), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G290), .B2(G16), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n733), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n734), .B2(new_n737), .ZN(new_n739));
  INV_X1    g314(.A(G305), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n740), .A2(new_n735), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G6), .B2(new_n735), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT32), .B(G1981), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n735), .A2(G23), .ZN(new_n744));
  INV_X1    g319(.A(G288), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(new_n735), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT33), .B(G1976), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT85), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n742), .A2(new_n743), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n749), .B2(new_n748), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n735), .A2(G22), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G166), .B2(new_n735), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(G1971), .Z(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n742), .B2(new_n743), .ZN(new_n755));
  OAI21_X1  g330(.A(KEYINPUT34), .B1(new_n751), .B2(new_n755), .ZN(new_n756));
  OR3_X1    g331(.A1(new_n751), .A2(KEYINPUT34), .A3(new_n755), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n739), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT36), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n735), .A2(G20), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT23), .Z(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G299), .B2(G16), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1956), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n722), .A2(G35), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G162), .B2(new_n722), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT29), .Z(new_n766));
  INV_X1    g341(.A(G2090), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n763), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT95), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n722), .A2(G26), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT28), .ZN(new_n771));
  AOI22_X1  g346(.A1(G128), .A2(new_n488), .B1(new_n666), .B2(G140), .ZN(new_n772));
  INV_X1    g347(.A(G104), .ZN(new_n773));
  AND3_X1   g348(.A1(new_n773), .A2(new_n459), .A3(KEYINPUT87), .ZN(new_n774));
  AOI21_X1  g349(.A(KEYINPUT87), .B1(new_n773), .B2(new_n459), .ZN(new_n775));
  OAI221_X1 g350(.A(G2104), .B1(G116), .B2(new_n459), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n777), .A2(KEYINPUT88), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(KEYINPUT88), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n780), .A2(G29), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n781), .A2(KEYINPUT89), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n781), .A2(KEYINPUT89), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n771), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G2067), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n722), .A2(G32), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n666), .A2(G141), .B1(G105), .B2(new_n656), .ZN(new_n788));
  NAND3_X1  g363(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT26), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n488), .B2(G129), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n787), .B1(new_n793), .B2(new_n722), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT27), .ZN(new_n795));
  INV_X1    g370(.A(G1996), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n653), .A2(G16), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G16), .B2(G19), .ZN(new_n799));
  INV_X1    g374(.A(G1341), .ZN(new_n800));
  NOR2_X1   g375(.A1(G5), .A2(G16), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT93), .Z(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G171), .B2(G16), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n799), .A2(new_n800), .B1(G1961), .B2(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT91), .B(G1966), .ZN(new_n805));
  NAND2_X1  g380(.A1(G168), .A2(G16), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G16), .B2(G21), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n722), .A2(G27), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G164), .B2(new_n722), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT94), .B(G2078), .ZN(new_n810));
  OAI221_X1 g385(.A(new_n804), .B1(new_n805), .B2(new_n807), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  OAI221_X1 g387(.A(new_n812), .B1(G1961), .B2(new_n803), .C1(new_n799), .C2(new_n800), .ZN(new_n813));
  NOR2_X1   g388(.A1(G4), .A2(G16), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT86), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n641), .B2(new_n735), .ZN(new_n816));
  INV_X1    g391(.A(G1348), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NOR4_X1   g393(.A1(new_n797), .A2(new_n811), .A3(new_n813), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n786), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(G29), .A2(G33), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT25), .Z(new_n823));
  INV_X1    g398(.A(G139), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n495), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n476), .A2(G127), .A3(new_n478), .ZN(new_n826));
  NAND2_X1  g401(.A1(G115), .A2(G2104), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n459), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n821), .B1(new_n829), .B2(G29), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n830), .A2(G2072), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT30), .B(G28), .ZN(new_n832));
  OR2_X1    g407(.A1(KEYINPUT31), .A2(G11), .ZN(new_n833));
  NAND2_X1  g408(.A1(KEYINPUT31), .A2(G11), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n832), .A2(new_n722), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n671), .B2(new_n722), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT92), .Z(new_n837));
  AOI211_X1 g412(.A(new_n831), .B(new_n837), .C1(new_n805), .C2(new_n807), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n766), .A2(new_n767), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT24), .ZN(new_n840));
  INV_X1    g415(.A(G34), .ZN(new_n841));
  AOI21_X1  g416(.A(G29), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n840), .B2(new_n841), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(G160), .B2(new_n722), .ZN(new_n844));
  OAI211_X1 g419(.A(new_n838), .B(new_n839), .C1(G2084), .C2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n830), .A2(G2072), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT90), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n844), .A2(G2084), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OR4_X1    g424(.A1(new_n769), .A2(new_n820), .A3(new_n845), .A4(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n759), .A2(new_n850), .ZN(G311));
  INV_X1    g426(.A(G311), .ZN(G150));
  NAND2_X1  g427(.A1(new_n642), .A2(G559), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT38), .ZN(new_n854));
  AOI22_X1  g429(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n855));
  INV_X1    g430(.A(G81), .ZN(new_n856));
  OAI22_X1  g431(.A1(new_n855), .A2(new_n517), .B1(new_n856), .B2(new_n523), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n858));
  INV_X1    g433(.A(G93), .ZN(new_n859));
  OAI22_X1  g434(.A1(new_n858), .A2(new_n517), .B1(new_n859), .B2(new_n523), .ZN(new_n860));
  INV_X1    g435(.A(G55), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n861), .B1(new_n531), .B2(new_n532), .ZN(new_n862));
  OAI22_X1  g437(.A1(new_n551), .A2(new_n857), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(G80), .A2(G543), .ZN(new_n864));
  INV_X1    g439(.A(G67), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n864), .B1(new_n554), .B2(new_n865), .ZN(new_n866));
  AOI22_X1  g441(.A1(new_n866), .A2(G651), .B1(new_n559), .B2(G93), .ZN(new_n867));
  OAI21_X1  g442(.A(G55), .B1(new_n589), .B2(new_n590), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n552), .A2(new_n560), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n863), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n854), .B(new_n871), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n872), .A2(KEYINPUT39), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(KEYINPUT39), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n873), .A2(new_n562), .A3(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n860), .A2(new_n862), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n876), .A2(new_n562), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT37), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT96), .ZN(G145));
  NAND2_X1  g455(.A1(new_n666), .A2(G142), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n488), .A2(G130), .ZN(new_n882));
  OAI21_X1  g457(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n883));
  INV_X1    g458(.A(G118), .ZN(new_n884));
  AOI22_X1  g459(.A1(new_n883), .A2(KEYINPUT98), .B1(new_n884), .B2(G2105), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(KEYINPUT98), .B2(new_n883), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n881), .A2(new_n882), .A3(new_n886), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n887), .A2(new_n659), .A3(new_n660), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n887), .B1(new_n659), .B2(new_n660), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n730), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n730), .A2(new_n890), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n892), .A2(KEYINPUT99), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(KEYINPUT99), .B1(new_n892), .B2(new_n893), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n829), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT97), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(new_n898), .A3(new_n792), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n508), .A2(new_n509), .ZN(new_n900));
  INV_X1    g475(.A(new_n501), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n793), .B1(new_n829), .B2(KEYINPUT97), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n899), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n902), .B1(new_n899), .B2(new_n903), .ZN(new_n905));
  OR3_X1    g480(.A1(new_n904), .A2(new_n905), .A3(new_n780), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n780), .B1(new_n904), .B2(new_n905), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n896), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT100), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n671), .B(new_n496), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(G160), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n896), .A2(new_n908), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(new_n910), .A3(new_n909), .ZN(new_n916));
  AOI21_X1  g491(.A(G37), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n906), .A2(new_n907), .A3(new_n893), .A4(new_n892), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n909), .A2(new_n918), .A3(new_n913), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(KEYINPUT101), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n921), .B(new_n922), .ZN(G395));
  AOI22_X1  g498(.A1(G54), .A2(new_n619), .B1(new_n637), .B2(new_n638), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n924), .A2(new_n583), .A3(new_n576), .A4(new_n634), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n641), .A2(G299), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n925), .A2(new_n926), .A3(KEYINPUT41), .ZN(new_n927));
  AOI21_X1  g502(.A(KEYINPUT41), .B1(new_n925), .B2(new_n926), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n871), .B(new_n651), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n925), .A2(new_n926), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n932), .B1(new_n934), .B2(new_n931), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(KEYINPUT42), .ZN(new_n936));
  NAND2_X1  g511(.A1(G290), .A2(new_n740), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n745), .B(G166), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n626), .A2(G305), .A3(new_n628), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n938), .B1(new_n937), .B2(new_n939), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XOR2_X1   g517(.A(new_n936), .B(new_n942), .Z(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(G868), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n944), .B1(G868), .B2(new_n876), .ZN(G295));
  OAI21_X1  g520(.A(new_n944), .B1(G868), .B2(new_n876), .ZN(G331));
  OAI21_X1  g521(.A(G171), .B1(new_n596), .B2(new_n597), .ZN(new_n947));
  OAI21_X1  g522(.A(G301), .B1(new_n533), .B2(new_n541), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n947), .A2(new_n863), .A3(new_n869), .A4(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n594), .A2(new_n595), .A3(new_n593), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT79), .B1(new_n533), .B2(new_n541), .ZN(new_n951));
  AOI21_X1  g526(.A(G301), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(G171), .A2(G168), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n870), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT104), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n949), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n870), .B(KEYINPUT104), .C1(new_n952), .C2(new_n953), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n956), .A2(new_n929), .A3(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT105), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n956), .A2(new_n929), .A3(KEYINPUT105), .A4(new_n957), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT106), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n949), .A2(new_n954), .A3(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n871), .A2(KEYINPUT106), .A3(new_n947), .A4(new_n948), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n934), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n962), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(G37), .B1(new_n968), .B2(new_n942), .ZN(new_n969));
  XOR2_X1   g544(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n970));
  INV_X1    g545(.A(KEYINPUT107), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n942), .B1(new_n934), .B2(new_n966), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n971), .B1(new_n962), .B2(new_n972), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n962), .A2(new_n972), .A3(new_n971), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n969), .B(new_n970), .C1(new_n973), .C2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT44), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(new_n966), .B2(new_n930), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n964), .A2(new_n929), .A3(KEYINPUT108), .A4(new_n965), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n956), .A2(new_n957), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n934), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n978), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(G37), .B1(new_n982), .B2(new_n942), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT109), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n983), .B(new_n984), .C1(new_n974), .C2(new_n973), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n983), .B1(new_n974), .B2(new_n973), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n986), .B1(new_n987), .B2(KEYINPUT109), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n976), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n969), .B1(new_n973), .B2(new_n974), .ZN(new_n990));
  INV_X1    g565(.A(new_n970), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n983), .B(new_n970), .C1(new_n974), .C2(new_n973), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT44), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT110), .B1(new_n989), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n988), .A2(new_n985), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n975), .A2(KEYINPUT44), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n992), .A2(new_n993), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n998), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n995), .A2(new_n1003), .ZN(G397));
  OAI211_X1 g579(.A(new_n472), .B(G40), .C1(new_n483), .C2(new_n484), .ZN(new_n1005));
  XOR2_X1   g580(.A(KEYINPUT111), .B(G1384), .Z(new_n1006));
  AND2_X1   g581(.A1(new_n902), .A2(new_n1006), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n1005), .A2(new_n1007), .A3(KEYINPUT45), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1008), .A2(G1996), .A3(new_n792), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT112), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n780), .A2(G2067), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n778), .A2(new_n785), .A3(new_n779), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n792), .A2(G1996), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1008), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n1010), .A2(new_n1015), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n730), .A2(new_n732), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n730), .A2(new_n732), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1008), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(G290), .B(G1986), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1020), .B1(new_n1008), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT63), .ZN(new_n1023));
  INV_X1    g598(.A(G1384), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n902), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(G8), .B1(new_n1005), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1976), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT52), .B1(G288), .B2(new_n1028), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1027), .B(new_n1029), .C1(new_n1028), .C2(G288), .ZN(new_n1030));
  NOR2_X1   g605(.A1(G288), .A2(new_n1028), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT52), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n1034));
  NOR3_X1   g609(.A1(G305), .A2(KEYINPUT115), .A3(G1981), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT115), .B1(G305), .B2(G1981), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n611), .B1(new_n1038), .B2(new_n616), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(new_n1038), .B2(new_n616), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n1036), .A2(new_n1037), .B1(G1981), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1034), .B1(new_n1041), .B2(KEYINPUT49), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(G1981), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1037), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1043), .B1(new_n1044), .B2(new_n1035), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT49), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1045), .A2(KEYINPUT117), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1042), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1026), .B1(new_n1041), .B2(KEYINPUT49), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1033), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G8), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n902), .A2(KEYINPUT45), .A3(new_n1006), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT45), .B1(new_n902), .B2(new_n1024), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n1052), .A2(new_n1005), .A3(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT113), .B(G1971), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n902), .A2(new_n1058), .A3(new_n1024), .ZN(new_n1059));
  NAND4_X1  g634(.A1(G160), .A2(G40), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1060));
  OAI22_X1  g635(.A1(new_n1054), .A2(new_n1056), .B1(new_n1060), .B2(G2090), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1051), .B1(new_n1061), .B2(KEYINPUT114), .ZN(new_n1062));
  NAND2_X1  g637(.A1(G303), .A2(G8), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1063), .B(KEYINPUT55), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1005), .A2(new_n1053), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1052), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1059), .A2(new_n1057), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1069), .A2(new_n1005), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1068), .A2(new_n1055), .B1(new_n1070), .B2(new_n767), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT114), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1062), .A2(new_n1065), .A3(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1064), .B1(new_n1071), .B2(new_n1051), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1050), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NOR3_X1   g651(.A1(new_n1069), .A2(new_n1005), .A3(G2084), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n902), .A2(KEYINPUT45), .A3(new_n1024), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1066), .A2(new_n1078), .ZN(new_n1079));
  AOI22_X1  g654(.A1(KEYINPUT118), .A2(new_n1077), .B1(new_n1079), .B2(new_n805), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n1060), .B2(G2084), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(G286), .A2(new_n1051), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1023), .B1(new_n1076), .B2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1074), .A2(KEYINPUT63), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT119), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1065), .B1(new_n1062), .B2(new_n1073), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1047), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT117), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1049), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1088), .B1(new_n1089), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(G8), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1061), .A2(KEYINPUT114), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1064), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1098), .A2(new_n1050), .A3(KEYINPUT119), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1087), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1086), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  AOI211_X1 g677(.A(KEYINPUT120), .B(new_n1087), .C1(new_n1095), .C2(new_n1099), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(G1961), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n1069), .B2(new_n1005), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1106), .B(KEYINPUT123), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1007), .A2(KEYINPUT45), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n482), .A2(G2105), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1110), .A2(G2078), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n472), .A2(G40), .A3(new_n1109), .A4(new_n1111), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1108), .A2(new_n1052), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G2078), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1054), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1113), .B1(new_n1115), .B2(new_n1110), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1107), .A2(new_n1116), .A3(G301), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT54), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1110), .B1(new_n1068), .B2(G2078), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1066), .A2(new_n1078), .A3(new_n1111), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1121), .A2(new_n1122), .A3(new_n1106), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(G171), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1124), .A2(new_n1117), .A3(KEYINPUT124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1077), .A2(KEYINPUT118), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1079), .A2(new_n805), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1082), .A2(new_n1126), .A3(new_n1127), .A4(G168), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(G8), .ZN(new_n1129));
  AOI21_X1  g704(.A(G168), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT51), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT51), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1128), .A2(new_n1132), .A3(G8), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1120), .A2(new_n1125), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(KEYINPUT54), .B1(new_n1123), .B2(G171), .ZN(new_n1135));
  AOI21_X1  g710(.A(G301), .B1(new_n1107), .B2(new_n1116), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1135), .B1(KEYINPUT125), .B2(new_n1136), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n1136), .A2(KEYINPUT125), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1076), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  OR3_X1    g714(.A1(new_n1005), .A2(G2067), .A3(new_n1025), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(KEYINPUT122), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1060), .A2(new_n817), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1140), .A2(KEYINPUT122), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n642), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g720(.A(KEYINPUT56), .B(G2072), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1054), .A2(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g722(.A(KEYINPUT121), .B(G1956), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1060), .A2(new_n1149), .ZN(new_n1150));
  XOR2_X1   g725(.A(G299), .B(KEYINPUT57), .Z(new_n1151));
  AND3_X1   g726(.A1(new_n1147), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1145), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1151), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1066), .A2(new_n796), .A3(new_n1067), .ZN(new_n1156));
  XOR2_X1   g731(.A(KEYINPUT58), .B(G1341), .Z(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(new_n1005), .B2(new_n1025), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n561), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT59), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1159), .B(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT61), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1162), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1151), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1147), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1166), .A2(new_n1167), .A3(KEYINPUT61), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1144), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT60), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .A4(new_n642), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1161), .A2(new_n1163), .A3(new_n1168), .A4(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1169), .A2(new_n641), .A3(new_n1170), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1171), .B1(new_n1174), .B2(new_n1145), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1155), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1134), .A2(new_n1139), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(KEYINPUT62), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT62), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1131), .A2(new_n1180), .A3(new_n1133), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1076), .A2(new_n1124), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1179), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1094), .A2(new_n1074), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1092), .A2(new_n1028), .A3(new_n745), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1185), .B1(new_n1044), .B2(new_n1035), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1184), .B1(new_n1186), .B2(new_n1027), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1177), .A2(new_n1183), .A3(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1022), .B1(new_n1104), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1008), .ZN(new_n1190));
  NOR3_X1   g765(.A1(new_n1190), .A2(G1986), .A3(G290), .ZN(new_n1191));
  XNOR2_X1  g766(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1191), .B(new_n1192), .ZN(new_n1193));
  AND3_X1   g768(.A1(new_n1016), .A2(new_n1019), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1190), .B1(new_n1195), .B2(new_n1012), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1008), .B1(new_n1013), .B2(new_n792), .ZN(new_n1197));
  XOR2_X1   g772(.A(new_n1197), .B(KEYINPUT126), .Z(new_n1198));
  NAND2_X1  g773(.A1(new_n1008), .A2(new_n796), .ZN(new_n1199));
  XOR2_X1   g774(.A(new_n1199), .B(KEYINPUT46), .Z(new_n1200));
  OAI21_X1  g775(.A(KEYINPUT47), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1201));
  OR3_X1    g776(.A1(new_n1198), .A2(KEYINPUT47), .A3(new_n1200), .ZN(new_n1202));
  AOI211_X1 g777(.A(new_n1194), .B(new_n1196), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1189), .A2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g779(.A1(new_n704), .A2(G319), .ZN(new_n1206));
  NOR3_X1   g780(.A1(G229), .A2(G401), .A3(new_n1206), .ZN(new_n1207));
  NAND3_X1  g781(.A1(new_n1207), .A2(new_n921), .A3(new_n999), .ZN(G225));
  INV_X1    g782(.A(G225), .ZN(G308));
endmodule


