//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n799,
    new_n800, new_n802, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n980, new_n981, new_n982, new_n983, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009, new_n1010;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT12), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208));
  INV_X1    g007(.A(G1gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT16), .ZN(new_n210));
  AND2_X1   g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n208), .A2(G1gat), .ZN(new_n212));
  OAI21_X1  g011(.A(G8gat), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n208), .A2(new_n210), .ZN(new_n214));
  INV_X1    g013(.A(G8gat), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n214), .B(new_n215), .C1(G1gat), .C2(new_n208), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G43gat), .A2(G50gat), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(G43gat), .A2(G50gat), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT91), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G43gat), .ZN(new_n222));
  INV_X1    g021(.A(G50gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT91), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n224), .A2(new_n225), .A3(new_n218), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n221), .A2(new_n226), .A3(KEYINPUT15), .ZN(new_n227));
  NAND2_X1  g026(.A1(G29gat), .A2(G36gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT14), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n229), .B(KEYINPUT92), .C1(G29gat), .C2(G36gat), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT92), .B1(G29gat), .B2(G36gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT14), .ZN(new_n232));
  NOR3_X1   g031(.A1(KEYINPUT92), .A2(G29gat), .A3(G36gat), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n228), .B(new_n230), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n224), .A2(new_n218), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT93), .B(KEYINPUT15), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n227), .B1(new_n234), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT15), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n239), .B1(new_n235), .B2(KEYINPUT91), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n230), .A2(new_n228), .ZN(new_n241));
  OR3_X1    g040(.A1(KEYINPUT92), .A2(G29gat), .A3(G36gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(KEYINPUT14), .A3(new_n231), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n240), .A2(new_n241), .A3(new_n226), .A4(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n238), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n217), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT17), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n238), .A2(new_n244), .A3(KEYINPUT17), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n246), .B1(new_n250), .B2(new_n217), .ZN(new_n251));
  NAND2_X1  g050(.A1(G229gat), .A2(G233gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT94), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT18), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n238), .A2(new_n244), .A3(KEYINPUT17), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT17), .B1(new_n238), .B2(new_n244), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n217), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n245), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n213), .A2(new_n216), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n257), .A2(KEYINPUT18), .A3(new_n253), .A4(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(new_n253), .B(KEYINPUT13), .Z(new_n262));
  NOR2_X1   g061(.A1(new_n258), .A2(new_n259), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n262), .B1(new_n263), .B2(new_n246), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n207), .B1(new_n254), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n257), .A2(new_n253), .A3(new_n260), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT18), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n269), .A2(new_n206), .A3(new_n264), .A4(new_n261), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(G225gat), .A2(G233gat), .ZN(new_n273));
  XOR2_X1   g072(.A(KEYINPUT79), .B(KEYINPUT5), .Z(new_n274));
  XOR2_X1   g073(.A(G127gat), .B(G134gat), .Z(new_n275));
  INV_X1    g074(.A(KEYINPUT1), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n276), .B1(G113gat), .B2(G120gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  XOR2_X1   g077(.A(KEYINPUT70), .B(G120gat), .Z(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G113gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n277), .ZN(new_n282));
  INV_X1    g081(.A(G113gat), .ZN(new_n283));
  INV_X1    g082(.A(G120gat), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(new_n275), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT76), .ZN(new_n288));
  NAND2_X1  g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT2), .ZN(new_n290));
  INV_X1    g089(.A(G155gat), .ZN(new_n291));
  INV_X1    g090(.A(G162gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n288), .A2(new_n290), .B1(new_n293), .B2(new_n289), .ZN(new_n294));
  INV_X1    g093(.A(G148gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n295), .A2(G141gat), .ZN(new_n296));
  INV_X1    g095(.A(G141gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(G148gat), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n290), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n297), .A2(G148gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n295), .A2(G141gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AND2_X1   g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n290), .B(new_n303), .C1(new_n306), .C2(new_n288), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n300), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT3), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n287), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT77), .B(KEYINPUT3), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n312), .B1(new_n300), .B2(new_n307), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n273), .B(new_n274), .C1(new_n310), .C2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT78), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n308), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT4), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n278), .A2(new_n280), .B1(new_n285), .B2(new_n275), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n300), .A2(KEYINPUT78), .A3(new_n307), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n317), .A2(new_n318), .A3(new_n319), .A4(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n308), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT4), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT80), .ZN(new_n324));
  AND3_X1   g123(.A1(new_n321), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n324), .B1(new_n321), .B2(new_n323), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n315), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n313), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n328), .B(new_n287), .C1(new_n309), .C2(new_n308), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n317), .A2(KEYINPUT4), .A3(new_n319), .A4(new_n320), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n322), .A2(new_n318), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n329), .A2(new_n330), .A3(new_n331), .A4(new_n273), .ZN(new_n332));
  INV_X1    g131(.A(new_n308), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n287), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n322), .ZN(new_n335));
  INV_X1    g134(.A(new_n273), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n274), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G1gat), .B(G29gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT0), .ZN(new_n340));
  XNOR2_X1  g139(.A(G57gat), .B(G85gat), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n340), .B(new_n341), .Z(new_n342));
  NAND4_X1  g141(.A1(new_n327), .A2(KEYINPUT81), .A3(new_n338), .A4(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT6), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n342), .B1(new_n327), .B2(new_n338), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT81), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n327), .A2(new_n338), .A3(new_n342), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n346), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n348), .B1(new_n351), .B2(KEYINPUT6), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G78gat), .B(G106gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(KEYINPUT31), .B(G50gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  XOR2_X1   g155(.A(new_n356), .B(KEYINPUT83), .Z(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  XOR2_X1   g157(.A(KEYINPUT87), .B(G22gat), .Z(new_n359));
  INV_X1    g158(.A(new_n320), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT78), .B1(new_n300), .B2(new_n307), .ZN(new_n361));
  XNOR2_X1  g160(.A(G197gat), .B(G204gat), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT22), .ZN(new_n363));
  INV_X1    g162(.A(G211gat), .ZN(new_n364));
  INV_X1    g163(.A(G218gat), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G211gat), .B(G218gat), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n368), .A2(new_n362), .A3(new_n366), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT29), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI22_X1  g171(.A1(new_n360), .A2(new_n361), .B1(new_n312), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n370), .A2(new_n371), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n375), .B1(new_n313), .B2(KEYINPUT29), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(G228gat), .ZN(new_n378));
  INV_X1    g177(.A(G233gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT84), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n377), .A2(KEYINPUT84), .A3(new_n381), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n333), .B1(new_n372), .B2(KEYINPUT3), .ZN(new_n386));
  OR2_X1    g185(.A1(new_n386), .A2(KEYINPUT85), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT29), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n328), .A2(KEYINPUT86), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT86), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n390), .B1(new_n313), .B2(KEYINPUT29), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(new_n375), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n381), .B1(new_n386), .B2(KEYINPUT85), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n387), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n359), .B1(new_n385), .B2(new_n394), .ZN(new_n395));
  AND3_X1   g194(.A1(new_n377), .A2(KEYINPUT84), .A3(new_n381), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n359), .B(new_n394), .C1(new_n396), .C2(new_n382), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n358), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n387), .A2(new_n393), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n383), .A2(new_n384), .B1(new_n400), .B2(new_n392), .ZN(new_n401));
  INV_X1    g200(.A(G22gat), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n397), .B(new_n356), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT35), .B1(new_n399), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT27), .ZN(new_n405));
  AOI211_X1 g204(.A(KEYINPUT28), .B(G190gat), .C1(new_n405), .C2(G183gat), .ZN(new_n406));
  AND2_X1   g205(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT68), .B1(new_n409), .B2(KEYINPUT27), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT67), .ZN(new_n411));
  INV_X1    g210(.A(G183gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n413), .A2(KEYINPUT68), .A3(KEYINPUT27), .A4(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n406), .B1(new_n410), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT69), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT26), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(G169gat), .ZN(new_n421));
  INV_X1    g220(.A(G176gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AND2_X1   g222(.A1(KEYINPUT69), .A2(KEYINPUT26), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n420), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(G169gat), .A2(G176gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT64), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT64), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(G169gat), .A3(G176gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n418), .A2(new_n419), .A3(new_n421), .A4(new_n422), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n425), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n405), .A2(G183gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n412), .A2(KEYINPUT27), .ZN(new_n434));
  INV_X1    g233(.A(G190gat), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n436), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n417), .A2(new_n432), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(G226gat), .A2(G233gat), .ZN(new_n439));
  AND3_X1   g238(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n441));
  NOR2_X1   g240(.A1(G183gat), .A2(G190gat), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT23), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n444), .A2(new_n421), .A3(new_n422), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n430), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT65), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n443), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n447), .A2(new_n430), .A3(KEYINPUT65), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT25), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n447), .A2(new_n430), .A3(KEYINPUT25), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n440), .B1(new_n409), .B2(new_n435), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT66), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n441), .B(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n453), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n438), .B(new_n439), .C1(new_n452), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n437), .A2(new_n432), .ZN(new_n459));
  INV_X1    g258(.A(new_n406), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n413), .A2(KEYINPUT27), .A3(new_n414), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT68), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n460), .B1(new_n463), .B2(new_n415), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT25), .ZN(new_n466));
  OR3_X1    g265(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n446), .A2(new_n445), .B1(new_n427), .B2(new_n429), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n467), .B1(new_n468), .B2(KEYINPUT65), .ZN(new_n469));
  INV_X1    g268(.A(new_n451), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n457), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n465), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n439), .A2(new_n388), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n458), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n375), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT74), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n448), .A2(new_n449), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n479), .A2(new_n451), .A3(new_n467), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n457), .B1(new_n480), .B2(new_n466), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n474), .B1(new_n481), .B2(new_n465), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n482), .A2(new_n374), .A3(new_n458), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n477), .A2(new_n478), .A3(new_n483), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n482), .A2(new_n374), .A3(new_n458), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT74), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(G8gat), .B(G36gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(G64gat), .B(G92gat), .ZN(new_n489));
  XOR2_X1   g288(.A(new_n488), .B(new_n489), .Z(new_n490));
  AOI21_X1  g289(.A(KEYINPUT30), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT30), .ZN(new_n492));
  INV_X1    g291(.A(new_n490), .ZN(new_n493));
  AOI211_X1 g292(.A(new_n492), .B(new_n493), .C1(new_n484), .C2(new_n486), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n484), .A2(new_n486), .A3(new_n493), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT75), .ZN(new_n496));
  NOR3_X1   g295(.A1(new_n491), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n487), .A2(KEYINPUT30), .A3(new_n490), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n498), .A2(KEYINPUT75), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n353), .B(new_n404), .C1(new_n497), .C2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n319), .B1(new_n481), .B2(new_n465), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n287), .B(new_n438), .C1(new_n452), .C2(new_n457), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(G227gat), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n504), .A2(new_n379), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT34), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT34), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n503), .A2(new_n509), .A3(new_n506), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n501), .A2(new_n505), .A3(new_n502), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT33), .ZN(new_n513));
  XNOR2_X1  g312(.A(G15gat), .B(G43gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(G71gat), .B(G99gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n512), .B(KEYINPUT32), .C1(new_n513), .C2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n516), .B1(new_n512), .B2(KEYINPUT32), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT71), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n512), .A2(new_n519), .A3(new_n513), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n519), .B1(new_n512), .B2(new_n513), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI211_X1 g321(.A(KEYINPUT73), .B(new_n511), .C1(new_n517), .C2(new_n522), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n522), .A2(new_n511), .A3(new_n517), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n511), .B1(new_n517), .B2(new_n522), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n523), .B1(new_n526), .B2(KEYINPUT73), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT90), .B1(new_n500), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n508), .A2(new_n510), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n512), .A2(KEYINPUT32), .ZN(new_n530));
  INV_X1    g329(.A(new_n516), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n521), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n512), .A2(new_n519), .A3(new_n513), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n517), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n529), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n522), .A2(new_n511), .A3(new_n517), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n537), .A2(KEYINPUT73), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT73), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n374), .B1(new_n482), .B2(new_n458), .ZN(new_n543));
  NOR3_X1   g342(.A1(new_n485), .A2(new_n543), .A3(KEYINPUT74), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n483), .A2(new_n478), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n490), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(new_n492), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n495), .A2(KEYINPUT75), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n547), .A2(new_n548), .A3(new_n498), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n498), .A2(KEYINPUT75), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n352), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT90), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n542), .A2(new_n551), .A3(new_n552), .A4(new_n404), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n399), .A2(new_n403), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n526), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT82), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n494), .A2(new_n496), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n499), .B1(new_n557), .B2(new_n547), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n556), .B1(new_n558), .B2(new_n352), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n549), .A2(new_n550), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n560), .A2(KEYINPUT82), .A3(new_n353), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n555), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT35), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n528), .B(new_n553), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n554), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n559), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT36), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n539), .A2(new_n567), .A3(new_n541), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n537), .A2(KEYINPUT72), .A3(KEYINPUT36), .A4(new_n538), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n537), .A2(KEYINPUT36), .A3(new_n538), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT72), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n568), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n334), .A2(new_n322), .A3(new_n273), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n574), .A2(KEYINPUT39), .ZN(new_n575));
  INV_X1    g374(.A(new_n329), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n321), .A2(new_n323), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT80), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n321), .A2(new_n323), .A3(new_n324), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n576), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n575), .B1(new_n580), .B2(new_n273), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n329), .B1(new_n325), .B2(new_n326), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT88), .B(KEYINPUT39), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n582), .A2(new_n336), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n581), .A2(new_n342), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT40), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n581), .A2(KEYINPUT40), .A3(new_n342), .A4(new_n584), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n588), .A2(new_n347), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n549), .A2(new_n550), .A3(new_n587), .A4(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT38), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT37), .B1(new_n484), .B2(new_n486), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT89), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT37), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n487), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n595), .A2(new_n490), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n591), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n594), .B1(new_n477), .B2(new_n483), .ZN(new_n598));
  NOR3_X1   g397(.A1(new_n598), .A2(KEYINPUT38), .A3(new_n490), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT89), .B1(new_n487), .B2(new_n594), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT89), .ZN(new_n601));
  AOI211_X1 g400(.A(new_n601), .B(KEYINPUT37), .C1(new_n484), .C2(new_n486), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n599), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n603), .A2(new_n352), .A3(new_n546), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n590), .B(new_n554), .C1(new_n597), .C2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n566), .A2(new_n573), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n272), .B1(new_n564), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(G64gat), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n608), .A2(G57gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(G57gat), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT9), .ZN(new_n611));
  NAND2_X1  g410(.A1(G71gat), .A2(G78gat), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n609), .A2(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(G71gat), .A2(G78gat), .ZN(new_n614));
  NOR2_X1   g413(.A1(G71gat), .A2(G78gat), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n609), .A2(new_n610), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n618), .B1(KEYINPUT9), .B2(new_n614), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT96), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT95), .ZN(new_n621));
  INV_X1    g420(.A(G71gat), .ZN(new_n622));
  INV_X1    g421(.A(G78gat), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(KEYINPUT95), .B1(G71gat), .B2(G78gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n620), .B1(new_n626), .B2(new_n612), .ZN(new_n627));
  AOI211_X1 g426(.A(KEYINPUT96), .B(new_n614), .C1(new_n624), .C2(new_n625), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n619), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT97), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI211_X1 g430(.A(KEYINPUT97), .B(new_n619), .C1(new_n627), .C2(new_n628), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n617), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n259), .B1(new_n633), .B2(KEYINPUT21), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(KEYINPUT21), .ZN(new_n635));
  NAND2_X1  g434(.A1(G231gat), .A2(G233gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(G127gat), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n637), .A2(G127gat), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n634), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n640), .ZN(new_n642));
  INV_X1    g441(.A(new_n634), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n642), .A2(new_n643), .A3(new_n638), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(new_n291), .ZN(new_n646));
  XNOR2_X1  g445(.A(G183gat), .B(G211gat), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n646), .B(new_n647), .Z(new_n648));
  AND3_X1   g447(.A1(new_n641), .A2(new_n644), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n648), .B1(new_n641), .B2(new_n644), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(G85gat), .A2(G92gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT7), .ZN(new_n653));
  NOR2_X1   g452(.A1(G85gat), .A2(G92gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(G99gat), .A2(G106gat), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n654), .B1(KEYINPUT8), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(G99gat), .B(G106gat), .Z(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n658), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n660), .A2(new_n653), .A3(new_n656), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n250), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n662), .ZN(new_n664));
  AND2_X1   g463(.A1(G232gat), .A2(G233gat), .ZN(new_n665));
  AOI22_X1  g464(.A1(new_n258), .A2(new_n664), .B1(KEYINPUT41), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(KEYINPUT102), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT102), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n663), .A2(new_n669), .A3(new_n666), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT101), .B(G190gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(G218gat), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n668), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n672), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n663), .A2(new_n669), .A3(new_n666), .A4(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT100), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n665), .A2(KEYINPUT41), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT98), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n679), .B(KEYINPUT99), .Z(new_n680));
  XOR2_X1   g479(.A(G134gat), .B(G162gat), .Z(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n673), .A2(new_n677), .A3(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n682), .B1(new_n673), .B2(new_n677), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(G230gat), .A2(G233gat), .ZN(new_n688));
  INV_X1    g487(.A(new_n625), .ZN(new_n689));
  NOR3_X1   g488(.A1(KEYINPUT95), .A2(G71gat), .A3(G78gat), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n612), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT96), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n626), .A2(new_n620), .A3(new_n612), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(KEYINPUT97), .B1(new_n694), .B2(new_n619), .ZN(new_n695));
  INV_X1    g494(.A(new_n632), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n616), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n662), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n633), .A2(new_n664), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n688), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT103), .B(KEYINPUT10), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n698), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  AOI211_X1 g501(.A(new_n617), .B(new_n662), .C1(new_n631), .C2(new_n632), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(KEYINPUT10), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n700), .B1(new_n705), .B2(new_n688), .ZN(new_n706));
  XNOR2_X1  g505(.A(G120gat), .B(G148gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(G176gat), .B(G204gat), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n707), .B(new_n708), .Z(new_n709));
  NAND2_X1  g508(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n709), .ZN(new_n711));
  INV_X1    g510(.A(new_n688), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n712), .B1(new_n702), .B2(new_n704), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n711), .B1(new_n713), .B2(new_n700), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n651), .A2(new_n687), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n607), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(new_n353), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(new_n209), .ZN(G1324gat));
  NOR2_X1   g518(.A1(new_n717), .A2(new_n560), .ZN(new_n720));
  OR2_X1    g519(.A1(new_n720), .A2(KEYINPUT104), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(KEYINPUT104), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n721), .A2(G8gat), .A3(new_n722), .ZN(new_n723));
  XOR2_X1   g522(.A(KEYINPUT16), .B(G8gat), .Z(new_n724));
  NAND3_X1  g523(.A1(new_n720), .A2(KEYINPUT42), .A3(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n724), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n726), .B1(new_n721), .B2(new_n722), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n723), .B(new_n725), .C1(new_n727), .C2(KEYINPUT42), .ZN(G1325gat));
  OAI21_X1  g527(.A(G15gat), .B1(new_n717), .B2(new_n573), .ZN(new_n729));
  OR2_X1    g528(.A1(new_n527), .A2(G15gat), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(new_n717), .B2(new_n730), .ZN(G1326gat));
  AND2_X1   g530(.A1(new_n607), .A2(new_n565), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n716), .ZN(new_n733));
  XNOR2_X1  g532(.A(KEYINPUT43), .B(G22gat), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1327gat));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n736));
  AND3_X1   g535(.A1(new_n559), .A2(new_n561), .A3(new_n565), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n605), .A2(new_n573), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT107), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n566), .A2(new_n740), .A3(new_n573), .A4(new_n605), .ZN(new_n741));
  INV_X1    g540(.A(new_n555), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n551), .A2(KEYINPUT82), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n558), .A2(new_n556), .A3(new_n352), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(KEYINPUT35), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n528), .A2(new_n553), .ZN(new_n747));
  AOI22_X1  g546(.A1(new_n739), .A2(new_n741), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n736), .B1(new_n748), .B2(new_n686), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n564), .A2(new_n606), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n750), .A2(KEYINPUT44), .A3(new_n687), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  XOR2_X1   g551(.A(new_n715), .B(KEYINPUT105), .Z(new_n753));
  NAND3_X1  g552(.A1(new_n651), .A2(new_n753), .A3(new_n271), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n754), .B(KEYINPUT106), .Z(new_n755));
  NAND2_X1  g554(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(G29gat), .B1(new_n756), .B2(new_n353), .ZN(new_n757));
  INV_X1    g556(.A(new_n651), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n758), .A2(new_n686), .A3(new_n715), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n607), .A2(new_n759), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n760), .A2(G29gat), .A3(new_n353), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n761), .B(KEYINPUT45), .Z(new_n762));
  NAND2_X1  g561(.A1(new_n757), .A2(new_n762), .ZN(G1328gat));
  OAI21_X1  g562(.A(G36gat), .B1(new_n756), .B2(new_n560), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n760), .A2(G36gat), .A3(new_n560), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT46), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(G1329gat));
  NOR2_X1   g566(.A1(new_n573), .A2(new_n222), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n749), .A2(new_n751), .A3(new_n755), .A4(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n222), .B1(new_n760), .B2(new_n527), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g571(.A1(new_n749), .A2(new_n565), .A3(new_n751), .A4(new_n755), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(G50gat), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n732), .A2(new_n223), .A3(new_n759), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT48), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n774), .A2(KEYINPUT48), .A3(new_n775), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(G1331gat));
  OAI211_X1 g579(.A(new_n272), .B(new_n686), .C1(new_n649), .C2(new_n650), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(new_n753), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(KEYINPUT108), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n748), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n352), .ZN(new_n785));
  XOR2_X1   g584(.A(KEYINPUT109), .B(G57gat), .Z(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(G1332gat));
  OR2_X1    g586(.A1(new_n748), .A2(new_n783), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT49), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n558), .B1(new_n789), .B2(new_n608), .ZN(new_n790));
  XOR2_X1   g589(.A(new_n790), .B(KEYINPUT110), .Z(new_n791));
  OAI21_X1  g590(.A(KEYINPUT111), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  OR4_X1    g591(.A1(KEYINPUT111), .A2(new_n748), .A3(new_n783), .A4(new_n791), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n794), .B(new_n795), .ZN(G1333gat));
  NAND3_X1  g595(.A1(new_n784), .A2(new_n622), .A3(new_n542), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n788), .A2(new_n573), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n797), .B1(new_n798), .B2(new_n622), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n799), .B(new_n800), .ZN(G1334gat));
  NAND2_X1  g600(.A1(new_n784), .A2(new_n565), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g602(.A1(new_n651), .A2(new_n272), .ZN(new_n804));
  INV_X1    g603(.A(new_n715), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n752), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(G85gat), .B1(new_n807), .B2(new_n353), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n353), .A2(new_n805), .A3(G85gat), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n739), .A2(new_n741), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n686), .B1(new_n810), .B2(new_n564), .ZN(new_n811));
  INV_X1    g610(.A(new_n804), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT51), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT51), .ZN(new_n814));
  NOR4_X1   g613(.A1(new_n748), .A2(new_n814), .A3(new_n686), .A4(new_n804), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n809), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n808), .A2(new_n816), .ZN(G1336gat));
  NAND4_X1  g616(.A1(new_n749), .A2(new_n558), .A3(new_n751), .A4(new_n806), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(G92gat), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n753), .A2(G92gat), .A3(new_n560), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n820), .B1(new_n813), .B2(new_n815), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n819), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT52), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n819), .A2(new_n821), .A3(new_n822), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(G1337gat));
  OAI21_X1  g626(.A(G99gat), .B1(new_n807), .B2(new_n573), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n527), .A2(G99gat), .A3(new_n805), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(new_n813), .B2(new_n815), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(G1338gat));
  NAND4_X1  g630(.A1(new_n749), .A2(new_n565), .A3(new_n751), .A4(new_n806), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(G106gat), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n753), .A2(G106gat), .A3(new_n554), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n834), .B1(new_n813), .B2(new_n815), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(KEYINPUT53), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n833), .A2(new_n835), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(G1339gat));
  NOR2_X1   g639(.A1(new_n781), .A2(new_n715), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n251), .A2(new_n253), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n263), .A2(new_n246), .A3(new_n262), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n205), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n844), .A2(new_n270), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n715), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n633), .A2(new_n664), .ZN(new_n847));
  INV_X1    g646(.A(new_n701), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n847), .A2(new_n703), .A3(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n704), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n688), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n702), .A2(new_n704), .A3(new_n712), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(KEYINPUT54), .A3(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n709), .B1(new_n713), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n853), .A2(new_n855), .A3(KEYINPUT55), .ZN(new_n856));
  AOI22_X1  g655(.A1(new_n706), .A2(new_n709), .B1(new_n266), .B2(new_n270), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT55), .B1(new_n853), .B2(new_n855), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n846), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n686), .ZN(new_n861));
  INV_X1    g660(.A(new_n685), .ZN(new_n862));
  AOI22_X1  g661(.A1(new_n862), .A2(new_n683), .B1(new_n706), .B2(new_n709), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n853), .A2(new_n855), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT55), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n863), .A2(new_n845), .A3(new_n866), .A4(new_n856), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n861), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n758), .B1(new_n868), .B2(KEYINPUT113), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT113), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n861), .A2(new_n870), .A3(new_n867), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n841), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NOR4_X1   g671(.A1(new_n872), .A2(new_n353), .A3(new_n558), .A4(new_n555), .ZN(new_n873));
  AOI21_X1  g672(.A(G113gat), .B1(new_n873), .B2(new_n271), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n872), .A2(new_n565), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n558), .A2(new_n353), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n875), .A2(new_n542), .A3(new_n876), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT114), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n272), .A2(new_n283), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n874), .B1(new_n878), .B2(new_n879), .ZN(G1340gat));
  INV_X1    g679(.A(new_n878), .ZN(new_n881));
  OAI21_X1  g680(.A(G120gat), .B1(new_n881), .B2(new_n753), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n805), .A2(new_n279), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n873), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(G1341gat));
  OAI21_X1  g684(.A(G127gat), .B1(new_n881), .B2(new_n651), .ZN(new_n886));
  INV_X1    g685(.A(G127gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n873), .A2(new_n887), .A3(new_n758), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n888), .ZN(G1342gat));
  OAI21_X1  g688(.A(G134gat), .B1(new_n881), .B2(new_n686), .ZN(new_n890));
  INV_X1    g689(.A(G134gat), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n873), .A2(new_n891), .A3(new_n687), .ZN(new_n892));
  XOR2_X1   g691(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n893));
  XNOR2_X1  g692(.A(new_n892), .B(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n890), .A2(new_n894), .ZN(G1343gat));
  AND2_X1   g694(.A1(new_n573), .A2(new_n876), .ZN(new_n896));
  INV_X1    g695(.A(new_n841), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n866), .A2(new_n856), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n710), .B(new_n845), .C1(new_n684), .C2(new_n685), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g699(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n901), .B1(new_n853), .B2(new_n855), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n846), .B1(new_n858), .B2(new_n902), .ZN(new_n903));
  OR2_X1    g702(.A1(new_n903), .A2(KEYINPUT117), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n687), .B1(new_n903), .B2(KEYINPUT117), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n900), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n897), .B1(new_n906), .B2(new_n758), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n565), .A2(KEYINPUT57), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n866), .A2(new_n856), .A3(new_n857), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n687), .B1(new_n910), .B2(new_n846), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT113), .B1(new_n911), .B2(new_n900), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(new_n651), .A3(new_n871), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n897), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT57), .B1(new_n914), .B2(new_n565), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n896), .B1(new_n909), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(G141gat), .B1(new_n916), .B2(new_n272), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n872), .A2(new_n353), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n573), .A2(new_n565), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n919), .A2(new_n560), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n271), .A2(new_n297), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT118), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n917), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g724(.A(new_n921), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n926), .A2(new_n295), .A3(new_n715), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n715), .B(new_n896), .C1(new_n909), .C2(new_n915), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n295), .A2(KEYINPUT59), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT119), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n930), .B(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT59), .ZN(new_n933));
  AOI21_X1  g732(.A(KEYINPUT57), .B1(new_n907), .B2(new_n565), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n934), .A2(KEYINPUT120), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n914), .A2(new_n908), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n936), .B1(new_n934), .B2(KEYINPUT120), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n715), .B(new_n896), .C1(new_n935), .C2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n933), .B1(new_n938), .B2(G148gat), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n927), .B1(new_n932), .B2(new_n939), .ZN(G1345gat));
  OAI21_X1  g739(.A(G155gat), .B1(new_n916), .B2(new_n651), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n926), .A2(new_n291), .A3(new_n758), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1346gat));
  NOR3_X1   g742(.A1(new_n916), .A2(new_n292), .A3(new_n686), .ZN(new_n944));
  AOI21_X1  g743(.A(G162gat), .B1(new_n926), .B2(new_n687), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n944), .A2(new_n945), .ZN(G1347gat));
  AOI21_X1  g745(.A(new_n352), .B1(new_n913), .B2(new_n897), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT121), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n558), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AOI211_X1 g748(.A(KEYINPUT121), .B(new_n352), .C1(new_n913), .C2(new_n897), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n949), .A2(new_n555), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n951), .A2(new_n421), .A3(new_n271), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n560), .A2(new_n352), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(new_n542), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT122), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n875), .A2(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(new_n271), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n958), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT123), .B1(new_n958), .B2(G169gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n952), .B1(new_n959), .B2(new_n960), .ZN(G1348gat));
  OAI21_X1  g760(.A(G176gat), .B1(new_n956), .B2(new_n753), .ZN(new_n962));
  OAI21_X1  g761(.A(KEYINPUT121), .B1(new_n872), .B2(new_n352), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n914), .A2(new_n948), .A3(new_n353), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n963), .A2(new_n558), .A3(new_n742), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n715), .A2(new_n422), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n962), .B1(new_n965), .B2(new_n966), .ZN(G1349gat));
  OAI22_X1  g766(.A1(new_n956), .A2(new_n651), .B1(new_n408), .B2(new_n407), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT124), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n433), .A2(new_n434), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n651), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n969), .B1(new_n951), .B2(new_n971), .ZN(new_n972));
  INV_X1    g771(.A(new_n971), .ZN(new_n973));
  NOR3_X1   g772(.A1(new_n965), .A2(KEYINPUT124), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n968), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(KEYINPUT60), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT60), .ZN(new_n977));
  OAI211_X1 g776(.A(new_n977), .B(new_n968), .C1(new_n972), .C2(new_n974), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n976), .A2(new_n978), .ZN(G1350gat));
  NAND3_X1  g778(.A1(new_n951), .A2(new_n435), .A3(new_n687), .ZN(new_n980));
  OAI21_X1  g779(.A(G190gat), .B1(new_n956), .B2(new_n686), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n981), .A2(KEYINPUT61), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n981), .A2(KEYINPUT61), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(G1351gat));
  OR2_X1    g783(.A1(new_n935), .A2(new_n937), .ZN(new_n985));
  AND2_X1   g784(.A1(new_n573), .A2(new_n953), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n985), .A2(new_n271), .A3(new_n986), .ZN(new_n987));
  XOR2_X1   g786(.A(KEYINPUT125), .B(G197gat), .Z(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g788(.A1(new_n963), .A2(new_n558), .A3(new_n919), .A4(new_n964), .ZN(new_n990));
  OR2_X1    g789(.A1(new_n272), .A2(new_n988), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(G1352gat));
  INV_X1    g791(.A(new_n753), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n985), .A2(new_n993), .A3(new_n986), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n994), .A2(G204gat), .ZN(new_n995));
  OR2_X1    g794(.A1(new_n805), .A2(G204gat), .ZN(new_n996));
  OAI21_X1  g795(.A(KEYINPUT62), .B1(new_n990), .B2(new_n996), .ZN(new_n997));
  OR3_X1    g796(.A1(new_n990), .A2(KEYINPUT62), .A3(new_n996), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n995), .A2(new_n997), .A3(new_n998), .ZN(G1353gat));
  OAI211_X1 g798(.A(new_n758), .B(new_n986), .C1(new_n935), .C2(new_n937), .ZN(new_n1000));
  OAI21_X1  g799(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n1001));
  INV_X1    g800(.A(new_n1001), .ZN(new_n1002));
  AND2_X1   g801(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n1003));
  AND3_X1   g802(.A1(new_n1000), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g803(.A(new_n1003), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n758), .A2(new_n364), .ZN(new_n1006));
  OAI22_X1  g805(.A1(new_n1004), .A2(new_n1005), .B1(new_n990), .B2(new_n1006), .ZN(G1354gat));
  NAND3_X1  g806(.A1(new_n985), .A2(new_n687), .A3(new_n986), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1008), .A2(G218gat), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n687), .A2(new_n365), .ZN(new_n1010));
  OAI21_X1  g809(.A(new_n1009), .B1(new_n990), .B2(new_n1010), .ZN(G1355gat));
endmodule


