//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 0 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202));
  AND2_X1   g001(.A1(G232gat), .A2(G233gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT41), .ZN(new_n204));
  INV_X1    g003(.A(G50gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G43gat), .ZN(new_n206));
  INV_X1    g005(.A(G43gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G50gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT87), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n206), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT15), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n205), .A2(KEYINPUT87), .A3(G43gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n206), .A2(new_n208), .A3(KEYINPUT15), .ZN(new_n214));
  INV_X1    g013(.A(G29gat), .ZN(new_n215));
  INV_X1    g014(.A(G36gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT14), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT14), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(G29gat), .B2(G36gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(G29gat), .A2(G36gat), .ZN(new_n220));
  AND3_X1   g019(.A1(new_n217), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n213), .A2(new_n214), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT88), .B1(new_n221), .B2(new_n214), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n213), .A2(KEYINPUT88), .A3(new_n214), .A4(new_n221), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT7), .ZN(new_n228));
  INV_X1    g027(.A(G85gat), .ZN(new_n229));
  INV_X1    g028(.A(G92gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G99gat), .A2(G106gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT8), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n229), .A2(new_n230), .ZN(new_n236));
  AND3_X1   g035(.A1(new_n235), .A2(KEYINPUT96), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT96), .B1(new_n235), .B2(new_n236), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n233), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(G99gat), .B(G106gat), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n235), .A2(new_n236), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT96), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n235), .A2(KEYINPUT96), .A3(new_n236), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n240), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(new_n247), .A3(new_n233), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n241), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n204), .B1(new_n227), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT17), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n226), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n224), .A2(KEYINPUT17), .A3(new_n225), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(new_n253), .A3(new_n249), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT97), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n252), .A2(KEYINPUT97), .A3(new_n253), .A4(new_n249), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n250), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G190gat), .B(G218gat), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n202), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(G134gat), .B(G162gat), .Z(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(KEYINPUT95), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n203), .A2(KEYINPUT41), .ZN(new_n264));
  XOR2_X1   g063(.A(new_n263), .B(new_n264), .Z(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n258), .A2(new_n260), .ZN(new_n268));
  AOI211_X1 g067(.A(new_n259), .B(new_n250), .C1(new_n256), .C2(new_n257), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  OAI22_X1  g070(.A1(new_n261), .A2(new_n266), .B1(new_n268), .B2(new_n269), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G64gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(G57gat), .ZN(new_n276));
  INV_X1    g075(.A(G57gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(G64gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT9), .ZN(new_n280));
  INV_X1    g079(.A(G71gat), .ZN(new_n281));
  INV_X1    g080(.A(G78gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(G71gat), .A2(G78gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AND2_X1   g084(.A1(new_n280), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT92), .B1(new_n277), .B2(G64gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT92), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(new_n275), .A3(G57gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n287), .A2(new_n289), .A3(new_n278), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT93), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT93), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n287), .A2(new_n289), .A3(new_n292), .A4(new_n278), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n283), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n284), .A2(KEYINPUT9), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n286), .B1(new_n294), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n298), .A2(KEYINPUT21), .ZN(new_n299));
  XOR2_X1   g098(.A(G127gat), .B(G155gat), .Z(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G1gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT16), .ZN(new_n303));
  INV_X1    g102(.A(G22gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G15gat), .ZN(new_n305));
  INV_X1    g104(.A(G15gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G22gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n303), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G15gat), .B(G22gat), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n308), .B1(G1gat), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G8gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT89), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n312), .B1(new_n309), .B2(G1gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n310), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  OAI221_X1 g113(.A(new_n308), .B1(new_n312), .B2(G8gat), .C1(G1gat), .C2(new_n309), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT90), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n314), .A2(KEYINPUT90), .A3(new_n315), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n320), .B1(KEYINPUT21), .B2(new_n298), .ZN(new_n321));
  XOR2_X1   g120(.A(new_n301), .B(new_n321), .Z(new_n322));
  NAND2_X1  g121(.A1(G231gat), .A2(G233gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n323), .B(KEYINPUT94), .ZN(new_n324));
  XOR2_X1   g123(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G183gat), .B(G211gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n326), .B(new_n327), .ZN(new_n328));
  XOR2_X1   g127(.A(new_n322), .B(new_n328), .Z(new_n329));
  NAND2_X1  g128(.A1(new_n274), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n247), .B1(new_n246), .B2(new_n233), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n231), .A2(new_n232), .ZN(new_n332));
  AOI211_X1 g131(.A(new_n240), .B(new_n332), .C1(new_n244), .C2(new_n245), .ZN(new_n333));
  AOI22_X1  g132(.A1(new_n291), .A2(new_n293), .B1(new_n295), .B2(new_n296), .ZN(new_n334));
  OAI22_X1  g133(.A1(new_n331), .A2(new_n333), .B1(new_n334), .B2(new_n286), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n294), .A2(new_n297), .ZN(new_n336));
  INV_X1    g135(.A(new_n286), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n336), .A2(new_n241), .A3(new_n248), .A4(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G230gat), .A2(G233gat), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT99), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT100), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n339), .A2(KEYINPUT99), .A3(new_n341), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT99), .B1(new_n339), .B2(new_n341), .ZN(new_n348));
  AOI211_X1 g147(.A(new_n343), .B(new_n340), .C1(new_n335), .C2(new_n338), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT100), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT10), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n338), .A3(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n298), .A2(KEYINPUT10), .A3(new_n248), .A4(new_n241), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n341), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G120gat), .B(G148gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(KEYINPUT101), .ZN(new_n356));
  XNOR2_X1  g155(.A(G176gat), .B(G204gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n347), .A2(new_n350), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n346), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n358), .B1(new_n361), .B2(new_n354), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT102), .B1(new_n330), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(G229gat), .A2(G233gat), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n252), .A2(new_n316), .A3(new_n253), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT91), .B1(new_n320), .B2(new_n226), .ZN(new_n367));
  AND3_X1   g166(.A1(new_n314), .A2(KEYINPUT90), .A3(new_n315), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT90), .B1(new_n314), .B2(new_n315), .ZN(new_n369));
  OAI211_X1 g168(.A(KEYINPUT91), .B(new_n226), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n365), .B(new_n366), .C1(new_n367), .C2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT18), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n226), .B1(new_n368), .B2(new_n369), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT91), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n370), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n378), .A2(KEYINPUT18), .A3(new_n365), .A4(new_n366), .ZN(new_n379));
  INV_X1    g178(.A(new_n320), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(new_n227), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n381), .B1(new_n367), .B2(new_n371), .ZN(new_n382));
  XOR2_X1   g181(.A(new_n365), .B(KEYINPUT13), .Z(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n374), .A2(new_n379), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT86), .ZN(new_n386));
  XNOR2_X1  g185(.A(G113gat), .B(G141gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(G197gat), .ZN(new_n388));
  XOR2_X1   g187(.A(KEYINPUT11), .B(G169gat), .Z(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT85), .B(KEYINPUT12), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n390), .B(new_n391), .Z(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n386), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n385), .A2(KEYINPUT86), .A3(new_n392), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT102), .ZN(new_n398));
  INV_X1    g197(.A(new_n363), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n274), .A2(new_n398), .A3(new_n329), .A4(new_n399), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n364), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G15gat), .B(G43gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(G71gat), .B(G99gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(G183gat), .ZN(new_n405));
  INV_X1    g204(.A(G190gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(G183gat), .A2(G190gat), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n407), .A2(KEYINPUT24), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT24), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n410), .A2(G183gat), .A3(G190gat), .ZN(new_n411));
  NOR2_X1   g210(.A1(G169gat), .A2(G176gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT23), .ZN(new_n413));
  NAND2_X1  g212(.A1(G169gat), .A2(G176gat), .ZN(new_n414));
  AND4_X1   g213(.A1(new_n409), .A2(new_n411), .A3(new_n413), .A4(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(G169gat), .ZN(new_n416));
  INV_X1    g215(.A(G176gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT23), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n418), .A2(KEYINPUT64), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT64), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n421), .B1(new_n412), .B2(KEYINPUT23), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT25), .B1(new_n415), .B2(new_n423), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n413), .A2(new_n411), .A3(new_n414), .ZN(new_n425));
  AND4_X1   g224(.A1(KEYINPUT25), .A2(new_n425), .A3(new_n423), .A4(new_n409), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT27), .B(G183gat), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n427), .A2(KEYINPUT28), .A3(new_n406), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT28), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT27), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(G183gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT65), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n406), .B(new_n433), .C1(new_n427), .C2(KEYINPUT65), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n429), .B1(new_n430), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT66), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n436), .B1(new_n418), .B2(KEYINPUT26), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT26), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n412), .A2(KEYINPUT66), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n414), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n441), .B1(KEYINPUT26), .B2(new_n418), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n408), .ZN(new_n444));
  OAI22_X1  g243(.A1(new_n424), .A2(new_n426), .B1(new_n435), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT1), .ZN(new_n446));
  INV_X1    g245(.A(G113gat), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n447), .A2(G120gat), .ZN(new_n448));
  INV_X1    g247(.A(G120gat), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n449), .A2(G113gat), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n446), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(G127gat), .ZN(new_n452));
  INV_X1    g251(.A(G134gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(G127gat), .A2(G134gat), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n454), .A2(new_n455), .B1(KEYINPUT67), .B2(new_n446), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n449), .A2(G113gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n447), .A2(G120gat), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT1), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n446), .A2(KEYINPUT67), .ZN(new_n461));
  INV_X1    g260(.A(new_n455), .ZN(new_n462));
  NOR2_X1   g261(.A1(G127gat), .A2(G134gat), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n457), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n445), .A2(KEYINPUT68), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(G227gat), .ZN(new_n468));
  INV_X1    g267(.A(G233gat), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n425), .A2(new_n423), .A3(new_n409), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT25), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n415), .A2(KEYINPUT25), .A3(new_n423), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n433), .A2(new_n406), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n405), .A2(KEYINPUT27), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT65), .B1(new_n432), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n430), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n428), .ZN(new_n479));
  AOI22_X1  g278(.A1(new_n440), .A2(new_n442), .B1(G183gat), .B2(G190gat), .ZN(new_n480));
  AOI22_X1  g279(.A1(new_n473), .A2(new_n474), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT68), .ZN(new_n482));
  OR2_X1    g281(.A1(new_n466), .A2(KEYINPUT68), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n467), .A2(new_n470), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT33), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n404), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(KEYINPUT32), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n485), .B(KEYINPUT32), .C1(new_n486), .C2(new_n404), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n467), .A2(new_n484), .ZN(new_n493));
  INV_X1    g292(.A(new_n470), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n492), .ZN(new_n496));
  AOI211_X1 g295(.A(new_n470), .B(new_n496), .C1(new_n467), .C2(new_n484), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n491), .A2(KEYINPUT70), .A3(new_n499), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n498), .A2(new_n489), .A3(new_n490), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n498), .B1(new_n489), .B2(new_n490), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT70), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n500), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT76), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT73), .ZN(new_n507));
  INV_X1    g306(.A(G155gat), .ZN(new_n508));
  INV_X1    g307(.A(G162gat), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(G155gat), .A2(G162gat), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT73), .B1(G155gat), .B2(G162gat), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G141gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(G148gat), .ZN(new_n515));
  INV_X1    g314(.A(G148gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(G141gat), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT2), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n516), .A2(KEYINPUT74), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT74), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(G148gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(new_n522), .A3(G141gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT2), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n524), .A2(new_n508), .A3(new_n509), .ZN(new_n525));
  AOI22_X1  g324(.A1(new_n523), .A2(new_n515), .B1(new_n511), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n506), .B1(new_n519), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n523), .A2(new_n515), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n525), .A2(new_n511), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n517), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n524), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n530), .A2(new_n534), .A3(KEYINPUT76), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n527), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G211gat), .B(G218gat), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n537), .A2(KEYINPUT71), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(KEYINPUT71), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G197gat), .B(G204gat), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT22), .ZN(new_n542));
  INV_X1    g341(.A(G211gat), .ZN(new_n543));
  INV_X1    g342(.A(G218gat), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n540), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n538), .A2(new_n545), .A3(new_n541), .A4(new_n539), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT29), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n536), .B1(new_n549), .B2(KEYINPUT3), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n547), .A2(new_n548), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT3), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n530), .A2(new_n534), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT29), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n550), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G228gat), .A2(G233gat), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n559), .B(KEYINPUT82), .Z(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n530), .A2(new_n534), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n562), .B1(new_n549), .B2(KEYINPUT3), .ZN(new_n563));
  INV_X1    g362(.A(new_n559), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n557), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G78gat), .B(G106gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(KEYINPUT31), .B(G50gat), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n567), .B(new_n568), .Z(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT83), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n304), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n569), .B1(new_n561), .B2(new_n565), .ZN(new_n574));
  NOR3_X1   g373(.A1(new_n574), .A2(KEYINPUT83), .A3(G22gat), .ZN(new_n575));
  OAI22_X1  g374(.A1(new_n573), .A2(new_n575), .B1(new_n570), .B2(new_n566), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n571), .A2(new_n572), .A3(new_n304), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n566), .A2(new_n570), .ZN(new_n578));
  OAI21_X1  g377(.A(G22gat), .B1(new_n574), .B2(KEYINPUT83), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n505), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G1gat), .B(G29gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT0), .ZN(new_n584));
  XNOR2_X1  g383(.A(G57gat), .B(G85gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n584), .B(new_n585), .Z(new_n586));
  NAND3_X1  g385(.A1(new_n527), .A2(new_n535), .A3(new_n466), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT4), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT4), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n466), .A2(new_n589), .A3(new_n530), .A4(new_n534), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n590), .A2(KEYINPUT77), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT77), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n587), .A2(new_n593), .A3(KEYINPUT4), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G225gat), .A2(G233gat), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n466), .B1(new_n562), .B2(KEYINPUT3), .ZN(new_n597));
  AOI21_X1  g396(.A(KEYINPUT75), .B1(new_n597), .B2(new_n554), .ZN(new_n598));
  OAI21_X1  g397(.A(KEYINPUT3), .B1(new_n519), .B2(new_n526), .ZN(new_n599));
  INV_X1    g398(.A(new_n466), .ZN(new_n600));
  AND4_X1   g399(.A1(KEYINPUT75), .A2(new_n599), .A3(new_n600), .A4(new_n554), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n596), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT78), .B1(new_n595), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n596), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n599), .A2(new_n600), .A3(new_n554), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT75), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n597), .A2(KEYINPUT75), .A3(new_n554), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n604), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT78), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n609), .A2(new_n610), .A3(new_n592), .A4(new_n594), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n562), .B(new_n466), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT5), .B1(new_n612), .B2(new_n596), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n603), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n587), .A2(new_n589), .ZN(new_n616));
  INV_X1    g415(.A(new_n562), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n617), .A2(KEYINPUT4), .A3(new_n466), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT5), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n620), .A2(new_n609), .A3(KEYINPUT79), .A4(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT79), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n616), .A2(new_n621), .A3(new_n618), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n623), .B1(new_n602), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n586), .B1(new_n615), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT6), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n615), .A2(new_n586), .A3(new_n626), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n627), .A2(KEYINPUT6), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G226gat), .A2(G233gat), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n634), .B1(new_n481), .B2(KEYINPUT29), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(KEYINPUT72), .ZN(new_n636));
  INV_X1    g435(.A(new_n634), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n445), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n551), .B(new_n636), .C1(new_n640), .C2(KEYINPUT72), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n552), .ZN(new_n642));
  XNOR2_X1  g441(.A(G8gat), .B(G36gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(G64gat), .B(G92gat), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n643), .B(new_n644), .Z(new_n645));
  NAND3_X1  g444(.A1(new_n641), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n645), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT72), .B1(new_n635), .B2(new_n638), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT72), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n445), .A2(new_n555), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n649), .B1(new_n650), .B2(new_n634), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n648), .A2(new_n651), .A3(new_n552), .ZN(new_n652));
  INV_X1    g451(.A(new_n642), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n647), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n646), .A2(new_n654), .A3(KEYINPUT30), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n652), .A2(new_n653), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT30), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n656), .A2(new_n657), .A3(new_n645), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  XOR2_X1   g459(.A(KEYINPUT84), .B(KEYINPUT35), .Z(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n582), .A2(new_n633), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT80), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n629), .B(new_n630), .C1(new_n627), .C2(new_n665), .ZN(new_n666));
  AOI211_X1 g465(.A(KEYINPUT80), .B(new_n586), .C1(new_n615), .C2(new_n626), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n632), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(new_n659), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(KEYINPUT81), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT81), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n668), .A2(new_n671), .A3(new_n659), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n491), .A2(new_n499), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n498), .A2(new_n489), .A3(new_n490), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n581), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n670), .A2(new_n672), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n664), .B1(new_n677), .B2(KEYINPUT35), .ZN(new_n678));
  INV_X1    g477(.A(new_n581), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n679), .B1(new_n670), .B2(new_n672), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n598), .A2(new_n601), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n604), .B1(new_n681), .B2(new_n619), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n586), .B1(new_n682), .B2(KEYINPUT39), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT39), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n685), .B1(new_n612), .B2(new_n596), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT40), .B1(new_n684), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n687), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT40), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n689), .A2(new_n683), .A3(new_n690), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n688), .A2(new_n691), .A3(new_n627), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n581), .B1(new_n692), .B2(new_n660), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT37), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n645), .B1(new_n656), .B2(new_n694), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n552), .B(new_n636), .C1(new_n640), .C2(KEYINPUT72), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n694), .B1(new_n639), .B2(new_n551), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT38), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  AOI22_X1  g497(.A1(new_n695), .A2(new_n698), .B1(new_n656), .B2(new_n645), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n641), .A2(new_n642), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n647), .B1(new_n700), .B2(KEYINPUT37), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n656), .A2(new_n694), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT38), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n699), .A2(new_n703), .A3(new_n631), .A4(new_n632), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n693), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n673), .A2(new_n504), .A3(new_n674), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n502), .A2(KEYINPUT70), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT36), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n675), .A2(KEYINPUT36), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n705), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n680), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n401), .B1(new_n678), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT103), .ZN(new_n714));
  INV_X1    g513(.A(new_n668), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g516(.A(KEYINPUT16), .B(G8gat), .Z(new_n718));
  AND3_X1   g517(.A1(new_n714), .A2(new_n660), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n311), .B1(new_n714), .B2(new_n660), .ZN(new_n720));
  OAI21_X1  g519(.A(KEYINPUT42), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(KEYINPUT42), .B2(new_n719), .ZN(G1325gat));
  INV_X1    g521(.A(new_n505), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n714), .A2(new_n306), .A3(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT104), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n675), .A2(KEYINPUT36), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n726), .B(new_n727), .C1(new_n505), .C2(KEYINPUT36), .ZN(new_n728));
  OAI21_X1  g527(.A(KEYINPUT104), .B1(new_n708), .B2(new_n709), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n306), .B1(new_n714), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(KEYINPUT105), .B1(new_n725), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n714), .A2(new_n731), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n734), .B(new_n724), .C1(new_n735), .C2(new_n306), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n733), .A2(new_n736), .ZN(G1326gat));
  NAND2_X1  g536(.A1(new_n714), .A2(new_n581), .ZN(new_n738));
  XNOR2_X1  g537(.A(KEYINPUT43), .B(G22gat), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(G1327gat));
  NOR3_X1   g539(.A1(new_n396), .A2(new_n329), .A3(new_n363), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n273), .B(new_n741), .C1(new_n678), .C2(new_n712), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n742), .A2(G29gat), .A3(new_n668), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n743), .B(KEYINPUT45), .Z(new_n744));
  NAND2_X1  g543(.A1(new_n677), .A2(KEYINPUT35), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n663), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n668), .A2(new_n671), .A3(new_n659), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n671), .B1(new_n668), .B2(new_n659), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n581), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  AOI22_X1  g548(.A1(new_n728), .A2(new_n729), .B1(new_n704), .B2(new_n693), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n751), .B1(new_n749), .B2(new_n750), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n746), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n754), .A2(new_n755), .A3(new_n273), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n273), .B1(new_n678), .B2(new_n712), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT44), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n741), .ZN(new_n760));
  OAI21_X1  g559(.A(G29gat), .B1(new_n760), .B2(new_n668), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n744), .A2(new_n761), .ZN(G1328gat));
  OAI21_X1  g561(.A(G36gat), .B1(new_n760), .B2(new_n659), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n742), .A2(G36gat), .A3(new_n659), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT46), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(G1329gat));
  OAI21_X1  g565(.A(new_n207), .B1(new_n742), .B2(new_n505), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n731), .A2(G43gat), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n767), .B1(new_n760), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(KEYINPUT47), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT47), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n771), .B(new_n767), .C1(new_n760), .C2(new_n768), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(G1330gat));
  NAND3_X1  g572(.A1(new_n759), .A2(new_n581), .A3(new_n741), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n774), .A2(G50gat), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n679), .A2(G50gat), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT48), .B1(new_n742), .B2(new_n777), .ZN(new_n778));
  OR3_X1    g577(.A1(new_n742), .A2(KEYINPUT107), .A3(new_n777), .ZN(new_n779));
  OAI21_X1  g578(.A(KEYINPUT107), .B1(new_n742), .B2(new_n777), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(new_n774), .B2(G50gat), .ZN(new_n782));
  OAI22_X1  g581(.A1(new_n775), .A2(new_n778), .B1(new_n782), .B2(KEYINPUT48), .ZN(G1331gat));
  XNOR2_X1  g582(.A(new_n668), .B(KEYINPUT108), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n330), .A2(new_n397), .A3(new_n399), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n754), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g586(.A1(new_n754), .A2(new_n785), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n659), .ZN(new_n789));
  NOR2_X1   g588(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n790));
  AND2_X1   g589(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(new_n789), .B2(new_n790), .ZN(G1333gat));
  OAI21_X1  g592(.A(G71gat), .B1(new_n788), .B2(new_n730), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n723), .A2(new_n281), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n788), .B2(new_n795), .ZN(new_n796));
  XOR2_X1   g595(.A(new_n796), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g596(.A1(new_n788), .A2(new_n679), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(new_n282), .ZN(G1335gat));
  NOR2_X1   g598(.A1(new_n397), .A2(new_n329), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n363), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n759), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(G85gat), .B1(new_n803), .B2(new_n668), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n754), .A2(new_n273), .A3(new_n800), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT51), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n715), .A2(new_n229), .A3(new_n363), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n804), .B1(new_n809), .B2(new_n810), .ZN(G1336gat));
  AND3_X1   g610(.A1(new_n805), .A2(KEYINPUT109), .A3(KEYINPUT51), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT51), .B1(new_n805), .B2(KEYINPUT109), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n659), .A2(G92gat), .A3(new_n399), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n801), .B1(new_n756), .B2(new_n758), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n230), .B1(new_n817), .B2(new_n660), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT52), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(G92gat), .B1(new_n803), .B2(new_n659), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n814), .B1(new_n807), .B2(new_n808), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n819), .A2(new_n823), .ZN(G1337gat));
  OAI21_X1  g623(.A(G99gat), .B1(new_n803), .B2(new_n730), .ZN(new_n825));
  OR3_X1    g624(.A1(new_n505), .A2(G99gat), .A3(new_n399), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n825), .B1(new_n809), .B2(new_n826), .ZN(G1338gat));
  NOR3_X1   g626(.A1(new_n679), .A2(G106gat), .A3(new_n399), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n812), .A2(new_n813), .A3(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(G106gat), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n831), .B1(new_n817), .B2(new_n581), .ZN(new_n832));
  OAI21_X1  g631(.A(KEYINPUT53), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(G106gat), .B1(new_n803), .B2(new_n679), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n828), .B1(new_n807), .B2(new_n808), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n833), .A2(new_n837), .ZN(G1339gat));
  INV_X1    g637(.A(new_n329), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT110), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n353), .A2(new_n341), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n841), .B1(new_n842), .B2(new_n352), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n352), .A2(new_n353), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n340), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n358), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n847), .B1(new_n354), .B2(new_n841), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n846), .A2(new_n848), .A3(KEYINPUT55), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n360), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT55), .B1(new_n846), .B2(new_n848), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n840), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n846), .A2(new_n848), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT55), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n855), .A2(KEYINPUT110), .A3(new_n360), .A4(new_n849), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n852), .A2(new_n394), .A3(new_n395), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n382), .A2(new_n383), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n365), .B1(new_n378), .B2(new_n366), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n390), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n374), .A2(new_n384), .A3(new_n379), .A4(new_n392), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n363), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n273), .B1(new_n857), .B2(new_n864), .ZN(new_n865));
  AND4_X1   g664(.A1(new_n273), .A2(new_n863), .A3(new_n852), .A4(new_n856), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n839), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n274), .A2(new_n396), .A3(new_n329), .A4(new_n399), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n869), .A2(new_n659), .A3(new_n784), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n676), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(KEYINPUT111), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n447), .A3(new_n397), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n869), .A2(new_n582), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n715), .A3(new_n659), .ZN(new_n875));
  OAI21_X1  g674(.A(G113gat), .B1(new_n875), .B2(new_n396), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n873), .A2(new_n876), .ZN(G1340gat));
  NAND3_X1  g676(.A1(new_n872), .A2(new_n449), .A3(new_n363), .ZN(new_n878));
  OAI21_X1  g677(.A(G120gat), .B1(new_n875), .B2(new_n399), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(G1341gat));
  NOR3_X1   g679(.A1(new_n875), .A2(new_n452), .A3(new_n839), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n871), .A2(KEYINPUT112), .A3(new_n839), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n882), .A2(G127gat), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT112), .B1(new_n871), .B2(new_n839), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(G1342gat));
  NAND4_X1  g684(.A1(new_n870), .A2(new_n453), .A3(new_n676), .A4(new_n273), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n886), .A2(KEYINPUT56), .ZN(new_n887));
  XOR2_X1   g686(.A(new_n887), .B(KEYINPUT113), .Z(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(KEYINPUT56), .ZN(new_n889));
  XOR2_X1   g688(.A(new_n889), .B(KEYINPUT114), .Z(new_n890));
  OAI21_X1  g689(.A(G134gat), .B1(new_n875), .B2(new_n274), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n888), .A2(new_n890), .A3(new_n891), .ZN(G1343gat));
  NOR2_X1   g691(.A1(new_n731), .A2(new_n679), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n870), .A2(new_n893), .ZN(new_n894));
  AND3_X1   g693(.A1(new_n894), .A2(new_n514), .A3(new_n397), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n895), .A2(KEYINPUT117), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(KEYINPUT117), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT58), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n731), .A2(new_n668), .A3(new_n660), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT57), .B1(new_n869), .B2(new_n581), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n581), .A2(KEYINPUT57), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n850), .A2(new_n851), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n394), .A2(new_n902), .A3(new_n395), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n273), .B1(new_n903), .B2(new_n864), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n839), .B1(new_n866), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n901), .B1(new_n905), .B2(new_n868), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n899), .B1(new_n900), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(G141gat), .B1(new_n907), .B2(new_n396), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n896), .A2(new_n897), .A3(new_n898), .A4(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT115), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  OAI211_X1 g710(.A(KEYINPUT115), .B(new_n899), .C1(new_n900), .C2(new_n906), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(new_n397), .A3(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT116), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n913), .A2(new_n914), .A3(G141gat), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n914), .B1(new_n913), .B2(G141gat), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n915), .A2(new_n916), .A3(new_n895), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n909), .B1(new_n917), .B2(new_n898), .ZN(G1344gat));
  NAND4_X1  g717(.A1(new_n894), .A2(new_n520), .A3(new_n522), .A4(new_n363), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT118), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n919), .B(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n364), .A2(new_n396), .A3(new_n400), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT119), .B1(new_n273), .B2(new_n902), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n923), .A2(new_n862), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n273), .A2(KEYINPUT119), .A3(new_n902), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n904), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n922), .B1(new_n926), .B2(new_n329), .ZN(new_n927));
  AOI21_X1  g726(.A(KEYINPUT57), .B1(new_n927), .B2(new_n581), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n901), .B1(new_n867), .B2(new_n868), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n363), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n730), .A2(new_n715), .A3(new_n659), .ZN(new_n931));
  OAI21_X1  g730(.A(G148gat), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n932), .A2(KEYINPUT59), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n911), .A2(new_n363), .A3(new_n912), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n520), .A2(new_n522), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT59), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n921), .B(KEYINPUT120), .C1(new_n933), .C2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT120), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n919), .B(KEYINPUT118), .ZN(new_n942));
  AOI22_X1  g741(.A1(KEYINPUT59), .A2(new_n932), .B1(new_n934), .B2(new_n938), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n940), .A2(new_n944), .ZN(G1345gat));
  NAND3_X1  g744(.A1(new_n894), .A2(new_n508), .A3(new_n329), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n911), .A2(new_n912), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n947), .A2(new_n329), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n946), .B1(new_n948), .B2(new_n508), .ZN(G1346gat));
  AOI21_X1  g748(.A(G162gat), .B1(new_n894), .B2(new_n273), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n274), .A2(new_n509), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n950), .B1(new_n947), .B2(new_n951), .ZN(G1347gat));
  NOR2_X1   g751(.A1(new_n784), .A2(new_n659), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n953), .A2(KEYINPUT121), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(KEYINPUT121), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(new_n874), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n957), .A2(new_n416), .A3(new_n396), .ZN(new_n958));
  AOI211_X1 g757(.A(new_n715), .B(new_n659), .C1(new_n867), .C2(new_n868), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n959), .A2(new_n676), .ZN(new_n960));
  AOI21_X1  g759(.A(G169gat), .B1(new_n960), .B2(new_n397), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n958), .A2(new_n961), .ZN(G1348gat));
  OAI21_X1  g761(.A(G176gat), .B1(new_n957), .B2(new_n399), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n960), .A2(new_n417), .A3(new_n363), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1349gat));
  INV_X1    g764(.A(KEYINPUT122), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(KEYINPUT60), .ZN(new_n967));
  XOR2_X1   g766(.A(new_n967), .B(KEYINPUT123), .Z(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  OAI21_X1  g768(.A(G183gat), .B1(new_n957), .B2(new_n839), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n960), .A2(new_n427), .A3(new_n329), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g771(.A(new_n972), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n966), .A2(KEYINPUT60), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n969), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI211_X1 g774(.A(new_n972), .B(new_n968), .C1(new_n966), .C2(KEYINPUT60), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(G1350gat));
  NAND3_X1  g776(.A1(new_n960), .A2(new_n406), .A3(new_n273), .ZN(new_n978));
  OAI21_X1  g777(.A(G190gat), .B1(new_n957), .B2(new_n274), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(KEYINPUT124), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT61), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT124), .ZN(new_n982));
  OAI211_X1 g781(.A(new_n982), .B(G190gat), .C1(new_n957), .C2(new_n274), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n980), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n981), .B1(new_n980), .B2(new_n983), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n978), .B1(new_n984), .B2(new_n985), .ZN(G1351gat));
  AND2_X1   g785(.A1(new_n959), .A2(new_n893), .ZN(new_n987));
  AOI21_X1  g786(.A(G197gat), .B1(new_n987), .B2(new_n397), .ZN(new_n988));
  AND3_X1   g787(.A1(new_n954), .A2(new_n730), .A3(new_n955), .ZN(new_n989));
  XNOR2_X1  g788(.A(new_n989), .B(KEYINPUT125), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n928), .A2(new_n929), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AND2_X1   g791(.A1(new_n397), .A2(G197gat), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n988), .B1(new_n992), .B2(new_n993), .ZN(G1352gat));
  OAI21_X1  g793(.A(G204gat), .B1(new_n990), .B2(new_n930), .ZN(new_n995));
  INV_X1    g794(.A(G204gat), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n987), .A2(new_n996), .A3(new_n363), .ZN(new_n997));
  XOR2_X1   g796(.A(new_n997), .B(KEYINPUT62), .Z(new_n998));
  NAND2_X1  g797(.A1(new_n995), .A2(new_n998), .ZN(G1353gat));
  NAND2_X1  g798(.A1(new_n989), .A2(new_n329), .ZN(new_n1000));
  NOR2_X1   g799(.A1(new_n1000), .A2(new_n991), .ZN(new_n1001));
  OR3_X1    g800(.A1(new_n1001), .A2(KEYINPUT63), .A3(new_n543), .ZN(new_n1002));
  OAI21_X1  g801(.A(KEYINPUT63), .B1(new_n1001), .B2(new_n543), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n987), .A2(new_n543), .A3(new_n329), .ZN(new_n1004));
  XNOR2_X1  g803(.A(new_n1004), .B(KEYINPUT126), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(G1354gat));
  AOI21_X1  g805(.A(G218gat), .B1(new_n987), .B2(new_n273), .ZN(new_n1007));
  XOR2_X1   g806(.A(new_n1007), .B(KEYINPUT127), .Z(new_n1008));
  NOR2_X1   g807(.A1(new_n274), .A2(new_n544), .ZN(new_n1009));
  AOI21_X1  g808(.A(new_n1008), .B1(new_n992), .B2(new_n1009), .ZN(G1355gat));
endmodule


