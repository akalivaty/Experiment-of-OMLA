

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580;

  XOR2_X1 U319 ( .A(n366), .B(n365), .Z(n287) );
  NOR2_X1 U320 ( .A1(n571), .A2(n399), .ZN(n400) );
  XNOR2_X1 U321 ( .A(n367), .B(n287), .ZN(n368) );
  XNOR2_X1 U322 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U323 ( .A(KEYINPUT72), .B(n550), .ZN(n533) );
  XNOR2_X1 U324 ( .A(n449), .B(n448), .ZN(n524) );
  XNOR2_X1 U325 ( .A(n454), .B(G190GAT), .ZN(n455) );
  XNOR2_X1 U326 ( .A(n456), .B(n455), .ZN(G1351GAT) );
  XOR2_X1 U327 ( .A(G141GAT), .B(G22GAT), .Z(n289) );
  XNOR2_X1 U328 ( .A(G50GAT), .B(G113GAT), .ZN(n288) );
  XNOR2_X1 U329 ( .A(n289), .B(n288), .ZN(n293) );
  XOR2_X1 U330 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n291) );
  XNOR2_X1 U331 ( .A(G197GAT), .B(KEYINPUT66), .ZN(n290) );
  XNOR2_X1 U332 ( .A(n291), .B(n290), .ZN(n292) );
  XNOR2_X1 U333 ( .A(n293), .B(n292), .ZN(n301) );
  XNOR2_X1 U334 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n294) );
  XNOR2_X1 U335 ( .A(n294), .B(KEYINPUT7), .ZN(n364) );
  XOR2_X1 U336 ( .A(G15GAT), .B(G1GAT), .Z(n394) );
  XOR2_X1 U337 ( .A(n364), .B(n394), .Z(n296) );
  NAND2_X1 U338 ( .A1(G229GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U339 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U340 ( .A(G169GAT), .B(G8GAT), .Z(n425) );
  XOR2_X1 U341 ( .A(n297), .B(n425), .Z(n299) );
  XNOR2_X1 U342 ( .A(G36GAT), .B(G29GAT), .ZN(n298) );
  XNOR2_X1 U343 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U344 ( .A(n301), .B(n300), .ZN(n567) );
  XOR2_X1 U345 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n432) );
  XOR2_X1 U346 ( .A(G120GAT), .B(G57GAT), .Z(n340) );
  XOR2_X1 U347 ( .A(G127GAT), .B(KEYINPUT0), .Z(n303) );
  XNOR2_X1 U348 ( .A(G113GAT), .B(KEYINPUT77), .ZN(n302) );
  XNOR2_X1 U349 ( .A(n303), .B(n302), .ZN(n436) );
  XOR2_X1 U350 ( .A(n340), .B(n436), .Z(n305) );
  NAND2_X1 U351 ( .A1(G225GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U353 ( .A(n306), .B(KEYINPUT4), .Z(n309) );
  XNOR2_X1 U354 ( .A(G29GAT), .B(G134GAT), .ZN(n307) );
  XNOR2_X1 U355 ( .A(n307), .B(G85GAT), .ZN(n363) );
  XNOR2_X1 U356 ( .A(n363), .B(KEYINPUT88), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U358 ( .A(KEYINPUT86), .B(KEYINPUT1), .Z(n311) );
  XNOR2_X1 U359 ( .A(G1GAT), .B(G162GAT), .ZN(n310) );
  XNOR2_X1 U360 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U361 ( .A(n313), .B(n312), .Z(n321) );
  XOR2_X1 U362 ( .A(KEYINPUT3), .B(G155GAT), .Z(n315) );
  XNOR2_X1 U363 ( .A(KEYINPUT2), .B(G148GAT), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U365 ( .A(G141GAT), .B(n316), .Z(n334) );
  XOR2_X1 U366 ( .A(KEYINPUT6), .B(KEYINPUT87), .Z(n318) );
  XNOR2_X1 U367 ( .A(KEYINPUT89), .B(KEYINPUT5), .ZN(n317) );
  XNOR2_X1 U368 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U369 ( .A(n334), .B(n319), .ZN(n320) );
  XNOR2_X1 U370 ( .A(n321), .B(n320), .ZN(n466) );
  XOR2_X1 U371 ( .A(KEYINPUT90), .B(n466), .Z(n563) );
  XOR2_X1 U372 ( .A(KEYINPUT85), .B(KEYINPUT24), .Z(n323) );
  XNOR2_X1 U373 ( .A(G218GAT), .B(G106GAT), .ZN(n322) );
  XNOR2_X1 U374 ( .A(n323), .B(n322), .ZN(n327) );
  XOR2_X1 U375 ( .A(KEYINPUT22), .B(KEYINPUT84), .Z(n325) );
  XNOR2_X1 U376 ( .A(KEYINPUT80), .B(KEYINPUT23), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U378 ( .A(n327), .B(n326), .Z(n332) );
  XOR2_X1 U379 ( .A(G50GAT), .B(G162GAT), .Z(n358) );
  XOR2_X1 U380 ( .A(G22GAT), .B(G78GAT), .Z(n386) );
  XOR2_X1 U381 ( .A(KEYINPUT81), .B(n386), .Z(n329) );
  NAND2_X1 U382 ( .A1(G228GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U383 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U384 ( .A(n358), .B(n330), .ZN(n331) );
  XNOR2_X1 U385 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U386 ( .A(n334), .B(n333), .ZN(n339) );
  XOR2_X1 U387 ( .A(KEYINPUT82), .B(G204GAT), .Z(n336) );
  XNOR2_X1 U388 ( .A(G197GAT), .B(G211GAT), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n336), .B(n335), .ZN(n338) );
  XOR2_X1 U390 ( .A(KEYINPUT83), .B(KEYINPUT21), .Z(n337) );
  XOR2_X1 U391 ( .A(n338), .B(n337), .Z(n423) );
  XOR2_X1 U392 ( .A(n339), .B(n423), .Z(n468) );
  AND2_X1 U393 ( .A1(n563), .A2(n468), .ZN(n430) );
  XOR2_X1 U394 ( .A(G71GAT), .B(KEYINPUT13), .Z(n393) );
  XOR2_X1 U395 ( .A(G176GAT), .B(G64GAT), .Z(n421) );
  XOR2_X1 U396 ( .A(n393), .B(n421), .Z(n342) );
  XOR2_X1 U397 ( .A(G99GAT), .B(G106GAT), .Z(n357) );
  XNOR2_X1 U398 ( .A(n340), .B(n357), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n355) );
  XOR2_X1 U400 ( .A(KEYINPUT67), .B(KEYINPUT69), .Z(n344) );
  NAND2_X1 U401 ( .A1(G230GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U402 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U403 ( .A(n345), .B(KEYINPUT68), .Z(n353) );
  XOR2_X1 U404 ( .A(G92GAT), .B(G85GAT), .Z(n347) );
  XNOR2_X1 U405 ( .A(G148GAT), .B(G78GAT), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U407 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n349) );
  XNOR2_X1 U408 ( .A(G204GAT), .B(KEYINPUT31), .ZN(n348) );
  XNOR2_X1 U409 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U410 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U411 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U412 ( .A(n355), .B(n354), .Z(n571) );
  XOR2_X1 U413 ( .A(KEYINPUT45), .B(KEYINPUT109), .Z(n356) );
  XNOR2_X1 U414 ( .A(KEYINPUT65), .B(n356), .ZN(n398) );
  XNOR2_X1 U415 ( .A(KEYINPUT36), .B(KEYINPUT99), .ZN(n372) );
  XNOR2_X1 U416 ( .A(n358), .B(n357), .ZN(n371) );
  XOR2_X1 U417 ( .A(G92GAT), .B(G218GAT), .Z(n360) );
  XNOR2_X1 U418 ( .A(G36GAT), .B(G190GAT), .ZN(n359) );
  XNOR2_X1 U419 ( .A(n360), .B(n359), .ZN(n418) );
  XNOR2_X1 U420 ( .A(n418), .B(KEYINPUT11), .ZN(n362) );
  AND2_X1 U421 ( .A1(G232GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n362), .B(n361), .ZN(n369) );
  XNOR2_X1 U423 ( .A(n364), .B(n363), .ZN(n367) );
  XOR2_X1 U424 ( .A(KEYINPUT64), .B(KEYINPUT10), .Z(n366) );
  XNOR2_X1 U425 ( .A(KEYINPUT71), .B(KEYINPUT9), .ZN(n365) );
  XNOR2_X1 U426 ( .A(n371), .B(n370), .ZN(n550) );
  NAND2_X1 U427 ( .A1(n372), .A2(n533), .ZN(n376) );
  INV_X1 U428 ( .A(n372), .ZN(n374) );
  INV_X1 U429 ( .A(n533), .ZN(n373) );
  NAND2_X1 U430 ( .A1(n374), .A2(n373), .ZN(n375) );
  NAND2_X1 U431 ( .A1(n376), .A2(n375), .ZN(n576) );
  XOR2_X1 U432 ( .A(KEYINPUT15), .B(KEYINPUT73), .Z(n378) );
  NAND2_X1 U433 ( .A1(G231GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U435 ( .A(KEYINPUT14), .B(KEYINPUT76), .Z(n380) );
  XNOR2_X1 U436 ( .A(G8GAT), .B(KEYINPUT12), .ZN(n379) );
  XNOR2_X1 U437 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U438 ( .A(n382), .B(n381), .Z(n388) );
  XOR2_X1 U439 ( .A(KEYINPUT74), .B(KEYINPUT75), .Z(n384) );
  XNOR2_X1 U440 ( .A(G57GAT), .B(G64GAT), .ZN(n383) );
  XNOR2_X1 U441 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U443 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U444 ( .A(G211GAT), .B(G155GAT), .Z(n390) );
  XNOR2_X1 U445 ( .A(G183GAT), .B(G127GAT), .ZN(n389) );
  XNOR2_X1 U446 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U447 ( .A(n392), .B(n391), .Z(n396) );
  XNOR2_X1 U448 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U449 ( .A(n396), .B(n395), .Z(n559) );
  INV_X1 U450 ( .A(n559), .ZN(n574) );
  NAND2_X1 U451 ( .A1(n576), .A2(n574), .ZN(n397) );
  XOR2_X1 U452 ( .A(n398), .B(n397), .Z(n399) );
  XNOR2_X1 U453 ( .A(n400), .B(KEYINPUT110), .ZN(n401) );
  NAND2_X1 U454 ( .A1(n401), .A2(n567), .ZN(n410) );
  XOR2_X1 U455 ( .A(KEYINPUT47), .B(KEYINPUT108), .Z(n408) );
  XNOR2_X1 U456 ( .A(KEYINPUT46), .B(KEYINPUT107), .ZN(n402) );
  XNOR2_X1 U457 ( .A(n402), .B(KEYINPUT106), .ZN(n404) );
  XOR2_X1 U458 ( .A(n571), .B(KEYINPUT41), .Z(n498) );
  INV_X1 U459 ( .A(n498), .ZN(n552) );
  NOR2_X1 U460 ( .A1(n552), .A2(n567), .ZN(n403) );
  XOR2_X1 U461 ( .A(n404), .B(n403), .Z(n405) );
  NOR2_X1 U462 ( .A1(n574), .A2(n405), .ZN(n406) );
  NAND2_X1 U463 ( .A1(n406), .A2(n550), .ZN(n407) );
  XNOR2_X1 U464 ( .A(n408), .B(n407), .ZN(n409) );
  NAND2_X1 U465 ( .A1(n410), .A2(n409), .ZN(n412) );
  XNOR2_X1 U466 ( .A(KEYINPUT111), .B(KEYINPUT48), .ZN(n411) );
  XNOR2_X1 U467 ( .A(n412), .B(n411), .ZN(n539) );
  XOR2_X1 U468 ( .A(KEYINPUT93), .B(KEYINPUT91), .Z(n414) );
  NAND2_X1 U469 ( .A1(G226GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U470 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U471 ( .A(n415), .B(KEYINPUT92), .Z(n420) );
  XOR2_X1 U472 ( .A(G183GAT), .B(KEYINPUT17), .Z(n417) );
  XNOR2_X1 U473 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n416) );
  XNOR2_X1 U474 ( .A(n417), .B(n416), .ZN(n447) );
  XNOR2_X1 U475 ( .A(n447), .B(n418), .ZN(n419) );
  XNOR2_X1 U476 ( .A(n420), .B(n419), .ZN(n422) );
  XOR2_X1 U477 ( .A(n422), .B(n421), .Z(n427) );
  INV_X1 U478 ( .A(n423), .ZN(n424) );
  XOR2_X1 U479 ( .A(n425), .B(n424), .Z(n426) );
  XOR2_X1 U480 ( .A(n427), .B(n426), .Z(n514) );
  XOR2_X1 U481 ( .A(n514), .B(KEYINPUT118), .Z(n428) );
  NOR2_X1 U482 ( .A1(n539), .A2(n428), .ZN(n429) );
  XNOR2_X1 U483 ( .A(n429), .B(KEYINPUT54), .ZN(n564) );
  NAND2_X1 U484 ( .A1(n430), .A2(n564), .ZN(n431) );
  XNOR2_X1 U485 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U486 ( .A(n433), .B(KEYINPUT55), .ZN(n450) );
  XOR2_X1 U487 ( .A(G190GAT), .B(G43GAT), .Z(n435) );
  NAND2_X1 U488 ( .A1(G227GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U489 ( .A(n435), .B(n434), .ZN(n437) );
  XOR2_X1 U490 ( .A(n437), .B(n436), .Z(n445) );
  XOR2_X1 U491 ( .A(G176GAT), .B(KEYINPUT79), .Z(n439) );
  XNOR2_X1 U492 ( .A(G99GAT), .B(G134GAT), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n443) );
  XOR2_X1 U494 ( .A(KEYINPUT20), .B(G71GAT), .Z(n441) );
  XNOR2_X1 U495 ( .A(G169GAT), .B(G15GAT), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U498 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U499 ( .A(n446), .B(G120GAT), .Z(n449) );
  XNOR2_X1 U500 ( .A(n447), .B(KEYINPUT78), .ZN(n448) );
  NAND2_X1 U501 ( .A1(n450), .A2(n524), .ZN(n558) );
  NOR2_X1 U502 ( .A1(n567), .A2(n558), .ZN(n453) );
  XNOR2_X1 U503 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n451) );
  XNOR2_X1 U504 ( .A(n451), .B(G169GAT), .ZN(n452) );
  XNOR2_X1 U505 ( .A(n453), .B(n452), .ZN(G1348GAT) );
  NOR2_X1 U506 ( .A1(n533), .A2(n558), .ZN(n456) );
  XNOR2_X1 U507 ( .A(KEYINPUT125), .B(KEYINPUT58), .ZN(n454) );
  INV_X1 U508 ( .A(n563), .ZN(n512) );
  NOR2_X1 U509 ( .A1(n567), .A2(n571), .ZN(n457) );
  XOR2_X1 U510 ( .A(KEYINPUT70), .B(n457), .Z(n488) );
  NAND2_X1 U511 ( .A1(n514), .A2(n524), .ZN(n458) );
  NAND2_X1 U512 ( .A1(n458), .A2(n468), .ZN(n459) );
  XNOR2_X1 U513 ( .A(n459), .B(KEYINPUT25), .ZN(n460) );
  XOR2_X1 U514 ( .A(KEYINPUT95), .B(n460), .Z(n464) );
  NOR2_X1 U515 ( .A1(n468), .A2(n524), .ZN(n461) );
  XNOR2_X1 U516 ( .A(n461), .B(KEYINPUT26), .ZN(n565) );
  INV_X1 U517 ( .A(n565), .ZN(n540) );
  XOR2_X1 U518 ( .A(n514), .B(KEYINPUT94), .Z(n462) );
  XNOR2_X1 U519 ( .A(n462), .B(KEYINPUT27), .ZN(n467) );
  NOR2_X1 U520 ( .A1(n540), .A2(n467), .ZN(n463) );
  NOR2_X1 U521 ( .A1(n464), .A2(n463), .ZN(n465) );
  NOR2_X1 U522 ( .A1(n466), .A2(n465), .ZN(n471) );
  NOR2_X1 U523 ( .A1(n563), .A2(n467), .ZN(n542) );
  XOR2_X1 U524 ( .A(KEYINPUT28), .B(n468), .Z(n519) );
  INV_X1 U525 ( .A(n519), .ZN(n469) );
  NAND2_X1 U526 ( .A1(n542), .A2(n469), .ZN(n522) );
  NOR2_X1 U527 ( .A1(n524), .A2(n522), .ZN(n470) );
  NOR2_X1 U528 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U529 ( .A(KEYINPUT96), .B(n472), .ZN(n484) );
  NAND2_X1 U530 ( .A1(n574), .A2(n533), .ZN(n473) );
  XNOR2_X1 U531 ( .A(KEYINPUT16), .B(n473), .ZN(n474) );
  OR2_X1 U532 ( .A1(n484), .A2(n474), .ZN(n499) );
  NOR2_X1 U533 ( .A1(n488), .A2(n499), .ZN(n481) );
  NAND2_X1 U534 ( .A1(n512), .A2(n481), .ZN(n477) );
  XOR2_X1 U535 ( .A(G1GAT), .B(KEYINPUT34), .Z(n475) );
  XNOR2_X1 U536 ( .A(KEYINPUT97), .B(n475), .ZN(n476) );
  XNOR2_X1 U537 ( .A(n477), .B(n476), .ZN(G1324GAT) );
  NAND2_X1 U538 ( .A1(n514), .A2(n481), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n478), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U540 ( .A(G15GAT), .B(KEYINPUT35), .Z(n480) );
  NAND2_X1 U541 ( .A1(n481), .A2(n524), .ZN(n479) );
  XNOR2_X1 U542 ( .A(n480), .B(n479), .ZN(G1326GAT) );
  NAND2_X1 U543 ( .A1(n519), .A2(n481), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n482), .B(KEYINPUT98), .ZN(n483) );
  XNOR2_X1 U545 ( .A(G22GAT), .B(n483), .ZN(G1327GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT39), .B(KEYINPUT101), .Z(n491) );
  XOR2_X1 U547 ( .A(KEYINPUT37), .B(KEYINPUT100), .Z(n487) );
  NOR2_X1 U548 ( .A1(n574), .A2(n484), .ZN(n485) );
  NAND2_X1 U549 ( .A1(n485), .A2(n576), .ZN(n486) );
  XNOR2_X1 U550 ( .A(n487), .B(n486), .ZN(n511) );
  NOR2_X1 U551 ( .A1(n488), .A2(n511), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n489), .B(KEYINPUT38), .ZN(n496) );
  NAND2_X1 U553 ( .A1(n496), .A2(n512), .ZN(n490) );
  XNOR2_X1 U554 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U555 ( .A(G29GAT), .B(n492), .Z(G1328GAT) );
  NAND2_X1 U556 ( .A1(n496), .A2(n514), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n493), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U558 ( .A1(n496), .A2(n524), .ZN(n494) );
  XNOR2_X1 U559 ( .A(n494), .B(KEYINPUT40), .ZN(n495) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  NAND2_X1 U561 ( .A1(n496), .A2(n519), .ZN(n497) );
  XNOR2_X1 U562 ( .A(n497), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT102), .B(KEYINPUT42), .Z(n501) );
  NAND2_X1 U564 ( .A1(n567), .A2(n498), .ZN(n510) );
  NOR2_X1 U565 ( .A1(n510), .A2(n499), .ZN(n507) );
  NAND2_X1 U566 ( .A1(n507), .A2(n512), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U568 ( .A(G57GAT), .B(n502), .Z(G1332GAT) );
  XOR2_X1 U569 ( .A(G64GAT), .B(KEYINPUT103), .Z(n504) );
  NAND2_X1 U570 ( .A1(n507), .A2(n514), .ZN(n503) );
  XNOR2_X1 U571 ( .A(n504), .B(n503), .ZN(G1333GAT) );
  NAND2_X1 U572 ( .A1(n507), .A2(n524), .ZN(n505) );
  XNOR2_X1 U573 ( .A(n505), .B(KEYINPUT104), .ZN(n506) );
  XNOR2_X1 U574 ( .A(G71GAT), .B(n506), .ZN(G1334GAT) );
  XOR2_X1 U575 ( .A(G78GAT), .B(KEYINPUT43), .Z(n509) );
  NAND2_X1 U576 ( .A1(n507), .A2(n519), .ZN(n508) );
  XNOR2_X1 U577 ( .A(n509), .B(n508), .ZN(G1335GAT) );
  NOR2_X1 U578 ( .A1(n511), .A2(n510), .ZN(n518) );
  NAND2_X1 U579 ( .A1(n518), .A2(n512), .ZN(n513) );
  XNOR2_X1 U580 ( .A(G85GAT), .B(n513), .ZN(G1336GAT) );
  NAND2_X1 U581 ( .A1(n514), .A2(n518), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n515), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U583 ( .A(G99GAT), .B(KEYINPUT105), .Z(n517) );
  NAND2_X1 U584 ( .A1(n518), .A2(n524), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n517), .B(n516), .ZN(G1338GAT) );
  NAND2_X1 U586 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n520), .B(KEYINPUT44), .ZN(n521) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(n521), .ZN(G1339GAT) );
  NOR2_X1 U589 ( .A1(n539), .A2(n522), .ZN(n523) );
  NAND2_X1 U590 ( .A1(n524), .A2(n523), .ZN(n534) );
  NOR2_X1 U591 ( .A1(n567), .A2(n534), .ZN(n525) );
  XOR2_X1 U592 ( .A(G113GAT), .B(n525), .Z(G1340GAT) );
  NOR2_X1 U593 ( .A1(n534), .A2(n552), .ZN(n529) );
  XOR2_X1 U594 ( .A(KEYINPUT112), .B(KEYINPUT49), .Z(n527) );
  XNOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT113), .ZN(n526) );
  XNOR2_X1 U596 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U597 ( .A(n529), .B(n528), .ZN(G1341GAT) );
  NOR2_X1 U598 ( .A1(n559), .A2(n534), .ZN(n531) );
  XNOR2_X1 U599 ( .A(KEYINPUT50), .B(KEYINPUT114), .ZN(n530) );
  XNOR2_X1 U600 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U601 ( .A(G127GAT), .B(n532), .Z(G1342GAT) );
  NOR2_X1 U602 ( .A1(n534), .A2(n533), .ZN(n538) );
  XOR2_X1 U603 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n536) );
  XNOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT116), .ZN(n535) );
  XNOR2_X1 U605 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U606 ( .A(n538), .B(n537), .ZN(G1343GAT) );
  NOR2_X1 U607 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n549) );
  NOR2_X1 U609 ( .A1(n567), .A2(n549), .ZN(n543) );
  XOR2_X1 U610 ( .A(G141GAT), .B(n543), .Z(G1344GAT) );
  NOR2_X1 U611 ( .A1(n549), .A2(n552), .ZN(n547) );
  XOR2_X1 U612 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n545) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n544) );
  XNOR2_X1 U614 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(G1345GAT) );
  NOR2_X1 U616 ( .A1(n559), .A2(n549), .ZN(n548) );
  XOR2_X1 U617 ( .A(G155GAT), .B(n548), .Z(G1346GAT) );
  NOR2_X1 U618 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U619 ( .A(G162GAT), .B(n551), .Z(G1347GAT) );
  NOR2_X1 U620 ( .A1(n552), .A2(n558), .ZN(n557) );
  XOR2_X1 U621 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n554) );
  XNOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n553) );
  XNOR2_X1 U623 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U624 ( .A(KEYINPUT56), .B(n555), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(G1349GAT) );
  NOR2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U627 ( .A(G183GAT), .B(n560), .Z(G1350GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n562) );
  XNOR2_X1 U629 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(n569) );
  AND2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n566) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n570) );
  NOR2_X1 U633 ( .A1(n567), .A2(n570), .ZN(n568) );
  XOR2_X1 U634 ( .A(n569), .B(n568), .Z(G1352GAT) );
  XOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .Z(n573) );
  INV_X1 U636 ( .A(n570), .ZN(n577) );
  NAND2_X1 U637 ( .A1(n577), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  NAND2_X1 U639 ( .A1(n577), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n579) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(n580), .ZN(G1355GAT) );
endmodule

