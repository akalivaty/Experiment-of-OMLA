//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n630,
    new_n633, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT64), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n464), .B(KEYINPUT66), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  AOI22_X1  g046(.A1(G101), .A2(new_n465), .B1(new_n471), .B2(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n473), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(new_n470), .A2(new_n463), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n471), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NAND2_X1  g060(.A1(new_n471), .A2(G138), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT4), .ZN(new_n487));
  OR2_X1    g062(.A1(new_n463), .A2(G114), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AOI22_X1  g065(.A1(new_n479), .A2(G126), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G164));
  INV_X1    g068(.A(G651), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT67), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT67), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G651), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT6), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n494), .B1(KEYINPUT68), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT6), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n498), .A2(KEYINPUT6), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(KEYINPUT5), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n504), .A2(KEYINPUT69), .A3(G543), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n503), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n496), .A2(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n494), .A2(KEYINPUT67), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT6), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n499), .A2(KEYINPUT68), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n502), .A2(new_n516), .A3(G651), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n515), .A2(G543), .A3(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G50), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n511), .A2(new_n512), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n521), .A2(new_n498), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n520), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND3_X1  g099(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n525));
  XOR2_X1   g100(.A(KEYINPUT70), .B(G51), .Z(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n518), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT71), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n529), .B(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n511), .ZN(new_n532));
  XOR2_X1   g107(.A(KEYINPUT73), .B(G89), .Z(new_n533));
  AOI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n528), .A2(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n511), .A2(new_n537), .B1(new_n518), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT74), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(new_n498), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  INV_X1    g120(.A(G43), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n511), .A2(new_n545), .B1(new_n518), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT75), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n498), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(KEYINPUT75), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n547), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT76), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT77), .Z(G188));
  INV_X1    g136(.A(G91), .ZN(new_n562));
  XNOR2_X1  g137(.A(KEYINPUT67), .B(G651), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n499), .A2(KEYINPUT68), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n501), .B2(KEYINPUT6), .ZN(new_n565));
  OAI22_X1  g140(.A1(new_n563), .A2(new_n499), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n567));
  AND3_X1   g142(.A1(new_n504), .A2(KEYINPUT69), .A3(G543), .ZN(new_n568));
  AOI21_X1  g143(.A(KEYINPUT69), .B1(new_n504), .B2(G543), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT78), .B1(new_n566), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT78), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n510), .A2(new_n515), .A3(new_n572), .A4(new_n517), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n562), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n510), .A2(G65), .ZN(new_n575));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n494), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n515), .A2(G53), .A3(G543), .A4(new_n517), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT9), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(G299));
  NAND2_X1  g156(.A1(new_n571), .A2(new_n573), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n582), .A2(G87), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n584));
  INV_X1    g159(.A(G49), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n518), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G288));
  INV_X1    g163(.A(new_n518), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G48), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n510), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n498), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n582), .A2(G86), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n592), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n593), .A2(KEYINPUT79), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(G72), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G60), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n570), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT80), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n498), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(new_n602), .B2(new_n601), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n532), .A2(G85), .B1(new_n589), .B2(G47), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  INV_X1    g182(.A(G54), .ZN(new_n608));
  NOR3_X1   g183(.A1(new_n566), .A2(new_n608), .A3(new_n507), .ZN(new_n609));
  OAI211_X1 g184(.A(G66), .B(new_n567), .C1(new_n568), .C2(new_n569), .ZN(new_n610));
  NAND2_X1  g185(.A1(G79), .A2(G543), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n494), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(KEYINPUT81), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n503), .A2(G54), .A3(G543), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT81), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n510), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n614), .B(new_n615), .C1(new_n494), .C2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g193(.A(KEYINPUT10), .B1(new_n582), .B2(G92), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT10), .ZN(new_n620));
  INV_X1    g195(.A(G92), .ZN(new_n621));
  AOI211_X1 g196(.A(new_n620), .B(new_n621), .C1(new_n571), .C2(new_n573), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n618), .B1(new_n619), .B2(new_n622), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n623), .A2(KEYINPUT82), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(KEYINPUT82), .ZN(new_n625));
  AND2_X1   g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n607), .B1(new_n626), .B2(G868), .ZN(G284));
  OAI21_X1  g202(.A(new_n607), .B1(new_n626), .B2(G868), .ZN(G321));
  INV_X1    g203(.A(G868), .ZN(new_n629));
  NAND2_X1  g204(.A1(G299), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(G168), .B2(new_n629), .ZN(G297));
  OAI21_X1  g206(.A(new_n630), .B1(G168), .B2(new_n629), .ZN(G280));
  INV_X1    g207(.A(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n626), .B1(new_n633), .B2(G860), .ZN(G148));
  NAND2_X1  g209(.A1(new_n626), .A2(new_n633), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(G868), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g213(.A(new_n470), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n465), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(KEYINPUT83), .B(KEYINPUT12), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT13), .B(G2100), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n479), .A2(G123), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT84), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n479), .A2(KEYINPUT84), .A3(G123), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n471), .A2(G135), .ZN(new_n649));
  OR3_X1    g224(.A1(new_n463), .A2(KEYINPUT85), .A3(G111), .ZN(new_n650));
  OAI21_X1  g225(.A(KEYINPUT85), .B1(new_n463), .B2(G111), .ZN(new_n651));
  OR2_X1    g226(.A1(G99), .A2(G2105), .ZN(new_n652));
  NAND4_X1  g227(.A1(new_n650), .A2(G2104), .A3(new_n651), .A4(new_n652), .ZN(new_n653));
  NAND4_X1  g228(.A1(new_n647), .A2(new_n648), .A3(new_n649), .A4(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT86), .B(G2096), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n644), .A2(new_n657), .A3(new_n658), .ZN(G156));
  XOR2_X1   g234(.A(KEYINPUT15), .B(G2435), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2438), .ZN(new_n661));
  XOR2_X1   g236(.A(G2427), .B(G2430), .Z(new_n662));
  OAI21_X1  g237(.A(KEYINPUT14), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT87), .Z(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2451), .B(G2454), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT16), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2443), .B(G2446), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1341), .B(G1348), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n673), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n674), .A2(G14), .A3(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G401));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G2067), .B(G2678), .Z(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G2072), .B(G2078), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT18), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n679), .A2(new_n680), .ZN(new_n685));
  AND3_X1   g260(.A1(new_n685), .A2(KEYINPUT17), .A3(new_n682), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n682), .B1(new_n685), .B2(KEYINPUT17), .ZN(new_n687));
  NOR3_X1   g262(.A1(new_n686), .A2(new_n687), .A3(new_n681), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G2096), .B(G2100), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(G227));
  XNOR2_X1  g266(.A(G1971), .B(G1976), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT19), .ZN(new_n693));
  XOR2_X1   g268(.A(G1956), .B(G2474), .Z(new_n694));
  XOR2_X1   g269(.A(G1961), .B(G1966), .Z(new_n695));
  OR2_X1    g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n693), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n693), .A2(new_n697), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  OAI221_X1 g277(.A(new_n698), .B1(new_n693), .B2(new_n696), .C1(new_n700), .C2(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n700), .B2(new_n702), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(G1991), .ZN(new_n705));
  INV_X1    g280(.A(G1996), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1981), .B(G1986), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n708), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n707), .B(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n710), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n711), .A2(new_n715), .ZN(G229));
  NAND2_X1  g291(.A1(new_n465), .A2(G105), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT97), .Z(new_n718));
  NAND2_X1  g293(.A1(new_n479), .A2(G129), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n471), .A2(G141), .ZN(new_n720));
  NAND3_X1  g295(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT26), .Z(new_n722));
  NAND3_X1  g297(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n718), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G29), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G29), .B2(G32), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT27), .B(G1996), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(G164), .A2(G29), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G27), .B2(G29), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT98), .B(G2078), .Z(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  AND2_X1   g307(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n726), .A2(new_n727), .ZN(new_n734));
  NOR3_X1   g309(.A1(new_n728), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT31), .B(G11), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT30), .B(G28), .Z(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n737), .B2(G29), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n655), .B2(G29), .ZN(new_n739));
  INV_X1    g314(.A(G29), .ZN(new_n740));
  AND2_X1   g315(.A1(KEYINPUT24), .A2(G34), .ZN(new_n741));
  NOR2_X1   g316(.A1(KEYINPUT24), .A2(G34), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT95), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G160), .B2(G29), .ZN(new_n746));
  OAI221_X1 g321(.A(new_n739), .B1(G2084), .B2(new_n746), .C1(new_n730), .C2(new_n732), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n740), .A2(G35), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G162), .B2(new_n740), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT29), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(G2090), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n740), .A2(G26), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n479), .A2(G128), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n471), .A2(G140), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n463), .A2(G116), .ZN(new_n756));
  OAI21_X1  g331(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n754), .B(new_n755), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n753), .B1(new_n758), .B2(G29), .ZN(new_n759));
  MUX2_X1   g334(.A(new_n753), .B(new_n759), .S(KEYINPUT28), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G2067), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n746), .A2(G2084), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT96), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G2090), .B2(new_n750), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n735), .A2(new_n752), .A3(new_n761), .A4(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G16), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G21), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G168), .B2(new_n766), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1966), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n740), .A2(G33), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT25), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n471), .A2(G139), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT93), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n639), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n463), .B2(new_n777), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT94), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n771), .B1(new_n779), .B2(new_n740), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G2072), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n766), .A2(G5), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G171), .B2(new_n766), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1961), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT23), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n766), .A2(G20), .ZN(new_n787));
  AOI211_X1 g362(.A(new_n786), .B(new_n787), .C1(G299), .C2(G16), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n786), .B2(new_n787), .ZN(new_n789));
  INV_X1    g364(.A(G1956), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n766), .A2(G19), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n553), .B2(new_n766), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT92), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT91), .B(G1341), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n770), .A2(new_n785), .A3(new_n791), .A4(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(G4), .A2(G16), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT90), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n624), .A2(new_n625), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n766), .ZN(new_n801));
  INV_X1    g376(.A(G1348), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n797), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT89), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT36), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(G16), .A2(G23), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n587), .B2(G16), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT33), .B(G1976), .Z(new_n810));
  AND2_X1   g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n766), .A2(G22), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G166), .B2(new_n766), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n813), .A2(G1971), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n809), .A2(new_n810), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n813), .A2(G1971), .ZN(new_n816));
  NOR4_X1   g391(.A1(new_n811), .A2(new_n814), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT32), .B(G1981), .Z(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n766), .B1(new_n596), .B2(new_n597), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n766), .A2(G6), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OR3_X1    g397(.A1(new_n820), .A2(new_n821), .A3(new_n819), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n817), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT34), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n817), .A2(new_n822), .A3(KEYINPUT34), .A4(new_n823), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(G290), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n829), .A2(new_n766), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(new_n766), .B2(G24), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(G1986), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n479), .A2(G119), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n471), .A2(G131), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n463), .A2(G107), .ZN(new_n835));
  OAI21_X1  g410(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n833), .B(new_n834), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  MUX2_X1   g412(.A(G25), .B(new_n837), .S(G29), .Z(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT35), .B(G1991), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n838), .B(new_n839), .Z(new_n840));
  AND2_X1   g415(.A1(new_n832), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n828), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n805), .A2(new_n806), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n807), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AOI211_X1 g419(.A(new_n805), .B(new_n806), .C1(new_n828), .C2(new_n841), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n804), .B1(new_n844), .B2(new_n845), .ZN(G150));
  NAND2_X1  g421(.A1(G150), .A2(KEYINPUT99), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT99), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n848), .B(new_n804), .C1(new_n844), .C2(new_n845), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(G311));
  AOI22_X1  g425(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n851), .A2(new_n498), .ZN(new_n852));
  XOR2_X1   g427(.A(KEYINPUT100), .B(G93), .Z(new_n853));
  NAND4_X1  g428(.A1(new_n510), .A2(new_n515), .A3(new_n517), .A4(new_n853), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n515), .A2(G55), .A3(G543), .A4(new_n517), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n854), .A2(KEYINPUT101), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(KEYINPUT101), .B1(new_n854), .B2(new_n855), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n852), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(G860), .ZN(new_n859));
  XOR2_X1   g434(.A(KEYINPUT104), .B(KEYINPUT37), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n858), .A2(KEYINPUT102), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n551), .A2(new_n552), .ZN(new_n863));
  INV_X1    g438(.A(new_n547), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT102), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n866), .B(new_n852), .C1(new_n856), .C2(new_n857), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n862), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n858), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n869), .A2(new_n866), .A3(new_n553), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT38), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n800), .A2(new_n633), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(G860), .B1(new_n874), .B2(KEYINPUT39), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(KEYINPUT39), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n875), .B1(new_n876), .B2(KEYINPUT103), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n876), .A2(KEYINPUT103), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n861), .B1(new_n877), .B2(new_n878), .ZN(G145));
  AND2_X1   g454(.A1(new_n779), .A2(KEYINPUT105), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n779), .A2(KEYINPUT105), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n492), .B(new_n758), .ZN(new_n882));
  INV_X1    g457(.A(new_n724), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n882), .B(new_n883), .ZN(new_n884));
  OR3_X1    g459(.A1(new_n880), .A2(new_n881), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n880), .A2(new_n884), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n471), .A2(G142), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n463), .A2(G118), .ZN(new_n889));
  OAI21_X1  g464(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n891), .B1(G130), .B2(new_n479), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n892), .B(KEYINPUT106), .Z(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(new_n837), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n642), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n887), .A2(new_n895), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n894), .B(new_n642), .Z(new_n897));
  NAND3_X1  g472(.A1(new_n897), .A2(new_n885), .A3(new_n886), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n477), .B(new_n484), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(new_n654), .ZN(new_n901));
  AOI21_X1  g476(.A(G37), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n898), .A2(KEYINPUT107), .ZN(new_n903));
  INV_X1    g478(.A(new_n901), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n896), .B(new_n904), .C1(new_n898), .C2(KEYINPUT107), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n902), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g482(.A1(G288), .A2(new_n829), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n587), .A2(G290), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(KEYINPUT111), .ZN(new_n911));
  NAND2_X1  g486(.A1(G305), .A2(G166), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n596), .A2(G303), .A3(new_n597), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT111), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n908), .A2(new_n916), .A3(new_n909), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n911), .A2(new_n914), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  XOR2_X1   g494(.A(new_n919), .B(KEYINPUT42), .Z(new_n920));
  XOR2_X1   g495(.A(new_n635), .B(new_n871), .Z(new_n921));
  AOI21_X1  g496(.A(new_n572), .B1(new_n503), .B2(new_n510), .ZN(new_n922));
  AND4_X1   g497(.A1(new_n572), .A2(new_n510), .A3(new_n515), .A4(new_n517), .ZN(new_n923));
  OAI21_X1  g498(.A(G92), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n620), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n582), .A2(KEYINPUT10), .A3(G92), .ZN(new_n926));
  AOI22_X1  g501(.A1(new_n925), .A2(new_n926), .B1(new_n617), .B2(new_n613), .ZN(new_n927));
  AOI21_X1  g502(.A(KEYINPUT108), .B1(new_n927), .B2(G299), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT9), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n579), .B(new_n930), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n931), .A2(new_n574), .A3(new_n577), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n623), .A2(new_n929), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT109), .B1(new_n928), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n929), .B1(new_n623), .B2(new_n932), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n925), .A2(new_n926), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n936), .A2(G299), .A3(KEYINPUT108), .A4(new_n618), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT109), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n935), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n623), .A2(new_n932), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n934), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  OR2_X1    g517(.A1(new_n921), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT112), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n934), .A2(KEYINPUT41), .A3(new_n939), .A4(new_n940), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT110), .ZN(new_n946));
  AOI22_X1  g521(.A1(new_n935), .A2(new_n937), .B1(new_n932), .B2(new_n623), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n946), .B1(new_n947), .B2(KEYINPUT41), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n940), .B1(new_n928), .B2(new_n933), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT41), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(KEYINPUT110), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n945), .A2(new_n948), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n921), .A2(new_n952), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n920), .A2(new_n943), .A3(new_n944), .A4(new_n953), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n943), .A2(new_n953), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n954), .B1(new_n955), .B2(new_n920), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n944), .B1(new_n955), .B2(new_n920), .ZN(new_n957));
  OAI21_X1  g532(.A(G868), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n858), .A2(new_n629), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(G295));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n959), .ZN(G331));
  AND3_X1   g536(.A1(new_n868), .A2(new_n870), .A3(G301), .ZN(new_n962));
  AOI21_X1  g537(.A(G301), .B1(new_n868), .B2(new_n870), .ZN(new_n963));
  OAI21_X1  g538(.A(G286), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n871), .A2(G171), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n868), .A2(new_n870), .A3(G301), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n965), .A2(G168), .A3(new_n966), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n952), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n919), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n964), .A2(new_n967), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n941), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n969), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT113), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n969), .A2(new_n972), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n919), .ZN(new_n977));
  INV_X1    g552(.A(G37), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n969), .A2(new_n970), .A3(KEYINPUT113), .A4(new_n972), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n975), .A2(new_n977), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT43), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(G37), .B1(new_n973), .B2(new_n974), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT114), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(new_n949), .B2(new_n950), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n947), .A2(KEYINPUT114), .A3(KEYINPUT41), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n968), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n987), .B(new_n972), .C1(new_n942), .C2(KEYINPUT41), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n919), .ZN(new_n989));
  AND4_X1   g564(.A1(KEYINPUT43), .A2(new_n983), .A3(new_n989), .A4(new_n979), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT44), .B1(new_n982), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n983), .A2(new_n989), .A3(new_n981), .A4(new_n979), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n991), .A2(new_n996), .ZN(G397));
  INV_X1    g572(.A(G1384), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n492), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(KEYINPUT115), .B(KEYINPUT45), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n472), .A2(G40), .A3(new_n476), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G2067), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n758), .B(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n1007), .B(KEYINPUT116), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n883), .A2(G1996), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n724), .A2(new_n706), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n837), .B(new_n839), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(G290), .B(G1986), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1005), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(G1384), .B1(new_n487), .B2(new_n491), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n1003), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(G8), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1018), .B1(G1976), .B2(new_n587), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1019), .B(new_n1020), .C1(G1976), .C2(new_n587), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(new_n1020), .B2(new_n1019), .ZN(new_n1022));
  OR2_X1    g597(.A1(G305), .A2(G1981), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n591), .A2(new_n498), .ZN(new_n1024));
  INV_X1    g599(.A(G86), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n590), .B1(new_n1025), .B2(new_n511), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1024), .B1(new_n1026), .B2(KEYINPUT118), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1027), .B1(KEYINPUT118), .B2(new_n1026), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(G1981), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1023), .A2(KEYINPUT49), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT119), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1023), .A2(KEYINPUT119), .A3(KEYINPUT49), .A4(new_n1029), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT49), .B1(new_n1023), .B2(new_n1029), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1035), .A2(new_n1018), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1022), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G8), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1016), .A2(KEYINPUT45), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1002), .A2(new_n1003), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G1971), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1004), .B1(new_n999), .B2(KEYINPUT50), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT50), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1016), .A2(new_n1044), .ZN(new_n1045));
  XOR2_X1   g620(.A(KEYINPUT117), .B(G2090), .Z(new_n1046));
  NAND3_X1  g621(.A1(new_n1043), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1038), .B1(new_n1042), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(G303), .A2(G8), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n1049), .B(KEYINPUT55), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1048), .B(new_n1050), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n1037), .A2(KEYINPUT126), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT126), .B1(new_n1037), .B2(new_n1051), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT123), .ZN(new_n1055));
  XNOR2_X1  g630(.A(KEYINPUT56), .B(G2072), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1002), .A2(new_n1003), .A3(new_n1039), .A4(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(G1956), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1055), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n999), .A2(KEYINPUT50), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1061), .A2(new_n1003), .A3(new_n1045), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n790), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1063), .A2(KEYINPUT123), .A3(new_n1057), .ZN(new_n1064));
  XNOR2_X1  g639(.A(G299), .B(KEYINPUT57), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1060), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1065), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(new_n1063), .A3(new_n1057), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1066), .A2(KEYINPUT61), .A3(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1002), .A2(new_n706), .A3(new_n1003), .A4(new_n1039), .ZN(new_n1070));
  XOR2_X1   g645(.A(KEYINPUT58), .B(G1341), .Z(new_n1071));
  NAND2_X1  g646(.A1(new_n1017), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n865), .A2(KEYINPUT124), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT59), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1073), .A2(new_n1077), .A3(new_n1074), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1017), .A2(G2067), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1079), .B1(new_n1062), .B2(new_n802), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n800), .A2(KEYINPUT60), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1076), .A2(new_n1078), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1080), .A2(new_n800), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1080), .A2(new_n800), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT60), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT61), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1068), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1067), .B1(new_n1063), .B2(new_n1057), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1086), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1069), .A2(new_n1082), .A3(new_n1085), .A4(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1084), .A2(KEYINPUT122), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1091), .A2(new_n1087), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1084), .A2(KEYINPUT122), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1090), .A2(new_n1066), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1004), .B1(new_n1016), .B2(new_n1000), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(KEYINPUT45), .B2(new_n1016), .ZN(new_n1098));
  INV_X1    g673(.A(G2078), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT53), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1002), .A2(new_n1099), .A3(new_n1003), .A4(new_n1039), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(G1961), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1062), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1101), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(G171), .ZN(new_n1108));
  OR2_X1    g683(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1109), .B1(new_n1110), .B2(KEYINPUT125), .ZN(new_n1111));
  OR3_X1    g686(.A1(new_n1102), .A2(KEYINPUT125), .A3(new_n1103), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1111), .A2(new_n1112), .A3(new_n1106), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1104), .A2(G301), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1096), .B(new_n1108), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  AND4_X1   g690(.A1(G301), .A2(new_n1101), .A3(new_n1104), .A4(new_n1106), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1116), .B1(new_n1113), .B2(G171), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1115), .B1(new_n1117), .B2(new_n1096), .ZN(new_n1118));
  INV_X1    g693(.A(G1966), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1098), .A2(new_n1119), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT121), .B(G2084), .Z(new_n1121));
  OAI21_X1  g696(.A(new_n1120), .B1(new_n1062), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(G8), .ZN(new_n1123));
  NOR2_X1   g698(.A1(G168), .A2(new_n1038), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1123), .A2(KEYINPUT51), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT51), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1128), .B(G8), .C1(new_n1122), .C2(G286), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1126), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1095), .A2(new_n1118), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1108), .B1(new_n1130), .B2(KEYINPUT62), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(KEYINPUT62), .B2(new_n1130), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1054), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1135));
  NOR2_X1   g710(.A1(G288), .A2(G1976), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  OAI211_X1 g712(.A(KEYINPUT120), .B(new_n1023), .C1(new_n1135), .C2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1137), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1023), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1139), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1138), .A2(G8), .A3(new_n1142), .A4(new_n1017), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1123), .A2(G286), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1037), .A2(new_n1051), .A3(new_n1144), .ZN(new_n1145));
  AOI211_X1 g720(.A(new_n1038), .B(new_n1050), .C1(new_n1042), .C2(new_n1047), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n1145), .A2(KEYINPUT63), .B1(new_n1037), .B2(new_n1146), .ZN(new_n1147));
  OR2_X1    g722(.A1(new_n1145), .A2(KEYINPUT63), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1143), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1015), .B1(new_n1134), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT46), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1005), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1151), .B1(new_n1152), .B2(G1996), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1005), .A2(KEYINPUT46), .A3(new_n706), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1008), .A2(new_n724), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1153), .B(new_n1154), .C1(new_n1152), .C2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1156), .B(KEYINPUT47), .ZN(new_n1157));
  NOR2_X1   g732(.A1(G290), .A2(G1986), .ZN(new_n1158));
  AOI21_X1  g733(.A(KEYINPUT48), .B1(new_n1005), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1159), .B1(new_n1013), .B2(new_n1005), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1005), .A2(KEYINPUT48), .A3(new_n1158), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n837), .A2(new_n839), .ZN(new_n1162));
  OAI22_X1  g737(.A1(new_n1011), .A2(new_n1162), .B1(G2067), .B2(new_n758), .ZN(new_n1163));
  AOI22_X1  g738(.A1(new_n1160), .A2(new_n1161), .B1(new_n1005), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1157), .A2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1165), .B(KEYINPUT127), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1150), .A2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g742(.A1(G227), .A2(new_n461), .ZN(new_n1169));
  NOR3_X1   g743(.A1(G229), .A2(G401), .A3(new_n1169), .ZN(new_n1170));
  AND3_X1   g744(.A1(new_n1170), .A2(new_n994), .A3(new_n906), .ZN(G308));
  NAND3_X1  g745(.A1(new_n1170), .A2(new_n994), .A3(new_n906), .ZN(G225));
endmodule


