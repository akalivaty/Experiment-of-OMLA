

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809;

  BUF_X1 U377 ( .A(n617), .Z(n354) );
  AND2_X1 U378 ( .A1(n443), .A2(n441), .ZN(n437) );
  AND2_X1 U379 ( .A1(n381), .A2(n379), .ZN(n378) );
  NAND2_X1 U380 ( .A1(n388), .A2(n386), .ZN(n606) );
  XNOR2_X1 U381 ( .A(n430), .B(KEYINPUT33), .ZN(n601) );
  XNOR2_X1 U382 ( .A(n736), .B(KEYINPUT6), .ZN(n612) );
  NAND2_X1 U383 ( .A1(n418), .A2(n417), .ZN(n578) );
  OR2_X1 U384 ( .A1(n771), .A2(G902), .ZN(n434) );
  AND2_X1 U385 ( .A1(n412), .A2(n368), .ZN(n359) );
  XNOR2_X1 U386 ( .A(n353), .B(n785), .ZN(n699) );
  XNOR2_X1 U387 ( .A(G110), .B(G107), .ZN(n477) );
  XNOR2_X1 U388 ( .A(G116), .B(G107), .ZN(n521) );
  INV_X2 U389 ( .A(G125), .ZN(n728) );
  XNOR2_X1 U390 ( .A(n373), .B(n485), .ZN(n353) );
  XNOR2_X2 U391 ( .A(n563), .B(n447), .ZN(n798) );
  OR2_X2 U392 ( .A1(n692), .A2(G902), .ZN(n556) );
  NAND2_X1 U393 ( .A1(n605), .A2(n604), .ZN(n749) );
  INV_X1 U394 ( .A(n612), .ZN(n666) );
  XNOR2_X2 U395 ( .A(n529), .B(KEYINPUT4), .ZN(n800) );
  NOR2_X1 U396 ( .A1(n629), .A2(n538), .ZN(n540) );
  NAND2_X1 U397 ( .A1(n425), .A2(n422), .ZN(n657) );
  XNOR2_X1 U398 ( .A(n526), .B(n449), .ZN(n561) );
  XNOR2_X1 U399 ( .A(n540), .B(n468), .ZN(n613) );
  NOR2_X1 U400 ( .A1(n600), .A2(n603), .ZN(n387) );
  AND2_X1 U401 ( .A1(n655), .A2(n746), .ZN(n405) );
  XNOR2_X1 U402 ( .A(n567), .B(n566), .ZN(n599) );
  AND2_X1 U403 ( .A1(n459), .A2(n458), .ZN(n457) );
  NOR2_X1 U404 ( .A1(n768), .A2(n769), .ZN(n415) );
  XNOR2_X1 U405 ( .A(n411), .B(n410), .ZN(n382) );
  NOR2_X1 U406 ( .A1(n400), .A2(n394), .ZN(n393) );
  XNOR2_X1 U407 ( .A(n374), .B(KEYINPUT40), .ZN(n713) );
  NOR2_X1 U408 ( .A1(n387), .A2(n390), .ZN(n386) );
  OR2_X1 U409 ( .A1(n601), .A2(n391), .ZN(n385) );
  NAND2_X1 U410 ( .A1(n599), .A2(n734), .ZN(n608) );
  INV_X1 U411 ( .A(n599), .ZN(n619) );
  XNOR2_X1 U412 ( .A(n477), .B(G104), .ZN(n545) );
  XOR2_X1 U413 ( .A(G137), .B(G140), .Z(n562) );
  XNOR2_X1 U414 ( .A(KEYINPUT16), .B(G122), .ZN(n478) );
  XNOR2_X1 U415 ( .A(G113), .B(KEYINPUT71), .ZN(n473) );
  XNOR2_X1 U416 ( .A(G119), .B(G116), .ZN(n474) );
  XNOR2_X1 U417 ( .A(G128), .B(KEYINPUT23), .ZN(n557) );
  INV_X1 U418 ( .A(n460), .ZN(n355) );
  AND2_X2 U419 ( .A1(n688), .A2(n689), .ZN(n780) );
  BUF_X1 U420 ( .A(n687), .Z(n790) );
  BUF_X1 U421 ( .A(n713), .Z(n356) );
  BUF_X1 U422 ( .A(n627), .Z(n357) );
  INV_X1 U423 ( .A(n619), .ZN(n358) );
  NAND2_X1 U424 ( .A1(n402), .A2(KEYINPUT44), .ZN(n401) );
  INV_X1 U425 ( .A(KEYINPUT66), .ZN(n402) );
  NAND2_X1 U426 ( .A1(n424), .A2(n682), .ZN(n423) );
  INV_X1 U427 ( .A(n490), .ZN(n424) );
  INV_X1 U428 ( .A(KEYINPUT10), .ZN(n448) );
  NAND2_X1 U429 ( .A1(n435), .A2(n790), .ZN(n688) );
  NAND2_X1 U430 ( .A1(n437), .A2(n436), .ZN(n435) );
  NAND2_X1 U431 ( .A1(n397), .A2(n395), .ZN(n394) );
  NAND2_X1 U432 ( .A1(n396), .A2(KEYINPUT66), .ZN(n395) );
  NOR2_X1 U433 ( .A1(G953), .A2(G237), .ZN(n550) );
  XOR2_X1 U434 ( .A(KEYINPUT105), .B(KEYINPUT107), .Z(n510) );
  XNOR2_X1 U435 ( .A(G140), .B(KEYINPUT106), .ZN(n509) );
  XOR2_X1 U436 ( .A(G122), .B(G104), .Z(n508) );
  NAND2_X1 U437 ( .A1(n427), .A2(n426), .ZN(n412) );
  NAND2_X1 U438 ( .A1(n490), .A2(n642), .ZN(n426) );
  NAND2_X1 U439 ( .A1(n699), .A2(n490), .ZN(n427) );
  AND2_X1 U440 ( .A1(n380), .A2(n681), .ZN(n379) );
  NAND2_X1 U441 ( .A1(n679), .A2(KEYINPUT88), .ZN(n380) );
  XNOR2_X1 U442 ( .A(n641), .B(KEYINPUT45), .ZN(n687) );
  OR2_X1 U443 ( .A1(n699), .A2(n423), .ZN(n422) );
  NAND2_X1 U444 ( .A1(n421), .A2(n420), .ZN(n419) );
  NAND2_X1 U445 ( .A1(n594), .A2(KEYINPUT19), .ZN(n420) );
  NAND2_X1 U446 ( .A1(n404), .A2(n368), .ZN(n403) );
  XNOR2_X1 U447 ( .A(n565), .B(KEYINPUT25), .ZN(n566) );
  INV_X1 U448 ( .A(n562), .ZN(n447) );
  INV_X1 U449 ( .A(KEYINPUT8), .ZN(n449) );
  XNOR2_X1 U450 ( .A(n373), .B(n542), .ZN(n549) );
  NOR2_X1 U451 ( .A1(n463), .A2(n784), .ZN(n462) );
  NOR2_X1 U452 ( .A1(n466), .A2(G210), .ZN(n463) );
  NAND2_X1 U453 ( .A1(n780), .A2(n371), .ZN(n464) );
  NAND2_X1 U454 ( .A1(n460), .A2(n703), .ZN(n455) );
  XNOR2_X1 U455 ( .A(n415), .B(KEYINPUT85), .ZN(n429) );
  INV_X1 U456 ( .A(n688), .ZN(n768) );
  INV_X1 U457 ( .A(KEYINPUT44), .ZN(n396) );
  NAND2_X1 U458 ( .A1(n399), .A2(n398), .ZN(n397) );
  INV_X1 U459 ( .A(n401), .ZN(n398) );
  INV_X1 U460 ( .A(KEYINPUT90), .ZN(n634) );
  XOR2_X1 U461 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n482) );
  INV_X1 U462 ( .A(n423), .ZN(n404) );
  XOR2_X1 U463 ( .A(KEYINPUT12), .B(KEYINPUT104), .Z(n504) );
  INV_X1 U464 ( .A(KEYINPUT11), .ZN(n505) );
  XNOR2_X1 U465 ( .A(G113), .B(G143), .ZN(n507) );
  XNOR2_X1 U466 ( .A(KEYINPUT70), .B(G131), .ZN(n541) );
  NAND2_X1 U467 ( .A1(G234), .A2(G237), .ZN(n493) );
  AND2_X1 U468 ( .A1(n439), .A2(KEYINPUT2), .ZN(n438) );
  INV_X1 U469 ( .A(KEYINPUT87), .ZN(n439) );
  NAND2_X1 U470 ( .A1(n442), .A2(KEYINPUT87), .ZN(n441) );
  INV_X1 U471 ( .A(KEYINPUT2), .ZN(n442) );
  NAND2_X1 U472 ( .A1(n666), .A2(n431), .ZN(n430) );
  XNOR2_X1 U473 ( .A(n520), .B(n519), .ZN(n605) );
  XNOR2_X1 U474 ( .A(n433), .B(n432), .ZN(n627) );
  INV_X1 U475 ( .A(KEYINPUT101), .ZN(n432) );
  NAND2_X1 U476 ( .A1(n377), .A2(KEYINPUT88), .ZN(n376) );
  XNOR2_X1 U477 ( .A(KEYINPUT95), .B(KEYINPUT3), .ZN(n475) );
  INV_X1 U478 ( .A(G128), .ZN(n486) );
  XNOR2_X1 U479 ( .A(G134), .B(G122), .ZN(n522) );
  XOR2_X1 U480 ( .A(KEYINPUT109), .B(KEYINPUT7), .Z(n523) );
  INV_X1 U481 ( .A(KEYINPUT84), .ZN(n453) );
  INV_X1 U482 ( .A(n658), .ZN(n390) );
  XNOR2_X1 U483 ( .A(n407), .B(n406), .ZN(n655) );
  NOR2_X1 U484 ( .A1(n419), .A2(n359), .ZN(n418) );
  XNOR2_X1 U485 ( .A(n692), .B(n691), .ZN(n693) );
  XNOR2_X1 U486 ( .A(n451), .B(n450), .ZN(n444) );
  XNOR2_X1 U487 ( .A(n798), .B(n446), .ZN(n445) );
  XNOR2_X1 U488 ( .A(n706), .B(n705), .ZN(n707) );
  NAND2_X1 U489 ( .A1(n613), .A2(n367), .ZN(n467) );
  NOR2_X1 U490 ( .A1(n583), .A2(n582), .ZN(n723) );
  NAND2_X1 U491 ( .A1(n369), .A2(n455), .ZN(n456) );
  INV_X1 U492 ( .A(KEYINPUT53), .ZN(n413) );
  AND2_X1 U493 ( .A1(n770), .A2(n789), .ZN(n428) );
  AND2_X1 U494 ( .A1(n409), .A2(n680), .ZN(n360) );
  AND2_X1 U495 ( .A1(n462), .A2(KEYINPUT56), .ZN(n361) );
  XOR2_X1 U496 ( .A(n555), .B(n554), .Z(n362) );
  XNOR2_X1 U497 ( .A(G119), .B(G110), .ZN(n363) );
  XOR2_X1 U498 ( .A(KEYINPUT99), .B(KEYINPUT24), .Z(n364) );
  AND2_X1 U499 ( .A1(n416), .A2(n633), .ZN(n365) );
  INV_X1 U500 ( .A(n679), .ZN(n409) );
  AND2_X1 U501 ( .A1(n616), .A2(KEYINPUT66), .ZN(n366) );
  NOR2_X1 U502 ( .A1(n614), .A2(n666), .ZN(n367) );
  AND2_X1 U503 ( .A1(n745), .A2(n492), .ZN(n368) );
  AND2_X1 U504 ( .A1(n464), .A2(n361), .ZN(n369) );
  AND2_X1 U505 ( .A1(n422), .A2(KEYINPUT19), .ZN(n370) );
  INV_X1 U506 ( .A(n603), .ZN(n391) );
  AND2_X1 U507 ( .A1(n466), .A2(G210), .ZN(n371) );
  AND2_X1 U508 ( .A1(n703), .A2(n465), .ZN(n372) );
  XNOR2_X1 U509 ( .A(n445), .B(n444), .ZN(n781) );
  INV_X1 U510 ( .A(G953), .ZN(n789) );
  INV_X1 U511 ( .A(KEYINPUT56), .ZN(n465) );
  XNOR2_X2 U512 ( .A(n800), .B(n488), .ZN(n373) );
  NAND2_X1 U513 ( .A1(n644), .A2(n723), .ZN(n374) );
  XNOR2_X2 U514 ( .A(n375), .B(KEYINPUT39), .ZN(n644) );
  NAND2_X2 U515 ( .A1(n656), .A2(n405), .ZN(n375) );
  NAND2_X2 U516 ( .A1(n378), .A2(n376), .ZN(n686) );
  INV_X1 U517 ( .A(n382), .ZN(n377) );
  NAND2_X1 U518 ( .A1(n382), .A2(n360), .ZN(n381) );
  NAND2_X1 U519 ( .A1(n365), .A2(n383), .ZN(n635) );
  NAND2_X1 U520 ( .A1(n393), .A2(n392), .ZN(n383) );
  NOR2_X1 U521 ( .A1(n617), .A2(n401), .ZN(n400) );
  XNOR2_X2 U522 ( .A(n467), .B(KEYINPUT32), .ZN(n617) );
  NAND2_X1 U523 ( .A1(n385), .A2(n384), .ZN(n388) );
  NAND2_X1 U524 ( .A1(n389), .A2(n601), .ZN(n384) );
  NAND2_X1 U525 ( .A1(n600), .A2(n603), .ZN(n389) );
  NAND2_X1 U526 ( .A1(n617), .A2(n616), .ZN(n636) );
  NAND2_X1 U527 ( .A1(n617), .A2(n366), .ZN(n392) );
  INV_X1 U528 ( .A(n616), .ZN(n399) );
  OR2_X1 U529 ( .A1(n699), .A2(n403), .ZN(n421) );
  INV_X1 U530 ( .A(KEYINPUT30), .ZN(n406) );
  NAND2_X1 U531 ( .A1(n736), .A2(n745), .ZN(n407) );
  XNOR2_X2 U532 ( .A(n408), .B(KEYINPUT77), .ZN(n656) );
  NAND2_X1 U533 ( .A1(n627), .A2(n610), .ZN(n408) );
  INV_X1 U534 ( .A(KEYINPUT48), .ZN(n410) );
  NAND2_X1 U535 ( .A1(n678), .A2(n677), .ZN(n411) );
  INV_X1 U536 ( .A(n412), .ZN(n425) );
  XNOR2_X1 U537 ( .A(n414), .B(n413), .ZN(G75) );
  NAND2_X1 U538 ( .A1(n429), .A2(n428), .ZN(n414) );
  NAND2_X1 U539 ( .A1(n637), .A2(KEYINPUT44), .ZN(n416) );
  NOR2_X2 U540 ( .A1(n609), .A2(n608), .ZN(n433) );
  XNOR2_X1 U541 ( .A(n454), .B(n453), .ZN(n452) );
  NOR2_X1 U542 ( .A1(n732), .A2(n608), .ZN(n431) );
  NAND2_X1 U543 ( .A1(n440), .A2(n438), .ZN(n436) );
  NAND2_X1 U544 ( .A1(n370), .A2(n425), .ZN(n417) );
  XNOR2_X2 U545 ( .A(n606), .B(KEYINPUT35), .ZN(n637) );
  INV_X1 U546 ( .A(n601), .ZN(n762) );
  XNOR2_X2 U547 ( .A(n434), .B(n548), .ZN(n609) );
  INV_X1 U548 ( .A(n686), .ZN(n440) );
  NAND2_X1 U549 ( .A1(n686), .A2(KEYINPUT87), .ZN(n443) );
  INV_X1 U550 ( .A(n644), .ZN(n643) );
  NAND2_X1 U551 ( .A1(n561), .A2(G221), .ZN(n446) );
  XNOR2_X2 U552 ( .A(n515), .B(n448), .ZN(n563) );
  XNOR2_X2 U553 ( .A(n728), .B(G146), .ZN(n515) );
  XNOR2_X1 U554 ( .A(n558), .B(KEYINPUT78), .ZN(n450) );
  XNOR2_X1 U555 ( .A(n560), .B(n363), .ZN(n451) );
  NAND2_X1 U556 ( .A1(n452), .A2(n440), .ZN(n685) );
  NAND2_X1 U557 ( .A1(n687), .A2(n642), .ZN(n454) );
  NAND2_X1 U558 ( .A1(n464), .A2(n462), .ZN(n461) );
  NAND2_X1 U559 ( .A1(n457), .A2(n456), .ZN(G51) );
  NAND2_X1 U560 ( .A1(n460), .A2(n372), .ZN(n458) );
  NAND2_X1 U561 ( .A1(n461), .A2(n465), .ZN(n459) );
  INV_X1 U562 ( .A(n780), .ZN(n460) );
  INV_X1 U563 ( .A(n703), .ZN(n466) );
  NAND2_X1 U564 ( .A1(n613), .A2(n612), .ZN(n618) );
  XNOR2_X1 U565 ( .A(n549), .B(n362), .ZN(n692) );
  NAND2_X1 U566 ( .A1(n685), .A2(n471), .ZN(n689) );
  OR2_X1 U567 ( .A1(n806), .A2(G952), .ZN(n709) );
  XOR2_X1 U568 ( .A(n539), .B(KEYINPUT74), .Z(n468) );
  OR2_X1 U569 ( .A1(G237), .A2(G902), .ZN(n469) );
  NAND2_X1 U570 ( .A1(n501), .A2(n500), .ZN(n470) );
  XNOR2_X1 U571 ( .A(KEYINPUT68), .B(n684), .ZN(n471) );
  NAND2_X1 U572 ( .A1(n639), .A2(n638), .ZN(n472) );
  XNOR2_X1 U573 ( .A(n506), .B(n505), .ZN(n514) );
  INV_X1 U574 ( .A(G475), .ZN(n518) );
  XNOR2_X1 U575 ( .A(n514), .B(n513), .ZN(n517) );
  XNOR2_X1 U576 ( .A(n518), .B(KEYINPUT13), .ZN(n519) );
  XNOR2_X1 U577 ( .A(n474), .B(n473), .ZN(n476) );
  XNOR2_X1 U578 ( .A(n476), .B(n475), .ZN(n555) );
  XNOR2_X1 U579 ( .A(n545), .B(n478), .ZN(n479) );
  XNOR2_X1 U580 ( .A(n555), .B(n479), .ZN(n785) );
  INV_X1 U581 ( .A(KEYINPUT64), .ZN(n480) );
  XNOR2_X2 U582 ( .A(n480), .B(G953), .ZN(n806) );
  NAND2_X1 U583 ( .A1(n806), .A2(G224), .ZN(n481) );
  XNOR2_X1 U584 ( .A(n482), .B(n481), .ZN(n484) );
  XNOR2_X1 U585 ( .A(n515), .B(KEYINPUT79), .ZN(n483) );
  XNOR2_X1 U586 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X2 U587 ( .A(KEYINPUT65), .B(G143), .ZN(n487) );
  XNOR2_X2 U588 ( .A(n487), .B(n486), .ZN(n529) );
  XNOR2_X1 U589 ( .A(KEYINPUT69), .B(G101), .ZN(n488) );
  XNOR2_X1 U590 ( .A(G902), .B(KEYINPUT15), .ZN(n682) );
  INV_X1 U591 ( .A(n682), .ZN(n642) );
  XNOR2_X1 U592 ( .A(KEYINPUT76), .B(n469), .ZN(n491) );
  AND2_X1 U593 ( .A1(n491), .A2(G210), .ZN(n490) );
  AND2_X1 U594 ( .A1(n491), .A2(G214), .ZN(n594) );
  INV_X1 U595 ( .A(n594), .ZN(n745) );
  INV_X1 U596 ( .A(KEYINPUT19), .ZN(n492) );
  NOR2_X1 U597 ( .A1(G898), .A2(n789), .ZN(n787) );
  NAND2_X1 U598 ( .A1(G902), .A2(n787), .ZN(n496) );
  NOR2_X1 U599 ( .A1(KEYINPUT96), .A2(n496), .ZN(n499) );
  XNOR2_X1 U600 ( .A(n493), .B(KEYINPUT14), .ZN(n731) );
  NAND2_X1 U601 ( .A1(n499), .A2(n731), .ZN(n495) );
  INV_X1 U602 ( .A(KEYINPUT96), .ZN(n494) );
  NAND2_X1 U603 ( .A1(n495), .A2(n494), .ZN(n501) );
  NAND2_X1 U604 ( .A1(G952), .A2(n789), .ZN(n571) );
  NAND2_X1 U605 ( .A1(n571), .A2(n496), .ZN(n497) );
  NAND2_X1 U606 ( .A1(n731), .A2(n497), .ZN(n498) );
  OR2_X1 U607 ( .A1(n499), .A2(n498), .ZN(n500) );
  NAND2_X1 U608 ( .A1(n578), .A2(n470), .ZN(n502) );
  XNOR2_X2 U609 ( .A(n502), .B(KEYINPUT0), .ZN(n629) );
  NAND2_X1 U610 ( .A1(G214), .A2(n550), .ZN(n503) );
  XNOR2_X1 U611 ( .A(n504), .B(n503), .ZN(n506) );
  XNOR2_X1 U612 ( .A(n508), .B(n507), .ZN(n512) );
  XNOR2_X1 U613 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U614 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U615 ( .A(n541), .B(n563), .Z(n516) );
  XNOR2_X1 U616 ( .A(n517), .B(n516), .ZN(n706) );
  NOR2_X1 U617 ( .A1(G902), .A2(n706), .ZN(n520) );
  XNOR2_X1 U618 ( .A(n521), .B(KEYINPUT9), .ZN(n525) );
  XNOR2_X1 U619 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U620 ( .A(n525), .B(n524), .Z(n528) );
  NAND2_X1 U621 ( .A1(n806), .A2(G234), .ZN(n526) );
  NAND2_X1 U622 ( .A1(G217), .A2(n561), .ZN(n527) );
  XNOR2_X1 U623 ( .A(n528), .B(n527), .ZN(n530) );
  XNOR2_X1 U624 ( .A(n529), .B(n530), .ZN(n778) );
  INV_X1 U625 ( .A(G902), .ZN(n531) );
  NAND2_X1 U626 ( .A1(n778), .A2(n531), .ZN(n532) );
  XNOR2_X1 U627 ( .A(n532), .B(G478), .ZN(n582) );
  INV_X1 U628 ( .A(n582), .ZN(n604) );
  INV_X1 U629 ( .A(n749), .ZN(n536) );
  NAND2_X1 U630 ( .A1(G234), .A2(n682), .ZN(n533) );
  XNOR2_X1 U631 ( .A(KEYINPUT20), .B(n533), .ZN(n564) );
  NAND2_X1 U632 ( .A1(n564), .A2(G221), .ZN(n535) );
  INV_X1 U633 ( .A(KEYINPUT21), .ZN(n534) );
  XNOR2_X1 U634 ( .A(n535), .B(n534), .ZN(n734) );
  NAND2_X1 U635 ( .A1(n536), .A2(n734), .ZN(n537) );
  XNOR2_X1 U636 ( .A(n537), .B(KEYINPUT110), .ZN(n538) );
  XNOR2_X1 U637 ( .A(KEYINPUT75), .B(KEYINPUT22), .ZN(n539) );
  XNOR2_X1 U638 ( .A(n541), .B(G134), .ZN(n799) );
  XNOR2_X1 U639 ( .A(n799), .B(G146), .ZN(n542) );
  NAND2_X1 U640 ( .A1(n806), .A2(G227), .ZN(n544) );
  XNOR2_X1 U641 ( .A(KEYINPUT97), .B(n562), .ZN(n543) );
  XNOR2_X1 U642 ( .A(n544), .B(n543), .ZN(n546) );
  XNOR2_X1 U643 ( .A(n545), .B(n546), .ZN(n547) );
  XNOR2_X1 U644 ( .A(n549), .B(n547), .ZN(n771) );
  INV_X1 U645 ( .A(G469), .ZN(n548) );
  XNOR2_X1 U646 ( .A(n609), .B(KEYINPUT1), .ZN(n732) );
  INV_X1 U647 ( .A(n732), .ZN(n623) );
  NAND2_X1 U648 ( .A1(n550), .A2(G210), .ZN(n551) );
  XNOR2_X1 U649 ( .A(n551), .B(G137), .ZN(n553) );
  XNOR2_X1 U650 ( .A(KEYINPUT102), .B(KEYINPUT5), .ZN(n552) );
  XNOR2_X1 U651 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X2 U652 ( .A(n556), .B(G472), .ZN(n736) );
  INV_X1 U653 ( .A(n736), .ZN(n626) );
  XNOR2_X1 U654 ( .A(n557), .B(KEYINPUT100), .ZN(n558) );
  XNOR2_X1 U655 ( .A(KEYINPUT72), .B(KEYINPUT98), .ZN(n559) );
  XNOR2_X1 U656 ( .A(n364), .B(n559), .ZN(n560) );
  NOR2_X1 U657 ( .A1(n781), .A2(G902), .ZN(n567) );
  NAND2_X1 U658 ( .A1(G217), .A2(n564), .ZN(n565) );
  NAND2_X1 U659 ( .A1(n626), .A2(n619), .ZN(n568) );
  NOR2_X1 U660 ( .A1(n623), .A2(n568), .ZN(n569) );
  NAND2_X1 U661 ( .A1(n613), .A2(n569), .ZN(n616) );
  XNOR2_X1 U662 ( .A(n616), .B(G110), .ZN(G12) );
  NOR2_X1 U663 ( .A1(G900), .A2(n806), .ZN(n570) );
  NAND2_X1 U664 ( .A1(G902), .A2(n570), .ZN(n572) );
  NAND2_X1 U665 ( .A1(n572), .A2(n571), .ZN(n573) );
  AND2_X1 U666 ( .A1(n573), .A2(n731), .ZN(n610) );
  NAND2_X1 U667 ( .A1(n734), .A2(n610), .ZN(n574) );
  NOR2_X1 U668 ( .A1(n574), .A2(n358), .ZN(n575) );
  NAND2_X1 U669 ( .A1(n736), .A2(n575), .ZN(n576) );
  XNOR2_X1 U670 ( .A(n576), .B(KEYINPUT28), .ZN(n577) );
  OR2_X1 U671 ( .A1(n577), .A2(n609), .ZN(n596) );
  INV_X1 U672 ( .A(n596), .ZN(n579) );
  AND2_X1 U673 ( .A1(n578), .A2(n579), .ZN(n672) );
  XNOR2_X1 U674 ( .A(n605), .B(KEYINPUT108), .ZN(n583) );
  AND2_X1 U675 ( .A1(n583), .A2(n582), .ZN(n725) );
  NAND2_X1 U676 ( .A1(n672), .A2(n725), .ZN(n581) );
  XOR2_X1 U677 ( .A(G128), .B(KEYINPUT29), .Z(n580) );
  XNOR2_X1 U678 ( .A(n581), .B(n580), .ZN(G30) );
  NAND2_X1 U679 ( .A1(n723), .A2(n672), .ZN(n584) );
  XNOR2_X1 U680 ( .A(n584), .B(G146), .ZN(G48) );
  INV_X1 U681 ( .A(n610), .ZN(n585) );
  NOR2_X1 U682 ( .A1(n585), .A2(n594), .ZN(n586) );
  NAND2_X1 U683 ( .A1(n734), .A2(n586), .ZN(n587) );
  NOR2_X1 U684 ( .A1(n587), .A2(n358), .ZN(n588) );
  NAND2_X1 U685 ( .A1(n723), .A2(n588), .ZN(n665) );
  NOR2_X1 U686 ( .A1(n665), .A2(n623), .ZN(n589) );
  NAND2_X1 U687 ( .A1(n589), .A2(n666), .ZN(n592) );
  INV_X1 U688 ( .A(KEYINPUT111), .ZN(n590) );
  XNOR2_X1 U689 ( .A(n590), .B(KEYINPUT43), .ZN(n591) );
  XNOR2_X1 U690 ( .A(n592), .B(n591), .ZN(n593) );
  INV_X1 U691 ( .A(n657), .ZN(n664) );
  AND2_X1 U692 ( .A1(n593), .A2(n664), .ZN(n679) );
  XOR2_X1 U693 ( .A(G140), .B(n679), .Z(G42) );
  XNOR2_X1 U694 ( .A(n657), .B(KEYINPUT38), .ZN(n607) );
  OR2_X1 U695 ( .A1(n607), .A2(n594), .ZN(n750) );
  NOR2_X1 U696 ( .A1(n750), .A2(n749), .ZN(n595) );
  XNOR2_X1 U697 ( .A(n595), .B(KEYINPUT41), .ZN(n761) );
  OR2_X1 U698 ( .A1(n761), .A2(n596), .ZN(n598) );
  XNOR2_X1 U699 ( .A(KEYINPUT112), .B(KEYINPUT42), .ZN(n597) );
  XNOR2_X1 U700 ( .A(n598), .B(n597), .ZN(n645) );
  XNOR2_X1 U701 ( .A(n645), .B(G137), .ZN(G39) );
  INV_X1 U702 ( .A(n629), .ZN(n600) );
  XNOR2_X1 U703 ( .A(KEYINPUT80), .B(KEYINPUT34), .ZN(n602) );
  XNOR2_X1 U704 ( .A(n602), .B(KEYINPUT73), .ZN(n603) );
  NOR2_X1 U705 ( .A1(n605), .A2(n604), .ZN(n658) );
  XOR2_X1 U706 ( .A(n637), .B(G122), .Z(G24) );
  INV_X1 U707 ( .A(n607), .ZN(n746) );
  INV_X1 U708 ( .A(n725), .ZN(n611) );
  OR2_X1 U709 ( .A1(n643), .A2(n611), .ZN(n681) );
  XNOR2_X1 U710 ( .A(n681), .B(G134), .ZN(G36) );
  NAND2_X1 U711 ( .A1(n623), .A2(n619), .ZN(n614) );
  XNOR2_X1 U712 ( .A(G119), .B(KEYINPUT126), .ZN(n615) );
  XNOR2_X1 U713 ( .A(n354), .B(n615), .ZN(G21) );
  XNOR2_X1 U714 ( .A(n618), .B(KEYINPUT89), .ZN(n621) );
  NOR2_X1 U715 ( .A1(n623), .A2(n619), .ZN(n620) );
  NAND2_X1 U716 ( .A1(n621), .A2(n620), .ZN(n714) );
  NOR2_X1 U717 ( .A1(n626), .A2(n608), .ZN(n622) );
  NAND2_X1 U718 ( .A1(n623), .A2(n622), .ZN(n740) );
  NOR2_X1 U719 ( .A1(n629), .A2(n740), .ZN(n625) );
  XNOR2_X1 U720 ( .A(KEYINPUT103), .B(KEYINPUT31), .ZN(n624) );
  XNOR2_X1 U721 ( .A(n625), .B(n624), .ZN(n726) );
  INV_X1 U722 ( .A(n726), .ZN(n630) );
  NAND2_X1 U723 ( .A1(n357), .A2(n626), .ZN(n628) );
  OR2_X1 U724 ( .A1(n629), .A2(n628), .ZN(n715) );
  NAND2_X1 U725 ( .A1(n630), .A2(n715), .ZN(n631) );
  OR2_X1 U726 ( .A1(n725), .A2(n723), .ZN(n671) );
  NAND2_X1 U727 ( .A1(n631), .A2(n671), .ZN(n632) );
  AND2_X1 U728 ( .A1(n714), .A2(n632), .ZN(n633) );
  XNOR2_X1 U729 ( .A(n635), .B(n634), .ZN(n640) );
  XNOR2_X1 U730 ( .A(n636), .B(KEYINPUT91), .ZN(n639) );
  NOR2_X1 U731 ( .A1(n637), .A2(KEYINPUT44), .ZN(n638) );
  NAND2_X1 U732 ( .A1(n640), .A2(n472), .ZN(n641) );
  NAND2_X1 U733 ( .A1(n713), .A2(n645), .ZN(n647) );
  INV_X1 U734 ( .A(KEYINPUT46), .ZN(n646) );
  XNOR2_X1 U735 ( .A(n647), .B(n646), .ZN(n678) );
  INV_X1 U736 ( .A(n671), .ZN(n751) );
  AND2_X1 U737 ( .A1(KEYINPUT83), .A2(KEYINPUT47), .ZN(n648) );
  NAND2_X1 U738 ( .A1(n751), .A2(n648), .ZN(n650) );
  INV_X1 U739 ( .A(KEYINPUT83), .ZN(n652) );
  NAND2_X1 U740 ( .A1(n671), .A2(n652), .ZN(n649) );
  NAND2_X1 U741 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U742 ( .A1(n651), .A2(n672), .ZN(n654) );
  INV_X1 U743 ( .A(KEYINPUT47), .ZN(n670) );
  NAND2_X1 U744 ( .A1(n652), .A2(n670), .ZN(n653) );
  NAND2_X1 U745 ( .A1(n654), .A2(n653), .ZN(n662) );
  AND2_X1 U746 ( .A1(n656), .A2(n655), .ZN(n660) );
  AND2_X1 U747 ( .A1(n658), .A2(n657), .ZN(n659) );
  AND2_X1 U748 ( .A1(n660), .A2(n659), .ZN(n722) );
  INV_X1 U749 ( .A(n722), .ZN(n661) );
  NAND2_X1 U750 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U751 ( .A(n663), .B(KEYINPUT82), .ZN(n676) );
  NOR2_X1 U752 ( .A1(n665), .A2(n664), .ZN(n667) );
  NAND2_X1 U753 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U754 ( .A(n668), .B(KEYINPUT36), .ZN(n669) );
  OR2_X1 U755 ( .A1(n669), .A2(n732), .ZN(n729) );
  AND2_X1 U756 ( .A1(n671), .A2(n670), .ZN(n673) );
  NAND2_X1 U757 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U758 ( .A1(n729), .A2(n674), .ZN(n675) );
  NOR2_X1 U759 ( .A1(n676), .A2(n675), .ZN(n677) );
  INV_X1 U760 ( .A(KEYINPUT88), .ZN(n680) );
  XOR2_X1 U761 ( .A(KEYINPUT86), .B(n682), .Z(n683) );
  NAND2_X1 U762 ( .A1(n683), .A2(KEYINPUT2), .ZN(n684) );
  NAND2_X1 U763 ( .A1(n780), .A2(G472), .ZN(n694) );
  XOR2_X1 U764 ( .A(KEYINPUT93), .B(KEYINPUT113), .Z(n690) );
  XNOR2_X1 U765 ( .A(n690), .B(KEYINPUT62), .ZN(n691) );
  XNOR2_X1 U766 ( .A(n694), .B(n693), .ZN(n695) );
  NAND2_X1 U767 ( .A1(n695), .A2(n709), .ZN(n698) );
  XNOR2_X1 U768 ( .A(KEYINPUT114), .B(KEYINPUT63), .ZN(n696) );
  XNOR2_X1 U769 ( .A(n696), .B(KEYINPUT94), .ZN(n697) );
  XNOR2_X1 U770 ( .A(n698), .B(n697), .ZN(G57) );
  XOR2_X1 U771 ( .A(KEYINPUT55), .B(KEYINPUT54), .Z(n701) );
  XNOR2_X1 U772 ( .A(KEYINPUT92), .B(KEYINPUT81), .ZN(n700) );
  XOR2_X1 U773 ( .A(n701), .B(n700), .Z(n702) );
  XNOR2_X1 U774 ( .A(n699), .B(n702), .ZN(n703) );
  INV_X1 U775 ( .A(n709), .ZN(n784) );
  NAND2_X1 U776 ( .A1(n780), .A2(G475), .ZN(n708) );
  XNOR2_X1 U777 ( .A(KEYINPUT67), .B(KEYINPUT121), .ZN(n704) );
  XNOR2_X1 U778 ( .A(n704), .B(KEYINPUT59), .ZN(n705) );
  XNOR2_X1 U779 ( .A(n708), .B(n707), .ZN(n710) );
  NAND2_X1 U780 ( .A1(n710), .A2(n709), .ZN(n712) );
  XOR2_X1 U781 ( .A(KEYINPUT122), .B(KEYINPUT60), .Z(n711) );
  XNOR2_X1 U782 ( .A(n712), .B(n711), .ZN(G60) );
  XNOR2_X1 U783 ( .A(n356), .B(G131), .ZN(G33) );
  XNOR2_X1 U784 ( .A(G101), .B(n714), .ZN(G3) );
  XOR2_X1 U785 ( .A(G104), .B(KEYINPUT115), .Z(n717) );
  INV_X1 U786 ( .A(n715), .ZN(n718) );
  NAND2_X1 U787 ( .A1(n718), .A2(n723), .ZN(n716) );
  XNOR2_X1 U788 ( .A(n717), .B(n716), .ZN(G6) );
  XOR2_X1 U789 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n720) );
  NAND2_X1 U790 ( .A1(n718), .A2(n725), .ZN(n719) );
  XNOR2_X1 U791 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X1 U792 ( .A(G107), .B(n721), .ZN(G9) );
  XOR2_X1 U793 ( .A(G143), .B(n722), .Z(G45) );
  NAND2_X1 U794 ( .A1(n726), .A2(n723), .ZN(n724) );
  XNOR2_X1 U795 ( .A(n724), .B(G113), .ZN(G15) );
  NAND2_X1 U796 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U797 ( .A(n727), .B(G116), .ZN(G18) );
  XNOR2_X1 U798 ( .A(n729), .B(n728), .ZN(n730) );
  XNOR2_X1 U799 ( .A(n730), .B(KEYINPUT37), .ZN(G27) );
  NAND2_X1 U800 ( .A1(G952), .A2(n731), .ZN(n760) );
  XOR2_X1 U801 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n743) );
  NAND2_X1 U802 ( .A1(n732), .A2(n608), .ZN(n733) );
  XNOR2_X1 U803 ( .A(n733), .B(KEYINPUT50), .ZN(n739) );
  NOR2_X1 U804 ( .A1(n734), .A2(n358), .ZN(n735) );
  XOR2_X1 U805 ( .A(KEYINPUT49), .B(n735), .Z(n737) );
  NOR2_X1 U806 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U807 ( .A1(n739), .A2(n738), .ZN(n741) );
  NAND2_X1 U808 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U809 ( .A(n743), .B(n742), .Z(n744) );
  NOR2_X1 U810 ( .A1(n744), .A2(n761), .ZN(n757) );
  NOR2_X1 U811 ( .A1(n746), .A2(n745), .ZN(n747) );
  XOR2_X1 U812 ( .A(KEYINPUT117), .B(n747), .Z(n748) );
  NOR2_X1 U813 ( .A1(n749), .A2(n748), .ZN(n754) );
  NOR2_X1 U814 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U815 ( .A(n752), .B(KEYINPUT118), .ZN(n753) );
  NOR2_X1 U816 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U817 ( .A1(n755), .A2(n762), .ZN(n756) );
  NOR2_X1 U818 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U819 ( .A(n758), .B(KEYINPUT52), .ZN(n759) );
  NOR2_X1 U820 ( .A1(n760), .A2(n759), .ZN(n764) );
  NOR2_X1 U821 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U822 ( .A1(n764), .A2(n763), .ZN(n765) );
  XOR2_X1 U823 ( .A(KEYINPUT119), .B(n765), .Z(n770) );
  INV_X1 U824 ( .A(n790), .ZN(n766) );
  NOR2_X1 U825 ( .A1(n766), .A2(n686), .ZN(n767) );
  NOR2_X1 U826 ( .A1(n767), .A2(KEYINPUT2), .ZN(n769) );
  NAND2_X1 U827 ( .A1(n355), .A2(G469), .ZN(n775) );
  XNOR2_X1 U828 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n772) );
  XOR2_X1 U829 ( .A(n772), .B(KEYINPUT57), .Z(n773) );
  XNOR2_X1 U830 ( .A(n771), .B(n773), .ZN(n774) );
  XNOR2_X1 U831 ( .A(n775), .B(n774), .ZN(n776) );
  NOR2_X1 U832 ( .A1(n784), .A2(n776), .ZN(G54) );
  NAND2_X1 U833 ( .A1(n780), .A2(G478), .ZN(n777) );
  XOR2_X1 U834 ( .A(n778), .B(n777), .Z(n779) );
  NOR2_X1 U835 ( .A1(n784), .A2(n779), .ZN(G63) );
  NAND2_X1 U836 ( .A1(n780), .A2(G217), .ZN(n782) );
  XNOR2_X1 U837 ( .A(n781), .B(n782), .ZN(n783) );
  NOR2_X1 U838 ( .A1(n784), .A2(n783), .ZN(G66) );
  XNOR2_X1 U839 ( .A(G101), .B(KEYINPUT124), .ZN(n786) );
  XNOR2_X1 U840 ( .A(n785), .B(n786), .ZN(n788) );
  NOR2_X1 U841 ( .A1(n788), .A2(n787), .ZN(n797) );
  NAND2_X1 U842 ( .A1(n790), .A2(n789), .ZN(n795) );
  XOR2_X1 U843 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n792) );
  NAND2_X1 U844 ( .A1(G224), .A2(G953), .ZN(n791) );
  XNOR2_X1 U845 ( .A(n792), .B(n791), .ZN(n793) );
  NAND2_X1 U846 ( .A1(n793), .A2(G898), .ZN(n794) );
  NAND2_X1 U847 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U848 ( .A(n797), .B(n796), .ZN(G69) );
  XOR2_X1 U849 ( .A(KEYINPUT125), .B(n798), .Z(n802) );
  XNOR2_X1 U850 ( .A(n800), .B(n799), .ZN(n801) );
  XNOR2_X1 U851 ( .A(n802), .B(n801), .ZN(n805) );
  XOR2_X1 U852 ( .A(G227), .B(n805), .Z(n803) );
  NAND2_X1 U853 ( .A1(G900), .A2(n803), .ZN(n804) );
  NAND2_X1 U854 ( .A1(n804), .A2(G953), .ZN(n809) );
  XOR2_X1 U855 ( .A(n805), .B(n686), .Z(n807) );
  NAND2_X1 U856 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U857 ( .A1(n809), .A2(n808), .ZN(G72) );
endmodule

