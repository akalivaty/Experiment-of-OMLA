//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 1 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 1 0 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n209), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  OR2_X1    g0020(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n212), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n223), .A2(new_n207), .ZN(new_n224));
  OAI21_X1  g0024(.A(G50), .B1(G58), .B2(G68), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT64), .Z(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT65), .Z(new_n227));
  AOI21_X1  g0027(.A(new_n222), .B1(new_n224), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G87), .B(G97), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  NOR2_X1   g0043(.A1(G223), .A2(G1698), .ZN(new_n244));
  INV_X1    g0044(.A(G226), .ZN(new_n245));
  AOI21_X1  g0045(.A(new_n244), .B1(new_n245), .B2(G1698), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT3), .B(G33), .ZN(new_n247));
  AOI22_X1  g0047(.A1(new_n246), .A2(new_n247), .B1(G33), .B2(G87), .ZN(new_n248));
  NAND2_X1  g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(G1), .A3(G13), .ZN(new_n250));
  OAI21_X1  g0050(.A(KEYINPUT74), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT66), .ZN(new_n252));
  AND2_X1   g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  OAI21_X1  g0053(.A(G274), .B1(new_n253), .B2(new_n223), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n252), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G274), .ZN(new_n257));
  AND2_X1   g0057(.A1(G1), .A2(G13), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n257), .B1(new_n258), .B2(new_n249), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  INV_X1    g0060(.A(G45), .ZN(new_n261));
  AOI21_X1  g0061(.A(G1), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n259), .A2(KEYINPUT66), .A3(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n253), .A2(new_n223), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(new_n262), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n256), .A2(new_n263), .B1(new_n265), .B2(G232), .ZN(new_n266));
  INV_X1    g0066(.A(G190), .ZN(new_n267));
  INV_X1    g0067(.A(new_n244), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT3), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G33), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT3), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n245), .A2(G1698), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n268), .A2(new_n270), .A3(new_n272), .A4(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G87), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT74), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(new_n277), .A3(new_n264), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n251), .A2(new_n266), .A3(new_n267), .A4(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G200), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n265), .A2(G232), .ZN(new_n281));
  NOR3_X1   g0081(.A1(new_n254), .A2(new_n252), .A3(new_n255), .ZN(new_n282));
  AOI21_X1  g0082(.A(KEYINPUT66), .B1(new_n259), .B2(new_n262), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n248), .A2(new_n250), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n280), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n279), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(G58), .B(G68), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n288), .A2(G20), .B1(G159), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n207), .A2(KEYINPUT7), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n291), .B1(new_n270), .B2(new_n272), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n271), .A2(KEYINPUT3), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n269), .A2(G33), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n207), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT7), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n292), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G68), .ZN(new_n298));
  OAI211_X1 g0098(.A(KEYINPUT16), .B(new_n290), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n223), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n288), .A2(G20), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n289), .A2(G159), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT73), .ZN(new_n305));
  AND3_X1   g0105(.A1(new_n270), .A2(new_n272), .A3(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n296), .A2(G20), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n307), .B1(new_n270), .B2(new_n305), .ZN(new_n308));
  AOI21_X1  g0108(.A(G20), .B1(new_n270), .B2(new_n272), .ZN(new_n309));
  OAI22_X1  g0109(.A1(new_n306), .A2(new_n308), .B1(new_n309), .B2(KEYINPUT7), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n304), .B1(new_n310), .B2(G68), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n299), .B(new_n301), .C1(new_n311), .C2(KEYINPUT16), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n206), .A2(G20), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT68), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n313), .B(new_n314), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT8), .B(G58), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G13), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n318), .A2(new_n207), .A3(G1), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(new_n301), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n317), .A2(new_n320), .B1(new_n316), .B2(new_n319), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n287), .A2(new_n312), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT17), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n321), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n310), .A2(G68), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n290), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT16), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n301), .ZN(new_n330));
  OAI22_X1  g0130(.A1(new_n309), .A2(KEYINPUT7), .B1(new_n247), .B2(new_n291), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n304), .B1(new_n331), .B2(G68), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n330), .B1(new_n332), .B2(KEYINPUT16), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n325), .B1(new_n329), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n334), .A2(KEYINPUT17), .A3(new_n287), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n324), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n299), .A2(new_n301), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT16), .B1(new_n326), .B2(new_n290), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n321), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n277), .B1(new_n276), .B2(new_n264), .ZN(new_n340));
  AOI211_X1 g0140(.A(KEYINPUT74), .B(new_n250), .C1(new_n274), .C2(new_n275), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n256), .A2(new_n263), .ZN(new_n343));
  INV_X1    g0143(.A(G179), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n343), .A2(new_n344), .A3(new_n281), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n343), .B(new_n281), .C1(new_n250), .C2(new_n248), .ZN(new_n346));
  INV_X1    g0146(.A(G169), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n342), .A2(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT18), .B1(new_n339), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n339), .A2(new_n348), .A3(KEYINPUT18), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n349), .B1(KEYINPUT75), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT75), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n339), .A2(new_n348), .A3(new_n352), .A4(KEYINPUT18), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n336), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n289), .A2(G50), .B1(G20), .B2(new_n298), .ZN(new_n355));
  INV_X1    g0155(.A(G77), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n207), .A2(G33), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n358), .A2(new_n301), .ZN(new_n359));
  OR2_X1    g0159(.A1(new_n359), .A2(KEYINPUT11), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n318), .A2(G1), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G20), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n330), .A2(new_n362), .A3(KEYINPUT70), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT70), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n319), .B2(new_n301), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n315), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(G68), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n319), .A2(new_n298), .ZN(new_n369));
  XNOR2_X1  g0169(.A(new_n369), .B(KEYINPUT12), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n359), .A2(KEYINPUT11), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n360), .A2(new_n368), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT14), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT13), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G33), .A2(G97), .ZN(new_n375));
  INV_X1    g0175(.A(G232), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G1698), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(G226), .B2(G1698), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n270), .A2(new_n272), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n375), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n256), .A2(new_n263), .B1(new_n380), .B2(new_n264), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT67), .ZN(new_n382));
  AND3_X1   g0182(.A1(new_n250), .A2(new_n382), .A3(new_n255), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n382), .B1(new_n250), .B2(new_n255), .ZN(new_n384));
  OAI21_X1  g0184(.A(G238), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n374), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n380), .A2(new_n264), .ZN(new_n387));
  AND4_X1   g0187(.A1(new_n374), .A2(new_n385), .A3(new_n343), .A4(new_n387), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n373), .B(G169), .C1(new_n386), .C2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n385), .A2(new_n343), .A3(new_n387), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT13), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n381), .A2(new_n374), .A3(new_n385), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n391), .A2(new_n392), .A3(G179), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n391), .A2(new_n392), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n373), .B1(new_n395), .B2(G169), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n372), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n395), .A2(G200), .ZN(new_n398));
  INV_X1    g0198(.A(new_n372), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n398), .B(new_n399), .C1(new_n267), .C2(new_n395), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n354), .A2(new_n402), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n383), .A2(new_n384), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(G226), .ZN(new_n405));
  NOR2_X1   g0205(.A1(G222), .A2(G1698), .ZN(new_n406));
  INV_X1    g0206(.A(G1698), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n407), .A2(G223), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n247), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n409), .B(new_n264), .C1(G77), .C2(new_n247), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n405), .A2(new_n343), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n347), .ZN(new_n412));
  INV_X1    g0212(.A(G50), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n315), .A2(new_n413), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(new_n320), .B1(new_n413), .B2(new_n319), .ZN(new_n415));
  INV_X1    g0215(.A(G150), .ZN(new_n416));
  INV_X1    g0216(.A(new_n289), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n316), .A2(new_n357), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(G58), .A2(G68), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n207), .B1(new_n419), .B2(new_n413), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n301), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n415), .A2(new_n421), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n412), .B(new_n422), .C1(G179), .C2(new_n411), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT71), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT9), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n415), .A2(new_n426), .A3(new_n421), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n426), .B1(new_n415), .B2(new_n421), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n425), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n429), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n431), .A2(KEYINPUT71), .A3(new_n427), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n411), .A2(G200), .ZN(new_n433));
  INV_X1    g0233(.A(new_n411), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT10), .B1(new_n434), .B2(G190), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n430), .A2(new_n432), .A3(new_n433), .A4(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n433), .B1(new_n267), .B2(new_n411), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n428), .A2(new_n429), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT10), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n424), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(G87), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT15), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT15), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G87), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(new_n357), .ZN(new_n446));
  OAI22_X1  g0246(.A1(new_n316), .A2(new_n417), .B1(new_n207), .B2(new_n356), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n301), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT69), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n448), .B(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n366), .A2(G77), .A3(new_n367), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(G77), .B2(new_n362), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n404), .A2(G244), .ZN(new_n454));
  NOR2_X1   g0254(.A1(G232), .A2(G1698), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n407), .A2(G238), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n247), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n457), .B(new_n264), .C1(G107), .C2(new_n247), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n454), .A2(new_n343), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G200), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n453), .B(new_n460), .C1(new_n267), .C2(new_n459), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n459), .A2(new_n347), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n454), .A2(new_n344), .A3(new_n343), .A4(new_n458), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n462), .B(new_n463), .C1(new_n450), .C2(new_n452), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n440), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT72), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT72), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n440), .A2(new_n468), .A3(new_n465), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n403), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT79), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n407), .A2(G238), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n379), .B2(new_n473), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n247), .A2(KEYINPUT79), .A3(G238), .A4(new_n407), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G116), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n270), .A2(new_n272), .A3(G244), .A4(G1698), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT80), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT80), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n247), .A2(new_n480), .A3(G244), .A4(G1698), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n264), .B1(new_n477), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G250), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n261), .A2(G1), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n264), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n486), .B1(new_n259), .B2(new_n485), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n483), .A2(new_n344), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT81), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n483), .A2(new_n487), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n347), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT82), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT19), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n207), .B1(new_n375), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n441), .A2(new_n202), .A3(new_n203), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n270), .A2(new_n272), .A3(new_n207), .A4(G68), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n493), .B1(new_n357), .B2(new_n202), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n301), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n442), .A2(new_n444), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n362), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n492), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  AOI211_X1 g0304(.A(KEYINPUT82), .B(new_n502), .C1(new_n499), .C2(new_n301), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n320), .B1(G1), .B2(new_n271), .ZN(new_n506));
  OAI22_X1  g0306(.A1(new_n504), .A2(new_n505), .B1(new_n445), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT81), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n483), .A2(new_n508), .A3(new_n344), .A4(new_n487), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n489), .A2(new_n491), .A3(new_n507), .A4(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n270), .A2(new_n272), .A3(G244), .A4(new_n407), .ZN(new_n511));
  XOR2_X1   g0311(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT4), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n515), .A2(G1698), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n516), .A2(new_n270), .A3(new_n272), .A4(G244), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n270), .A2(new_n272), .A3(G250), .A4(G1698), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G283), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n264), .B1(new_n514), .B2(new_n520), .ZN(new_n521));
  AND2_X1   g0321(.A1(KEYINPUT5), .A2(G41), .ZN(new_n522));
  NOR2_X1   g0322(.A1(KEYINPUT5), .A2(G41), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n485), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n524), .A2(G257), .A3(new_n250), .ZN(new_n525));
  XNOR2_X1  g0325(.A(KEYINPUT5), .B(G41), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n259), .A2(new_n485), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n521), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n347), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n513), .A2(new_n518), .A3(new_n517), .A4(new_n519), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n528), .B1(new_n532), .B2(new_n264), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n344), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT6), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT76), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT76), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT6), .ZN(new_n538));
  NAND2_X1  g0338(.A1(G97), .A2(G107), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n536), .A2(new_n538), .B1(new_n204), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n202), .A2(G107), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n541), .A2(new_n536), .A3(new_n538), .ZN(new_n542));
  OAI21_X1  g0342(.A(G20), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n289), .A2(G77), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n310), .A2(G107), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n330), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n319), .A2(new_n202), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n506), .B2(new_n202), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n531), .B(new_n534), .C1(new_n547), .C2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n506), .A2(new_n441), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n500), .A2(new_n503), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT82), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n500), .A2(new_n492), .A3(new_n503), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n551), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n490), .A2(G200), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n483), .A2(G190), .A3(new_n487), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT78), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n533), .B2(new_n280), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n291), .B1(new_n293), .B2(KEYINPUT73), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n270), .A2(new_n272), .A3(new_n305), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n296), .A2(new_n295), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n544), .B(new_n543), .C1(new_n563), .C2(new_n203), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n549), .B1(new_n564), .B2(new_n301), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n250), .B1(new_n566), .B2(new_n513), .ZN(new_n567));
  OAI211_X1 g0367(.A(KEYINPUT78), .B(G200), .C1(new_n567), .C2(new_n528), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n533), .A2(G190), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n560), .A2(new_n565), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n510), .A2(new_n550), .A3(new_n558), .A4(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT21), .ZN(new_n572));
  INV_X1    g0372(.A(G116), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(new_n206), .B2(G33), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n363), .A2(new_n365), .A3(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n361), .A2(G20), .A3(new_n573), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n300), .A2(new_n223), .B1(G20), .B2(new_n573), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n519), .B(new_n207), .C1(G33), .C2(new_n202), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n578), .A2(KEYINPUT20), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT20), .B1(new_n578), .B2(new_n579), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n577), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n576), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(G303), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n250), .B1(new_n379), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(G257), .A2(G1698), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n407), .A2(G264), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n247), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n524), .A2(G270), .A3(new_n250), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n589), .A2(new_n527), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(G169), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n572), .B1(new_n583), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n264), .B1(new_n485), .B2(new_n526), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n594), .A2(G270), .B1(new_n585), .B2(new_n588), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n595), .A2(G190), .A3(new_n527), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n591), .A2(G200), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n583), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n575), .B(new_n577), .C1(new_n581), .C2(new_n580), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n599), .A2(KEYINPUT21), .A3(G169), .A4(new_n591), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n599), .A2(G179), .A3(new_n527), .A4(new_n595), .ZN(new_n601));
  AND4_X1   g0401(.A1(new_n593), .A2(new_n598), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n527), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n524), .A2(G264), .A3(new_n250), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT85), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n524), .A2(KEYINPUT85), .A3(G264), .A4(new_n250), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n603), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n270), .A2(new_n272), .A3(G257), .A4(G1698), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT84), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n484), .A2(G1698), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n247), .A2(new_n611), .B1(G33), .B2(G294), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n609), .A2(KEYINPUT84), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n264), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n608), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(G169), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n608), .A2(new_n615), .A3(G179), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n270), .A2(new_n272), .A3(new_n207), .A4(G87), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(KEYINPUT22), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT22), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n247), .A2(new_n622), .A3(new_n207), .A4(G87), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT23), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n625), .B1(G20), .B2(new_n203), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n476), .A2(G20), .ZN(new_n628));
  AND2_X1   g0428(.A1(KEYINPUT83), .A2(KEYINPUT24), .ZN(new_n629));
  NOR4_X1   g0429(.A1(new_n626), .A2(new_n627), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(KEYINPUT83), .A2(KEYINPUT24), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n624), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n631), .B1(new_n624), .B2(new_n630), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n301), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT25), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n362), .B2(G107), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n319), .A2(KEYINPUT25), .A3(new_n203), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(new_n506), .B2(new_n203), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n634), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n619), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n616), .A2(G190), .ZN(new_n643));
  AOI21_X1  g0443(.A(G200), .B1(new_n608), .B2(new_n615), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n634), .B(new_n640), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n602), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n471), .A2(new_n571), .A3(new_n646), .ZN(G372));
  AND3_X1   g0447(.A1(new_n339), .A2(KEYINPUT18), .A3(new_n348), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n648), .A2(new_n349), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n397), .A2(new_n464), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n324), .A2(new_n335), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n400), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n650), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n436), .A2(new_n439), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n424), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n491), .A2(new_n507), .A3(new_n488), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n558), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n657), .B1(new_n659), .B2(new_n550), .ZN(new_n660));
  INV_X1    g0460(.A(new_n534), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n533), .A2(G169), .ZN(new_n662));
  NOR3_X1   g0462(.A1(new_n661), .A2(new_n565), .A3(new_n662), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n510), .A2(new_n663), .A3(new_n558), .A4(KEYINPUT26), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n593), .A2(new_n601), .A3(new_n600), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n642), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n558), .A2(new_n658), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n570), .A2(new_n550), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n668), .A2(new_n669), .A3(new_n670), .A4(new_n645), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n665), .A2(new_n658), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n656), .B1(new_n471), .B2(new_n673), .ZN(G369));
  NAND2_X1  g0474(.A1(new_n361), .A2(new_n207), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G213), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n642), .A2(new_n680), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n617), .A2(new_n618), .B1(new_n634), .B2(new_n640), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n680), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT87), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n641), .A2(new_n680), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n642), .A2(new_n645), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n680), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n666), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n681), .B1(new_n687), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n599), .A2(new_n680), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n602), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n667), .B2(new_n692), .ZN(new_n694));
  XOR2_X1   g0494(.A(KEYINPUT86), .B(G330), .Z(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n687), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n691), .A2(new_n698), .ZN(G399));
  INV_X1    g0499(.A(new_n210), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n495), .A2(G116), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G1), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n226), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n704), .B1(new_n705), .B2(new_n702), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  AND4_X1   g0507(.A1(KEYINPUT26), .A2(new_n663), .A3(new_n558), .A4(new_n658), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n510), .A2(new_n663), .A3(new_n558), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n708), .B1(new_n657), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n670), .A2(new_n645), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n558), .B(new_n658), .C1(new_n682), .C2(new_n666), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n658), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OAI211_X1 g0513(.A(KEYINPUT29), .B(new_n688), .C1(new_n710), .C2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n673), .A2(new_n680), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n714), .B1(new_n715), .B2(KEYINPUT29), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n608), .A2(new_n615), .A3(G179), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n483), .A2(new_n487), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n521), .A2(new_n529), .A3(new_n595), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n717), .A2(new_n718), .A3(KEYINPUT30), .A4(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n533), .A2(new_n483), .A3(new_n487), .A4(new_n595), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(new_n618), .ZN(new_n723));
  AOI21_X1  g0523(.A(G179), .B1(new_n595), .B2(new_n527), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n490), .A2(new_n616), .A3(new_n530), .A4(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n720), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n680), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT31), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n726), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT88), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n571), .A2(new_n680), .ZN(new_n733));
  INV_X1    g0533(.A(new_n646), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR4_X1   g0535(.A1(new_n646), .A2(new_n571), .A3(KEYINPUT88), .A4(new_n680), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n731), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n696), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n716), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n707), .B1(new_n739), .B2(G1), .ZN(G364));
  NOR2_X1   g0540(.A1(new_n318), .A2(G20), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n206), .B1(new_n741), .B2(G45), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n702), .A2(KEYINPUT89), .A3(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT89), .ZN(new_n744));
  INV_X1    g0544(.A(new_n742), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n744), .B1(new_n701), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n697), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n749), .B1(new_n696), .B2(new_n694), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n700), .A2(new_n379), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G355), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(G116), .B2(new_n210), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n227), .A2(new_n261), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n700), .A2(new_n247), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n756), .B1(new_n242), .B2(G45), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n753), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G13), .A2(G33), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G20), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n223), .B1(G20), .B2(new_n347), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n748), .B1(new_n758), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n207), .A2(new_n344), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G200), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n767), .A2(KEYINPUT90), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(KEYINPUT90), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n267), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G326), .ZN(new_n773));
  INV_X1    g0573(.A(G294), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n267), .A2(G179), .A3(G200), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n207), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n772), .A2(new_n773), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n777), .A2(KEYINPUT92), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(KEYINPUT92), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n768), .A2(new_n267), .A3(new_n769), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(KEYINPUT33), .B(G317), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n207), .A2(G179), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n784), .A2(G190), .A3(G200), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n784), .A2(new_n267), .A3(G200), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n786), .A2(G303), .B1(new_n788), .B2(G283), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n766), .A2(G190), .A3(new_n280), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n247), .B1(new_n791), .B2(G322), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G190), .A2(G200), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n766), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n784), .A2(new_n793), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G311), .A2(new_n795), .B1(new_n797), .B2(G329), .ZN(new_n798));
  AND3_X1   g0598(.A1(new_n789), .A2(new_n792), .A3(new_n798), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n778), .A2(new_n779), .A3(new_n783), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n788), .A2(G107), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n797), .A2(G159), .ZN(new_n802));
  XNOR2_X1  g0602(.A(KEYINPUT91), .B(KEYINPUT32), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n801), .B1(new_n202), .B2(new_n776), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(new_n441), .B2(new_n785), .ZN(new_n806));
  INV_X1    g0606(.A(G58), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n247), .B1(new_n794), .B2(new_n356), .C1(new_n807), .C2(new_n790), .ZN(new_n808));
  NOR3_X1   g0608(.A1(new_n804), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n809), .B1(new_n413), .B2(new_n772), .C1(new_n298), .C2(new_n780), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n800), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n765), .B1(new_n811), .B2(new_n762), .ZN(new_n812));
  INV_X1    g0612(.A(new_n761), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n812), .B1(new_n694), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n750), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(G396));
  NOR2_X1   g0616(.A1(new_n762), .A2(new_n759), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n748), .B1(G77), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT93), .ZN(new_n820));
  INV_X1    g0620(.A(G283), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n772), .A2(new_n584), .B1(new_n821), .B2(new_n780), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n247), .B1(new_n797), .B2(G311), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n823), .B1(new_n573), .B2(new_n794), .C1(new_n774), .C2(new_n790), .ZN(new_n824));
  INV_X1    g0624(.A(new_n776), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n825), .A2(G97), .B1(new_n788), .B2(G87), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n203), .B2(new_n785), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n822), .A2(new_n824), .A3(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(G132), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n247), .B1(new_n796), .B2(new_n829), .C1(new_n413), .C2(new_n785), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n776), .A2(new_n807), .B1(new_n787), .B2(new_n298), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n791), .A2(G143), .B1(new_n795), .B2(G159), .ZN(new_n832));
  INV_X1    g0632(.A(G137), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n832), .B1(new_n416), .B2(new_n780), .C1(new_n772), .C2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT34), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n830), .B(new_n831), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n834), .A2(new_n835), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n828), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n762), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n464), .A2(new_n680), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n680), .B1(new_n450), .B2(new_n452), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n461), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n840), .B1(new_n842), .B2(new_n464), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n820), .B1(new_n838), .B2(new_n839), .C1(new_n760), .C2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n465), .A2(new_n688), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n673), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n715), .B2(new_n843), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n748), .B1(new_n848), .B2(new_n738), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n848), .A2(new_n738), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n844), .B1(new_n850), .B2(new_n851), .ZN(G384));
  OR2_X1    g0652(.A1(new_n540), .A2(new_n542), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n853), .A2(KEYINPUT35), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(KEYINPUT35), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n854), .A2(G116), .A3(new_n224), .A4(new_n855), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT36), .Z(new_n857));
  OAI211_X1 g0657(.A(new_n226), .B(G77), .C1(new_n807), .C2(new_n298), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n413), .A2(G68), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n206), .B(G13), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  XOR2_X1   g0661(.A(KEYINPUT96), .B(KEYINPUT40), .Z(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n372), .A2(new_n680), .ZN(new_n864));
  AND3_X1   g0664(.A1(new_n397), .A2(new_n400), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n864), .B1(new_n397), .B2(new_n400), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n843), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n737), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT38), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n332), .A2(KEYINPUT16), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n321), .B1(new_n337), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n678), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n350), .A2(KEYINPUT75), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n339), .A2(new_n348), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT18), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n875), .A2(new_n353), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n874), .B1(new_n879), .B2(new_n652), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT37), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n334), .A2(new_n287), .B1(new_n872), .B2(new_n873), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n872), .A2(new_n348), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n339), .A2(new_n873), .ZN(new_n885));
  AND4_X1   g0685(.A1(new_n881), .A2(new_n876), .A3(new_n885), .A4(new_n322), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n870), .B1(new_n880), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n874), .A2(new_n322), .ZN(new_n889));
  INV_X1    g0689(.A(new_n883), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT37), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n876), .A2(new_n885), .A3(new_n881), .A4(new_n322), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(KEYINPUT38), .B(new_n893), .C1(new_n354), .C2(new_n874), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n888), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n863), .B1(new_n869), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT97), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n670), .A2(new_n558), .A3(new_n510), .A4(new_n688), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT88), .B1(new_n898), .B2(new_n646), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n733), .A2(new_n732), .A3(new_n734), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n867), .B1(new_n901), .B2(new_n731), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n888), .A2(new_n894), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT97), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n904), .A2(new_n905), .A3(new_n863), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n897), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT40), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n876), .A2(new_n885), .A3(new_n322), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT37), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(KEYINPUT95), .A3(new_n892), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n324), .B(new_n335), .C1(new_n648), .C2(new_n349), .ZN(new_n912));
  INV_X1    g0712(.A(new_n885), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT95), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n909), .A2(new_n915), .A3(KEYINPUT37), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n911), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n870), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n908), .B1(new_n918), .B2(new_n894), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n902), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n907), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n470), .A2(new_n737), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n695), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n921), .B2(new_n922), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT39), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n892), .A2(KEYINPUT95), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n926), .A2(new_n910), .B1(new_n913), .B2(new_n912), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT38), .B1(new_n927), .B2(new_n916), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n880), .A2(new_n887), .A3(new_n870), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n925), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n888), .A2(new_n894), .A3(KEYINPUT39), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n397), .A2(new_n680), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT94), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n840), .B(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n845), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n936), .B1(new_n672), .B2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n865), .A2(new_n866), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n939), .A2(new_n903), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n650), .B2(new_n873), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n934), .A2(new_n943), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n470), .B(new_n714), .C1(new_n715), .C2(KEYINPUT29), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n656), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n944), .B(new_n946), .Z(new_n947));
  OR2_X1    g0747(.A1(new_n924), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(G1), .B1(new_n318), .B2(G20), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n948), .A2(KEYINPUT98), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n924), .A2(new_n947), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(KEYINPUT98), .B1(new_n948), .B2(new_n949), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n861), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT99), .Z(G367));
  OAI21_X1  g0755(.A(new_n670), .B1(new_n565), .B2(new_n688), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n956), .A2(new_n642), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n680), .B1(new_n957), .B2(new_n550), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n687), .A2(new_n690), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n663), .A2(new_n680), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n956), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n963), .A2(KEYINPUT42), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(KEYINPUT42), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n958), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n698), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT102), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n967), .A2(new_n968), .A3(new_n961), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n555), .A2(new_n688), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n970), .A2(new_n491), .A3(new_n507), .A4(new_n488), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n659), .B2(new_n970), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n973), .A2(KEYINPUT101), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(KEYINPUT102), .B1(new_n698), .B2(new_n962), .ZN(new_n976));
  AND3_X1   g0776(.A1(new_n969), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n975), .B1(new_n969), .B2(new_n976), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT100), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n973), .A2(KEYINPUT101), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OR4_X1    g0782(.A1(new_n966), .A2(new_n977), .A3(new_n978), .A4(new_n982), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n966), .A2(new_n982), .B1(new_n977), .B2(new_n978), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n701), .B(KEYINPUT41), .Z(new_n985));
  INV_X1    g0785(.A(KEYINPUT45), .ZN(new_n986));
  INV_X1    g0786(.A(new_n681), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n959), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n986), .B1(new_n988), .B2(new_n962), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n691), .A2(KEYINPUT45), .A3(new_n961), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n988), .A2(KEYINPUT44), .A3(new_n962), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT44), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n691), .B2(new_n961), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n991), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n967), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n684), .A2(new_n686), .A3(new_n689), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n959), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(new_n697), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n991), .A2(new_n698), .A3(new_n995), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n997), .A2(new_n739), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n985), .B1(new_n1002), .B2(new_n739), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n983), .B(new_n984), .C1(new_n1003), .C2(new_n745), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n763), .B1(new_n210), .B2(new_n445), .C1(new_n756), .C2(new_n235), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n748), .A2(new_n1005), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(G143), .A2(new_n771), .B1(new_n781), .B2(G159), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n794), .A2(new_n413), .B1(new_n796), .B2(new_n833), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n379), .B(new_n1008), .C1(G150), .C2(new_n791), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n785), .A2(new_n807), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n787), .A2(new_n356), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n1010), .B(new_n1011), .C1(G68), .C2(new_n825), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1007), .A2(new_n1009), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n786), .A2(G116), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT46), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(KEYINPUT103), .B(G317), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n247), .B1(new_n797), .B2(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n791), .A2(G303), .B1(new_n795), .B2(G283), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n825), .A2(G107), .B1(new_n788), .B2(G97), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1015), .A2(new_n1017), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n771), .A2(G311), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n774), .B2(new_n780), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1013), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT47), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1006), .B1(new_n1024), .B2(new_n762), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n972), .A2(new_n813), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1004), .A2(new_n1027), .ZN(G387));
  INV_X1    g0828(.A(new_n703), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n751), .A2(new_n1029), .B1(new_n203), .B2(new_n700), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n232), .A2(new_n261), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n316), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n413), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT50), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n703), .B(new_n261), .C1(new_n298), .C2(new_n356), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n755), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1030), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n747), .B1(new_n1037), .B2(new_n763), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n687), .B2(new_n813), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n780), .A2(new_n316), .B1(new_n298), .B2(new_n794), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT105), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n379), .B1(new_n797), .B2(G150), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n356), .B2(new_n785), .C1(new_n202), .C2(new_n787), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT104), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n790), .A2(new_n413), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n776), .A2(new_n445), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1045), .B(new_n1046), .C1(new_n771), .C2(G159), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1041), .A2(new_n1044), .A3(new_n1047), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n776), .A2(new_n821), .B1(new_n785), .B2(new_n774), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1049), .A2(KEYINPUT106), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(KEYINPUT106), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n781), .A2(G311), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n791), .A2(new_n1016), .B1(new_n795), .B2(G303), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(KEYINPUT107), .B(G322), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1052), .B(new_n1053), .C1(new_n772), .C2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT48), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1050), .B(new_n1051), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT108), .Z(new_n1058));
  NAND2_X1  g0858(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1058), .A2(KEYINPUT49), .A3(new_n1059), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n379), .B1(new_n796), .B2(new_n773), .C1(new_n573), .C2(new_n787), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT109), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(KEYINPUT49), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1048), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1039), .B1(new_n1065), .B2(new_n762), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n1000), .B2(new_n745), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n739), .A2(new_n1000), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n701), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n739), .A2(new_n1000), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1067), .B1(new_n1069), .B2(new_n1070), .ZN(G393));
  INV_X1    g0871(.A(new_n1001), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n698), .B1(new_n991), .B2(new_n995), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1068), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1074), .A2(new_n1002), .A3(new_n701), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n755), .A2(new_n239), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1076), .B(new_n763), .C1(new_n202), .C2(new_n210), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n771), .A2(G150), .B1(G159), .B2(new_n791), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT51), .Z(new_n1079));
  AOI22_X1  g0879(.A1(new_n786), .A2(G68), .B1(new_n797), .B2(G143), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT110), .Z(new_n1081));
  NOR2_X1   g0881(.A1(new_n780), .A2(new_n413), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n776), .A2(new_n356), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n247), .B1(new_n794), .B2(new_n316), .C1(new_n441), .C2(new_n787), .ZN(new_n1084));
  NOR4_X1   g0884(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n771), .A2(G317), .B1(G311), .B2(new_n791), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT52), .Z(new_n1087));
  OAI221_X1 g0887(.A(new_n379), .B1(new_n796), .B2(new_n1054), .C1(new_n774), .C2(new_n794), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n801), .B1(new_n821), .B2(new_n785), .C1(new_n573), .C2(new_n776), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n1088), .B(new_n1089), .C1(G303), .C2(new_n781), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n1079), .A2(new_n1085), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n748), .B(new_n1077), .C1(new_n1091), .C2(new_n839), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT111), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n761), .B2(new_n962), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1094), .B1(new_n1095), .B2(new_n745), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1075), .A2(new_n1096), .ZN(G390));
  OAI21_X1  g0897(.A(new_n933), .B1(new_n938), .B2(new_n940), .ZN(new_n1098));
  AOI21_X1  g0898(.A(KEYINPUT39), .B1(new_n918), .B2(new_n894), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n888), .A2(new_n894), .A3(KEYINPUT39), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n688), .B(new_n843), .C1(new_n710), .C2(new_n713), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n936), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n941), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n933), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n918), .B2(new_n894), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n737), .A2(new_n696), .A3(new_n843), .A4(new_n941), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1101), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n932), .A2(new_n1098), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n737), .A2(new_n868), .A3(G330), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n745), .B(new_n1110), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT116), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n760), .B1(new_n930), .B2(new_n931), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n771), .A2(G128), .B1(G132), .B2(new_n791), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT113), .ZN(new_n1117));
  INV_X1    g0917(.A(G125), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT54), .B(G143), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n247), .B1(new_n796), .B2(new_n1118), .C1(new_n794), .C2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(G159), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n776), .A2(new_n1121), .B1(new_n787), .B2(new_n413), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n785), .A2(new_n416), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT53), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1123), .B(new_n1125), .C1(new_n833), .C2(new_n780), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n379), .B1(new_n794), .B2(new_n202), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(G294), .B2(new_n797), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n786), .A2(G87), .B1(new_n788), .B2(G68), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1128), .B(new_n1129), .C1(new_n772), .C2(new_n821), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n776), .A2(new_n356), .B1(new_n790), .B2(new_n573), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n781), .A2(G107), .B1(KEYINPUT114), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(KEYINPUT114), .B2(new_n1131), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n1117), .A2(new_n1126), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n762), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n747), .B1(new_n316), .B2(new_n817), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(KEYINPUT115), .B1(new_n1115), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n759), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT115), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1139), .A2(new_n1140), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n1113), .A2(new_n1114), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1114), .B1(new_n1113), .B2(new_n1142), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT112), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1110), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1104), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n729), .A2(new_n730), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n899), .B2(new_n900), .ZN(new_n1150));
  INV_X1    g0950(.A(G330), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n843), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1148), .B(new_n1109), .C1(new_n1153), .C2(new_n941), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n737), .A2(new_n696), .A3(new_n843), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n1155), .A2(new_n940), .B1(new_n1156), .B2(new_n868), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1154), .B1(new_n1157), .B2(new_n938), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n470), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n945), .A2(new_n656), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1147), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1101), .A2(new_n1108), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1112), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1166), .A2(new_n1158), .A3(new_n1110), .A4(new_n1161), .ZN(new_n1167));
  AND4_X1   g0967(.A1(new_n1146), .A2(new_n1163), .A3(new_n701), .A4(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n702), .B1(new_n1147), .B2(new_n1162), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1146), .B1(new_n1169), .B2(new_n1167), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1145), .B1(new_n1168), .B2(new_n1170), .ZN(G378));
  INV_X1    g0971(.A(KEYINPUT57), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n1167), .B2(new_n1161), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1151), .B1(new_n919), .B2(new_n902), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n905), .B1(new_n904), .B2(new_n863), .ZN(new_n1175));
  AOI211_X1 g0975(.A(KEYINPUT97), .B(new_n862), .C1(new_n902), .C2(new_n903), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1174), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT119), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n440), .B(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n422), .A2(new_n873), .ZN(new_n1181));
  XOR2_X1   g0981(.A(new_n1181), .B(KEYINPUT118), .Z(new_n1182));
  XNOR2_X1  g0982(.A(new_n1180), .B(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1177), .A2(new_n1184), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1174), .B(new_n1183), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1185), .A2(new_n944), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n944), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1173), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n701), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n944), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1183), .B1(new_n907), .B2(new_n1174), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1186), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1192), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n1187), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1167), .A2(new_n1161), .ZN(new_n1197));
  AOI21_X1  g0997(.A(KEYINPUT57), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1191), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1184), .A2(new_n759), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n748), .B1(G50), .B2(new_n818), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(G33), .A2(G41), .ZN(new_n1202));
  AOI211_X1 g1002(.A(G50), .B(new_n1202), .C1(new_n379), .C2(new_n260), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n787), .A2(new_n807), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1205), .B1(new_n356), .B2(new_n785), .C1(new_n298), .C2(new_n776), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n260), .B(new_n379), .C1(new_n790), .C2(new_n203), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n445), .A2(new_n794), .B1(new_n796), .B2(new_n821), .ZN(new_n1208));
  NOR3_X1   g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n202), .B2(new_n780), .C1(new_n573), .C2(new_n772), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT58), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1203), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n785), .A2(new_n1119), .ZN(new_n1213));
  INV_X1    g1013(.A(G128), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n790), .A2(new_n1214), .B1(new_n794), .B2(new_n833), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1213), .B(new_n1215), .C1(G150), .C2(new_n825), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1216), .B1(new_n829), .B2(new_n780), .C1(new_n772), .C2(new_n1118), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(KEYINPUT59), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1202), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(KEYINPUT117), .B(G124), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1219), .B1(new_n797), .B2(new_n1220), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1218), .B(new_n1221), .C1(new_n1121), .C2(new_n787), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1217), .A2(KEYINPUT59), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1212), .B1(new_n1211), .B2(new_n1210), .C1(new_n1222), .C2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1201), .B1(new_n1224), .B2(new_n762), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1196), .A2(new_n745), .B1(new_n1200), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1199), .A2(new_n1226), .ZN(G375));
  INV_X1    g1027(.A(new_n985), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1150), .A2(new_n695), .A3(new_n1152), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1112), .B1(new_n1229), .B2(new_n941), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(new_n939), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1231), .A2(new_n1160), .A3(new_n1154), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1162), .A2(new_n1228), .A3(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n940), .A2(new_n759), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n748), .B1(G68), .B2(new_n818), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(G294), .A2(new_n771), .B1(new_n781), .B2(G116), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n794), .A2(new_n203), .B1(new_n796), .B2(new_n584), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n247), .B(new_n1237), .C1(G283), .C2(new_n791), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n1011), .B(new_n1046), .C1(G97), .C2(new_n786), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1236), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n247), .B1(new_n796), .B2(new_n1214), .C1(new_n416), .C2(new_n794), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1205), .B1(new_n413), .B2(new_n776), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(G159), .C2(new_n786), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1243), .B(KEYINPUT120), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n771), .A2(G132), .B1(G137), .B2(new_n791), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1245), .B1(new_n780), .B2(new_n1119), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1240), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT121), .ZN(new_n1248));
  OR2_X1    g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n839), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1235), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1158), .A2(new_n745), .B1(new_n1234), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1233), .A2(new_n1252), .ZN(G381));
  OR2_X1    g1053(.A1(G393), .A2(G396), .ZN(new_n1254));
  OR4_X1    g1054(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1169), .A2(new_n1167), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1256), .A2(new_n1142), .A3(new_n1113), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  OR4_X1    g1058(.A1(G375), .A2(new_n1255), .A3(G381), .A4(new_n1258), .ZN(G407));
  INV_X1    g1059(.A(G375), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n679), .A2(G213), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1260), .A2(new_n1257), .A3(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(G407), .A2(G213), .A3(new_n1263), .ZN(G409));
  INV_X1    g1064(.A(KEYINPUT126), .ZN(new_n1265));
  OAI211_X1 g1065(.A(G378), .B(new_n1226), .C1(new_n1191), .C2(new_n1198), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1228), .B(new_n1197), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n745), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1200), .A2(new_n1225), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1267), .A2(new_n1268), .A3(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1257), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1262), .B1(new_n1266), .B2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1104), .B1(new_n1229), .B2(new_n941), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n737), .A2(G330), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n940), .B1(new_n1274), .B2(new_n1152), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n939), .A2(new_n1230), .B1(new_n1273), .B2(new_n1275), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1276), .A2(KEYINPUT122), .A3(KEYINPUT60), .A4(new_n1160), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1231), .A2(KEYINPUT60), .A3(new_n1160), .A4(new_n1154), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT122), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT60), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1232), .A2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n702), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1277), .A2(new_n1280), .A3(new_n1282), .A4(new_n1283), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n1284), .A2(G384), .A3(new_n1252), .ZN(new_n1285));
  AOI21_X1  g1085(.A(G384), .B1(new_n1284), .B2(new_n1252), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1272), .A2(KEYINPUT63), .A3(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(KEYINPUT63), .B1(new_n1272), .B2(new_n1287), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(G393), .B(new_n815), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1004), .A2(new_n1027), .A3(G390), .ZN(new_n1292));
  AOI21_X1  g1092(.A(G390), .B1(new_n1004), .B2(new_n1027), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1291), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT61), .ZN(new_n1295));
  INV_X1    g1095(.A(G390), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n983), .A2(new_n984), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1002), .A2(new_n739), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1228), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1297), .B1(new_n1299), .B2(new_n742), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1027), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1296), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1004), .A2(new_n1027), .A3(G390), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1302), .A2(new_n1290), .A3(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1294), .A2(new_n1295), .A3(new_n1304), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(new_n1288), .A2(new_n1289), .A3(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(G2897), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1261), .A2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1308), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1284), .A2(new_n1252), .ZN(new_n1310));
  INV_X1    g1110(.A(G384), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1284), .A2(G384), .A3(new_n1252), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT123), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1261), .B1(new_n1314), .B2(new_n1307), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(new_n1314), .B2(new_n1307), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1312), .A2(new_n1313), .A3(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT124), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1309), .A2(new_n1317), .A3(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1318), .B1(new_n1309), .B2(new_n1317), .ZN(new_n1320));
  OAI21_X1  g1120(.A(KEYINPUT125), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1316), .ZN(new_n1322));
  NOR3_X1   g1122(.A1(new_n1285), .A2(new_n1286), .A3(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1308), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1324), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1325));
  OAI21_X1  g1125(.A(KEYINPUT124), .B1(new_n1323), .B2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT125), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1309), .A2(new_n1317), .A3(new_n1318), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1326), .A2(new_n1327), .A3(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1266), .A2(new_n1271), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1261), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1321), .A2(new_n1329), .A3(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1265), .B1(new_n1306), .B2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT63), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1330), .A2(new_n1261), .A3(new_n1287), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1305), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1272), .A2(KEYINPUT63), .A3(new_n1287), .ZN(new_n1337));
  AND4_X1   g1137(.A1(new_n1265), .A2(new_n1336), .A3(new_n1332), .A4(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1326), .A2(new_n1328), .ZN(new_n1339));
  AOI21_X1  g1139(.A(KEYINPUT61), .B1(new_n1339), .B2(new_n1331), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1335), .A2(KEYINPUT62), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT62), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1272), .A2(new_n1342), .A3(new_n1287), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1340), .A2(KEYINPUT127), .A3(new_n1341), .A4(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1294), .A2(new_n1304), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  AND4_X1   g1146(.A1(new_n1342), .A2(new_n1330), .A3(new_n1261), .A4(new_n1287), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1342), .B1(new_n1272), .B2(new_n1287), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(KEYINPUT127), .B1(new_n1349), .B2(new_n1340), .ZN(new_n1350));
  OAI22_X1  g1150(.A1(new_n1333), .A2(new_n1338), .B1(new_n1346), .B2(new_n1350), .ZN(G405));
  NAND2_X1  g1151(.A1(G375), .A2(new_n1257), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1352), .A2(new_n1266), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1353), .A2(new_n1287), .ZN(new_n1354));
  OAI211_X1 g1154(.A(new_n1352), .B(new_n1266), .C1(new_n1286), .C2(new_n1285), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1354), .A2(new_n1355), .ZN(new_n1356));
  XNOR2_X1  g1156(.A(new_n1356), .B(new_n1345), .ZN(G402));
endmodule


