//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 1 0 0 0 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1325, new_n1326, new_n1327,
    new_n1328, new_n1329, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1389,
    new_n1390, new_n1391, new_n1392, new_n1393;
  OR2_X1    g0000(.A1(KEYINPUT64), .A2(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(KEYINPUT64), .A2(G50), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n208));
  INV_X1    g0008(.A(G68), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n208), .B1(new_n209), .B2(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n207), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT66), .ZN(new_n218));
  INV_X1    g0018(.A(KEYINPUT1), .ZN(new_n219));
  OR2_X1    g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n219), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n207), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT0), .Z(new_n224));
  AND2_X1   g0024(.A1(KEYINPUT65), .A2(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(KEYINPUT65), .A2(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(G58), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(new_n209), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n224), .B1(new_n229), .B2(new_n233), .ZN(new_n234));
  AND3_X1   g0034(.A1(new_n220), .A2(new_n221), .A3(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XOR2_X1   g0045(.A(G50), .B(G58), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  INV_X1    g0051(.A(KEYINPUT16), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT7), .ZN(new_n253));
  AND2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n253), .B1(new_n227), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT3), .B(G33), .ZN(new_n258));
  INV_X1    g0058(.A(G20), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n253), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n257), .A2(new_n209), .A3(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT75), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G58), .A2(G68), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n259), .B1(new_n231), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G159), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n263), .B1(new_n265), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n264), .ZN(new_n271));
  OAI21_X1  g0071(.A(G20), .B1(new_n271), .B2(new_n202), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G20), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G159), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n272), .A2(KEYINPUT75), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n252), .B1(new_n262), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT76), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n228), .ZN(new_n281));
  OR2_X1    g0081(.A1(KEYINPUT65), .A2(G20), .ZN(new_n282));
  NAND2_X1  g0082(.A1(KEYINPUT65), .A2(G20), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n253), .B1(new_n284), .B2(new_n258), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT74), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n256), .A2(new_n286), .A3(KEYINPUT7), .A4(new_n259), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n259), .A2(KEYINPUT7), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT74), .B1(new_n258), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n285), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G68), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n265), .A2(new_n269), .A3(new_n263), .ZN(new_n292));
  AOI21_X1  g0092(.A(KEYINPUT75), .B1(new_n272), .B2(new_n274), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n291), .A2(KEYINPUT16), .A3(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(KEYINPUT7), .B1(new_n284), .B2(new_n258), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n256), .A2(new_n253), .A3(new_n259), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(G68), .A3(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n298), .A2(new_n270), .A3(new_n275), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n299), .A2(KEYINPUT76), .A3(new_n252), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n279), .A2(new_n281), .A3(new_n295), .A4(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(KEYINPUT69), .A2(G58), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n302), .B(KEYINPUT8), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  OR2_X1    g0104(.A1(KEYINPUT67), .A2(G1), .ZN(new_n305));
  NAND2_X1  g0105(.A1(KEYINPUT67), .A2(G1), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n305), .A2(G13), .A3(G20), .A4(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  AND2_X1   g0108(.A1(KEYINPUT67), .A2(G1), .ZN(new_n309));
  NOR2_X1   g0109(.A1(KEYINPUT67), .A2(G1), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n281), .B1(new_n311), .B2(G20), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n308), .B1(new_n312), .B2(new_n304), .ZN(new_n313));
  INV_X1    g0113(.A(G200), .ZN(new_n314));
  INV_X1    g0114(.A(G274), .ZN(new_n315));
  AND2_X1   g0115(.A1(G1), .A2(G13), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G33), .A2(G41), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G1), .ZN(new_n319));
  NOR2_X1   g0119(.A1(G41), .A2(G45), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n318), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n316), .A2(new_n317), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT67), .B(G1), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(new_n320), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n322), .B1(new_n325), .B2(new_n237), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G223), .ZN(new_n328));
  INV_X1    g0128(.A(G1698), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n258), .B(new_n330), .C1(G226), .C2(new_n329), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G33), .A2(G87), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n323), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n314), .B1(new_n327), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n323), .B1(new_n331), .B2(new_n332), .ZN(new_n337));
  INV_X1    g0137(.A(G190), .ZN(new_n338));
  NOR3_X1   g0138(.A1(new_n337), .A2(new_n326), .A3(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n301), .A2(new_n313), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT17), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n341), .B(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT18), .ZN(new_n344));
  INV_X1    g0144(.A(new_n313), .ZN(new_n345));
  AOI211_X1 g0145(.A(new_n278), .B(KEYINPUT16), .C1(new_n294), .C2(new_n298), .ZN(new_n346));
  AOI21_X1  g0146(.A(KEYINPUT76), .B1(new_n299), .B2(new_n252), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n281), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n276), .B1(new_n290), .B2(G68), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n349), .B1(new_n350), .B2(KEYINPUT16), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n345), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n327), .A2(new_n335), .A3(G179), .ZN(new_n353));
  OAI21_X1  g0153(.A(G169), .B1(new_n337), .B2(new_n326), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n344), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  AOI211_X1 g0157(.A(new_n344), .B(new_n356), .C1(new_n301), .C2(new_n313), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n357), .B1(new_n358), .B2(KEYINPUT77), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n356), .B1(new_n301), .B2(new_n313), .ZN(new_n360));
  NOR3_X1   g0160(.A1(new_n360), .A2(KEYINPUT77), .A3(KEYINPUT18), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n343), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n363), .A2(KEYINPUT78), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n363), .A2(KEYINPUT78), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n258), .A2(G222), .A3(new_n329), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n256), .A2(G77), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n258), .A2(G1698), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n366), .B(new_n367), .C1(new_n368), .C2(new_n328), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n334), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n318), .A2(new_n319), .A3(new_n321), .ZN(new_n371));
  INV_X1    g0171(.A(new_n325), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n371), .B1(new_n372), .B2(G226), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT68), .ZN(new_n374));
  AND3_X1   g0174(.A1(new_n370), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n374), .B1(new_n370), .B2(new_n373), .ZN(new_n376));
  OAI21_X1  g0176(.A(G190), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n370), .A2(new_n373), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT68), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n370), .A2(new_n373), .A3(new_n374), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n379), .A2(G200), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n303), .A2(G33), .A3(new_n227), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n273), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n281), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n307), .A2(G50), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n386), .B1(G50), .B2(new_n312), .ZN(new_n387));
  AND3_X1   g0187(.A1(new_n385), .A2(KEYINPUT9), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT9), .B1(new_n385), .B2(new_n387), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n377), .A2(new_n381), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT10), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT10), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n377), .A2(new_n381), .A3(new_n390), .A4(new_n393), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G179), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n375), .B2(new_n376), .ZN(new_n397));
  INV_X1    g0197(.A(G169), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n379), .A2(new_n398), .A3(new_n380), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n385), .A2(new_n387), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n397), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n258), .A2(G232), .A3(new_n329), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n256), .A2(G107), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n402), .B(new_n403), .C1(new_n368), .C2(new_n210), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n334), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n371), .B1(new_n372), .B2(G244), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G200), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n284), .A2(G77), .ZN(new_n409));
  XNOR2_X1  g0209(.A(KEYINPUT8), .B(G58), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n227), .A2(G33), .ZN(new_n411));
  XNOR2_X1  g0211(.A(KEYINPUT15), .B(G87), .ZN(new_n412));
  OAI221_X1 g0212(.A(new_n409), .B1(new_n267), .B2(new_n410), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n281), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT70), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n307), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n311), .A2(KEYINPUT70), .A3(G13), .A4(G20), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(G77), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n414), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n405), .A2(new_n406), .A3(G190), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n416), .A2(new_n417), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n312), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(new_n419), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n408), .A2(new_n421), .A3(new_n422), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n421), .A2(new_n426), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n405), .A2(new_n406), .A3(new_n396), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n407), .A2(new_n398), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n401), .A2(new_n427), .A3(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n395), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT14), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT13), .ZN(new_n435));
  OAI211_X1 g0235(.A(G238), .B(new_n323), .C1(new_n324), .C2(new_n320), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n322), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT71), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n436), .A2(new_n322), .A3(KEYINPUT71), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n237), .A2(G1698), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(G226), .B2(G1698), .ZN(new_n443));
  INV_X1    g0243(.A(G97), .ZN(new_n444));
  OAI22_X1  g0244(.A1(new_n443), .A2(new_n256), .B1(new_n266), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n334), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n435), .B1(new_n441), .B2(new_n446), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n436), .A2(new_n322), .A3(KEYINPUT71), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT71), .B1(new_n436), .B2(new_n322), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n435), .B(new_n446), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n434), .B(G169), .C1(new_n447), .C2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT73), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(G169), .B1(new_n447), .B2(new_n451), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT14), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT13), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n450), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n459), .A2(KEYINPUT73), .A3(new_n434), .A4(G169), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n458), .A2(G179), .A3(new_n450), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n454), .A2(new_n456), .A3(new_n460), .A4(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n209), .B1(new_n424), .B2(KEYINPUT12), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT72), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT12), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(G68), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n418), .A2(new_n467), .B1(new_n466), .B2(new_n307), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n464), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n468), .ZN(new_n470));
  OAI21_X1  g0270(.A(KEYINPUT72), .B1(new_n470), .B2(new_n463), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n273), .A2(G50), .B1(G20), .B2(new_n209), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(new_n411), .B2(new_n419), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n281), .ZN(new_n474));
  XNOR2_X1  g0274(.A(new_n474), .B(KEYINPUT11), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n469), .A2(new_n471), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n462), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n459), .A2(new_n338), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n314), .B1(new_n458), .B2(new_n450), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n476), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n433), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  NOR3_X1   g0282(.A1(new_n364), .A2(new_n365), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT86), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n266), .A2(G97), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G283), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n484), .B1(new_n284), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n227), .A2(KEYINPUT86), .A3(new_n485), .A4(new_n486), .ZN(new_n489));
  INV_X1    g0289(.A(G116), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n280), .A2(new_n228), .B1(G20), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  XOR2_X1   g0292(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n311), .A2(G33), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n281), .A2(new_n490), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n423), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n416), .A2(new_n417), .A3(new_n490), .ZN(new_n498));
  NOR2_X1   g0298(.A1(KEYINPUT87), .A2(KEYINPUT20), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n488), .A2(new_n489), .A3(new_n499), .A4(new_n491), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n494), .A2(new_n497), .A3(new_n498), .A4(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n329), .A2(G264), .ZN(new_n502));
  NOR2_X1   g0302(.A1(G257), .A2(G1698), .ZN(new_n503));
  OAI22_X1  g0303(.A1(new_n502), .A2(new_n503), .B1(new_n254), .B2(new_n255), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n504), .B(new_n334), .C1(G303), .C2(new_n258), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n305), .A2(G45), .A3(new_n306), .ZN(new_n506));
  AND2_X1   g0306(.A1(KEYINPUT5), .A2(G41), .ZN(new_n507));
  NOR2_X1   g0307(.A1(KEYINPUT5), .A2(G41), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g0309(.A(G270), .B(new_n323), .C1(new_n506), .C2(new_n509), .ZN(new_n510));
  XNOR2_X1  g0310(.A(KEYINPUT5), .B(G41), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n318), .A2(new_n311), .A3(new_n511), .A4(G45), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n505), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n513), .A2(G169), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n501), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT21), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT89), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n515), .A2(KEYINPUT89), .A3(new_n516), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n501), .A2(new_n514), .A3(KEYINPUT21), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n505), .A2(G179), .A3(new_n510), .A4(new_n512), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n501), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT88), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT88), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n501), .A2(new_n527), .A3(new_n524), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n522), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n521), .A2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n513), .A2(G200), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n338), .B2(new_n513), .ZN(new_n533));
  OR2_X1    g0333(.A1(new_n533), .A2(new_n501), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT79), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT6), .ZN(new_n536));
  AND2_X1   g0336(.A1(G97), .A2(G107), .ZN(new_n537));
  NOR2_X1   g0337(.A1(G97), .A2(G107), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(G107), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n540), .A2(KEYINPUT6), .A3(G97), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n227), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n267), .A2(new_n419), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n535), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n543), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n540), .A2(KEYINPUT6), .A3(G97), .ZN(new_n546));
  XNOR2_X1  g0346(.A(G97), .B(G107), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n546), .B1(new_n547), .B2(new_n536), .ZN(new_n548));
  OAI211_X1 g0348(.A(KEYINPUT79), .B(new_n545), .C1(new_n548), .C2(new_n227), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n296), .A2(G107), .A3(new_n297), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n544), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n281), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n307), .A2(G97), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n495), .A2(new_n349), .A3(new_n307), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n553), .B1(new_n555), .B2(G97), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(G244), .B(new_n329), .C1(new_n254), .C2(new_n255), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT4), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n258), .A2(KEYINPUT4), .A3(G244), .A4(new_n329), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n258), .A2(G250), .A3(G1698), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n560), .A2(new_n561), .A3(new_n486), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n334), .ZN(new_n564));
  OAI211_X1 g0364(.A(G257), .B(new_n323), .C1(new_n506), .C2(new_n509), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n512), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT80), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT80), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n565), .A2(new_n568), .A3(new_n512), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n564), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n398), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n334), .A2(new_n563), .B1(new_n566), .B2(KEYINPUT80), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n572), .A2(new_n396), .A3(new_n569), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n557), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(KEYINPUT81), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT81), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n557), .A2(new_n571), .A3(new_n573), .A4(new_n576), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n564), .A2(new_n567), .A3(new_n569), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G190), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n570), .A2(G200), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n579), .A2(new_n552), .A3(new_n556), .A4(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n575), .A2(new_n577), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n227), .A2(new_n258), .A3(G87), .ZN(new_n583));
  NOR2_X1   g0383(.A1(KEYINPUT90), .A2(KEYINPUT22), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(KEYINPUT23), .A2(G107), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n586), .B1(new_n587), .B2(G20), .ZN(new_n588));
  NOR2_X1   g0388(.A1(KEYINPUT23), .A2(G107), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n588), .B1(new_n284), .B2(new_n589), .ZN(new_n590));
  XOR2_X1   g0390(.A(KEYINPUT90), .B(KEYINPUT22), .Z(new_n591));
  NAND4_X1  g0391(.A1(new_n591), .A2(G87), .A3(new_n227), .A4(new_n258), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n585), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT24), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT24), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n585), .A2(new_n590), .A3(new_n595), .A4(new_n592), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n349), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n307), .A2(G107), .ZN(new_n598));
  XNOR2_X1  g0398(.A(new_n598), .B(KEYINPUT25), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n540), .B2(new_n554), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(G250), .B(new_n329), .C1(new_n254), .C2(new_n255), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT92), .ZN(new_n603));
  OR2_X1    g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n602), .A2(new_n603), .B1(G33), .B2(G294), .ZN(new_n605));
  OAI211_X1 g0405(.A(G257), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT91), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n604), .B(new_n605), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n334), .ZN(new_n611));
  INV_X1    g0411(.A(new_n506), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n334), .B1(new_n612), .B2(new_n511), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(G264), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n611), .A2(new_n512), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G200), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n610), .A2(new_n334), .B1(G264), .B2(new_n613), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n617), .A2(G190), .A3(new_n512), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n601), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n282), .A2(G33), .A3(G97), .A4(new_n283), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT19), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g0422(.A(new_n622), .B(KEYINPUT85), .ZN(new_n623));
  NAND3_X1  g0423(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n282), .A2(new_n283), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT84), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n538), .A2(new_n211), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n284), .A2(new_n256), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n625), .A2(new_n627), .ZN(new_n630));
  AOI22_X1  g0430(.A1(G68), .A2(new_n629), .B1(new_n630), .B2(KEYINPUT84), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n623), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n632), .A2(new_n281), .B1(new_n418), .B2(new_n412), .ZN(new_n633));
  OAI211_X1 g0433(.A(G244), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n634));
  OAI211_X1 g0434(.A(G238), .B(new_n329), .C1(new_n254), .C2(new_n255), .ZN(new_n635));
  NAND2_X1  g0435(.A1(G33), .A2(G116), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT83), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n634), .A2(new_n635), .A3(KEYINPUT83), .A4(new_n636), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n323), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n212), .B1(new_n316), .B2(new_n317), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n506), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(KEYINPUT82), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT82), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n506), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n612), .A2(new_n318), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n641), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(G190), .ZN(new_n651));
  OAI21_X1  g0451(.A(G200), .B1(new_n641), .B2(new_n649), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n555), .A2(G87), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n633), .A2(new_n651), .A3(new_n652), .A4(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT85), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n622), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n629), .A2(G68), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n630), .A2(KEYINPUT84), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(new_n658), .A3(new_n628), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n281), .B1(new_n656), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n418), .A2(new_n412), .ZN(new_n661));
  INV_X1    g0461(.A(new_n412), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n555), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n660), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n650), .A2(new_n396), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n398), .B1(new_n641), .B2(new_n649), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n619), .A2(new_n654), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n601), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n617), .A2(new_n396), .A3(new_n512), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n615), .A2(new_n398), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n582), .A2(new_n668), .A3(new_n672), .ZN(new_n673));
  AND4_X1   g0473(.A1(new_n483), .A2(new_n531), .A3(new_n534), .A4(new_n673), .ZN(G372));
  AOI211_X1 g0474(.A(new_n480), .B(new_n343), .C1(new_n477), .C2(new_n431), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n360), .A2(KEYINPUT18), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(new_n358), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n392), .A2(KEYINPUT94), .A3(new_n394), .ZN(new_n678));
  AOI21_X1  g0478(.A(KEYINPUT94), .B1(new_n392), .B2(new_n394), .ZN(new_n679));
  OAI22_X1  g0479(.A1(new_n675), .A2(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n401), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n667), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n582), .A2(new_n668), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n521), .A2(new_n685), .A3(new_n529), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n683), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT93), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n574), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n557), .A2(new_n571), .A3(new_n573), .A4(KEYINPUT93), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n689), .A2(new_n667), .A3(new_n654), .A4(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT26), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n654), .A2(new_n667), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n575), .A2(new_n577), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(new_n695), .A3(KEYINPUT26), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n687), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n483), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n682), .A2(new_n699), .ZN(G369));
  NAND2_X1  g0500(.A1(new_n227), .A2(G13), .ZN(new_n701));
  OR3_X1    g0501(.A1(new_n701), .A2(KEYINPUT27), .A3(new_n324), .ZN(new_n702));
  OAI21_X1  g0502(.A(KEYINPUT27), .B1(new_n701), .B2(new_n324), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G213), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(G343), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n530), .A2(new_n501), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT95), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n501), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n521), .A2(new_n529), .A3(new_n534), .A4(new_n709), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n707), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n708), .B1(new_n707), .B2(new_n710), .ZN(new_n712));
  OAI21_X1  g0512(.A(G330), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n601), .B1(new_n398), .B2(new_n615), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n706), .B1(new_n597), .B2(new_n600), .ZN(new_n716));
  AOI22_X1  g0516(.A1(new_n715), .A2(new_n670), .B1(new_n619), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n685), .A2(new_n706), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT96), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n706), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n672), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT96), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n619), .A2(new_n716), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n685), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n721), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n719), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n714), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n706), .B1(new_n521), .B2(new_n529), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n719), .A2(new_n725), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(KEYINPUT97), .B1(new_n730), .B2(new_n721), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(KEYINPUT97), .A3(new_n721), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n728), .B1(new_n731), .B2(new_n733), .ZN(G399));
  INV_X1    g0534(.A(new_n222), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G41), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n319), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n627), .A2(G116), .ZN(new_n738));
  AOI22_X1  g0538(.A1(new_n737), .A2(new_n738), .B1(new_n233), .B2(new_n736), .ZN(new_n739));
  XOR2_X1   g0539(.A(new_n739), .B(KEYINPUT28), .Z(new_n740));
  NAND2_X1  g0540(.A1(new_n698), .A2(new_n720), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT99), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT29), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n706), .B1(new_n687), .B2(new_n697), .ZN(new_n745));
  OAI21_X1  g0545(.A(KEYINPUT99), .B1(new_n745), .B2(KEYINPUT29), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n684), .A2(new_n686), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n667), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n691), .A2(new_n692), .ZN(new_n750));
  AOI21_X1  g0550(.A(KEYINPUT26), .B1(new_n694), .B2(new_n695), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  OAI211_X1 g0552(.A(KEYINPUT29), .B(new_n720), .C1(new_n749), .C2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(KEYINPUT100), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n750), .A2(new_n751), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n687), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT100), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n756), .A2(new_n757), .A3(KEYINPUT29), .A4(new_n720), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n747), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G330), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT30), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n572), .A2(new_n611), .A3(new_n569), .A4(new_n614), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n639), .A2(new_n640), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(new_n334), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n644), .A2(new_n646), .B1(new_n318), .B2(new_n612), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n765), .A2(new_n524), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n762), .B1(new_n763), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n513), .A2(new_n396), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n769), .B1(new_n572), .B2(new_n569), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n765), .A2(KEYINPUT98), .A3(new_n766), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT98), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(new_n641), .B2(new_n649), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n770), .A2(new_n615), .A3(new_n771), .A4(new_n773), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n641), .A2(new_n649), .A3(new_n523), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n775), .A2(new_n617), .A3(KEYINPUT30), .A4(new_n578), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n768), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(new_n706), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT31), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AND4_X1   g0580(.A1(new_n521), .A2(new_n529), .A3(new_n534), .A4(new_n720), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n780), .B1(new_n673), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n778), .A2(new_n779), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n761), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n760), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n740), .B1(new_n787), .B2(G1), .ZN(G364));
  OR2_X1    g0588(.A1(new_n711), .A2(new_n712), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n761), .ZN(new_n791));
  INV_X1    g0591(.A(new_n701), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G45), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(new_n737), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n791), .A2(new_n713), .A3(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n794), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n258), .A2(new_n222), .ZN(new_n797));
  INV_X1    g0597(.A(G355), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n797), .A2(new_n798), .B1(G116), .B2(new_n222), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n256), .A2(new_n222), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT101), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G45), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n802), .B1(new_n803), .B2(new_n233), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n247), .A2(G45), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n799), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(G13), .A2(G33), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(G20), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n228), .B1(G20), .B2(new_n398), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n796), .B1(new_n806), .B2(new_n812), .ZN(new_n813));
  NOR4_X1   g0613(.A1(new_n227), .A2(G179), .A3(G190), .A4(new_n314), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n815), .A2(KEYINPUT103), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(KEYINPUT103), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(new_n540), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n227), .A2(new_n396), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(G200), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n338), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n819), .B1(G50), .B2(new_n822), .ZN(new_n823));
  NOR4_X1   g0623(.A1(new_n259), .A2(new_n338), .A3(new_n314), .A4(G179), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n825), .A2(KEYINPUT102), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(KEYINPUT102), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(new_n211), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n338), .A2(G200), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n820), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(G190), .A2(G200), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n820), .A2(new_n832), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n230), .A2(new_n831), .B1(new_n833), .B2(new_n419), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n829), .A2(new_n834), .ZN(new_n835));
  OR3_X1    g0635(.A1(new_n821), .A2(KEYINPUT104), .A3(G190), .ZN(new_n836));
  OAI21_X1  g0636(.A(KEYINPUT104), .B1(new_n821), .B2(G190), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(G68), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n227), .B1(new_n396), .B2(new_n830), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(new_n444), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT32), .ZN(new_n842));
  NOR3_X1   g0642(.A1(G179), .A2(G190), .A3(G200), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n284), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n842), .B1(new_n844), .B2(new_n268), .ZN(new_n845));
  INV_X1    g0645(.A(new_n844), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n846), .A2(KEYINPUT32), .A3(G159), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n256), .B(new_n841), .C1(new_n845), .C2(new_n847), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n823), .A2(new_n835), .A3(new_n839), .A4(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n818), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n850), .A2(G283), .B1(G329), .B2(new_n846), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT105), .ZN(new_n852));
  INV_X1    g0652(.A(G311), .ZN(new_n853));
  INV_X1    g0653(.A(G294), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n833), .A2(new_n853), .B1(new_n840), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n828), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n855), .B1(new_n856), .B2(G303), .ZN(new_n857));
  INV_X1    g0657(.A(G322), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n256), .B1(new_n831), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(G326), .B2(new_n822), .ZN(new_n860));
  INV_X1    g0660(.A(new_n838), .ZN(new_n861));
  XOR2_X1   g0661(.A(KEYINPUT33), .B(G317), .Z(new_n862));
  OAI211_X1 g0662(.A(new_n857), .B(new_n860), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n849), .B1(new_n852), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n813), .B1(new_n864), .B2(new_n810), .ZN(new_n865));
  INV_X1    g0665(.A(new_n809), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n865), .B1(new_n789), .B2(new_n866), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n795), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(G396));
  NAND2_X1  g0669(.A1(new_n414), .A2(new_n420), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n706), .B1(new_n870), .B2(new_n425), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n421), .A2(new_n426), .B1(new_n398), .B2(new_n407), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n427), .A2(new_n871), .B1(new_n872), .B2(new_n429), .ZN(new_n873));
  AND4_X1   g0673(.A1(new_n428), .A2(new_n429), .A3(new_n430), .A4(new_n720), .ZN(new_n874));
  NOR3_X1   g0674(.A1(new_n873), .A2(KEYINPUT107), .A3(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT107), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n427), .A2(new_n871), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n431), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n872), .A2(new_n429), .A3(new_n720), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n876), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n745), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT108), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n875), .B2(new_n880), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT107), .B1(new_n873), .B2(new_n874), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n878), .A2(new_n876), .A3(new_n879), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n886), .A2(KEYINPUT108), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n883), .B1(new_n745), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n796), .B1(new_n890), .B2(new_n785), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n785), .B2(new_n890), .ZN(new_n892));
  INV_X1    g0692(.A(new_n810), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n808), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n796), .B1(G77), .B2(new_n894), .ZN(new_n895));
  OAI22_X1  g0695(.A1(new_n490), .A2(new_n833), .B1(new_n831), .B2(new_n854), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n850), .A2(G87), .ZN(new_n897));
  INV_X1    g0697(.A(new_n841), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n822), .A2(G303), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n258), .B1(new_n846), .B2(G311), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n897), .A2(new_n898), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  AOI211_X1 g0701(.A(new_n896), .B(new_n901), .C1(G107), .C2(new_n856), .ZN(new_n902));
  INV_X1    g0702(.A(G283), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n861), .A2(KEYINPUT106), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n836), .A2(KEYINPUT106), .A3(new_n837), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n902), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n833), .ZN(new_n908));
  INV_X1    g0708(.A(new_n831), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n908), .A2(G159), .B1(new_n909), .B2(G143), .ZN(new_n910));
  INV_X1    g0710(.A(G137), .ZN(new_n911));
  INV_X1    g0711(.A(new_n822), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(G150), .B2(new_n838), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n914), .A2(KEYINPUT34), .ZN(new_n915));
  INV_X1    g0715(.A(G132), .ZN(new_n916));
  INV_X1    g0716(.A(G50), .ZN(new_n917));
  OAI221_X1 g0717(.A(new_n258), .B1(new_n916), .B2(new_n844), .C1(new_n828), .C2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n818), .A2(new_n209), .ZN(new_n919));
  INV_X1    g0719(.A(new_n840), .ZN(new_n920));
  AOI211_X1 g0720(.A(new_n918), .B(new_n919), .C1(G58), .C2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n914), .A2(KEYINPUT34), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n915), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n907), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n895), .B1(new_n924), .B2(new_n810), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n808), .B2(new_n882), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n892), .A2(new_n926), .ZN(G384));
  INV_X1    g0727(.A(new_n548), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n928), .A2(KEYINPUT35), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(KEYINPUT35), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n929), .A2(new_n930), .A3(G116), .A4(new_n229), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n931), .B(KEYINPUT36), .Z(new_n932));
  NAND3_X1  g0732(.A1(new_n233), .A2(G77), .A3(new_n264), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n201), .A2(new_n203), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(G68), .ZN(new_n936));
  AOI211_X1 g0736(.A(G13), .B(new_n311), .C1(new_n933), .C2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n932), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n747), .A2(new_n759), .A3(new_n483), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n939), .A2(new_n682), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n351), .B1(KEYINPUT16), .B2(new_n350), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n313), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n355), .ZN(new_n943));
  INV_X1    g0743(.A(new_n704), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n943), .A2(new_n945), .A3(new_n341), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(KEYINPUT37), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n301), .A2(new_n313), .A3(new_n340), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n948), .A2(new_n360), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT37), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n301), .A2(new_n313), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n944), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n949), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n947), .A2(new_n953), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n954), .B(KEYINPUT38), .C1(new_n363), .C2(new_n945), .ZN(new_n955));
  XOR2_X1   g0755(.A(KEYINPUT109), .B(KEYINPUT38), .Z(new_n956));
  AOI21_X1  g0756(.A(new_n950), .B1(new_n949), .B2(new_n952), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n951), .A2(new_n355), .ZN(new_n958));
  AND4_X1   g0758(.A1(new_n950), .A2(new_n958), .A3(new_n952), .A4(new_n341), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n341), .B(KEYINPUT17), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n360), .A2(KEYINPUT18), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n357), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n952), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n956), .B1(new_n960), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n955), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT39), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n954), .B1(new_n363), .B2(new_n945), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT38), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n971), .A2(KEYINPUT39), .A3(new_n955), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n462), .A2(new_n476), .A3(new_n720), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n968), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n476), .A2(new_n706), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n477), .A2(new_n481), .A3(new_n976), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n476), .B(new_n706), .C1(new_n462), .C2(new_n480), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n980), .B1(new_n883), .B2(new_n879), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n971), .A2(new_n955), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n677), .A2(new_n704), .ZN(new_n984));
  AND3_X1   g0784(.A1(new_n975), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n940), .B(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n956), .ZN(new_n987));
  INV_X1    g0787(.A(new_n952), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n677), .B2(new_n343), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n958), .A2(new_n952), .A3(new_n341), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(KEYINPUT37), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n953), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n987), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(KEYINPUT77), .B1(new_n360), .B2(KEYINPUT18), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n994), .A2(new_n676), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n961), .B1(new_n995), .B2(new_n361), .ZN(new_n996));
  INV_X1    g0796(.A(new_n945), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n996), .A2(new_n997), .B1(new_n953), .B2(new_n947), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n993), .B1(new_n998), .B2(KEYINPUT38), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n881), .B1(new_n977), .B2(new_n978), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n781), .A2(new_n684), .A3(new_n685), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT110), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n778), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n777), .A2(KEYINPUT110), .A3(new_n706), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1003), .A2(new_n779), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n780), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1001), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1000), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(KEYINPUT40), .B1(new_n999), .B2(new_n1008), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n1000), .A2(new_n1007), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT40), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n996), .A2(new_n997), .ZN(new_n1012));
  AOI21_X1  g0812(.A(KEYINPUT38), .B1(new_n1012), .B2(new_n954), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n955), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1010), .B(new_n1011), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1009), .A2(new_n1015), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n483), .A2(new_n1007), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n761), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n1017), .B2(new_n1016), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n986), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n311), .B2(new_n792), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n986), .A2(new_n1019), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n938), .B1(new_n1021), .B2(new_n1022), .ZN(G367));
  NAND2_X1  g0823(.A1(new_n801), .A2(new_n243), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n812), .B1(new_n735), .B2(new_n662), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n794), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n633), .A2(new_n653), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n706), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n694), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n667), .B2(new_n1028), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n828), .A2(new_n490), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT46), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n909), .A2(G303), .B1(new_n920), .B2(G107), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n903), .B2(new_n833), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(KEYINPUT111), .B(G317), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n258), .B1(new_n846), .B2(new_n1036), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n444), .B2(new_n815), .C1(new_n912), .C2(new_n853), .ZN(new_n1038));
  NOR3_X1   g0838(.A1(new_n1032), .A2(new_n1034), .A3(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n854), .B2(new_n906), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n833), .A2(new_n935), .B1(new_n911), .B2(new_n844), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n822), .A2(G143), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n258), .B1(new_n815), .B2(new_n419), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT112), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1042), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1041), .B(new_n1045), .C1(new_n1044), .C2(new_n1043), .ZN(new_n1046));
  INV_X1    g0846(.A(G150), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n828), .A2(new_n230), .B1(new_n1047), .B2(new_n831), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(G68), .B2(new_n920), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1046), .B(new_n1049), .C1(new_n906), .C2(new_n268), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1040), .A2(new_n1050), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT47), .Z(new_n1052));
  OAI221_X1 g0852(.A(new_n1026), .B1(new_n866), .B2(new_n1030), .C1(new_n1052), .C2(new_n893), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n736), .B(KEYINPUT41), .Z(new_n1054));
  INV_X1    g0854(.A(new_n695), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n557), .A2(new_n706), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1055), .A2(new_n581), .A3(new_n1056), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n574), .A2(new_n720), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n733), .B2(new_n731), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT45), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  OAI211_X1 g0862(.A(KEYINPUT45), .B(new_n1059), .C1(new_n733), .C2(new_n731), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n731), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1059), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1065), .A2(new_n732), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT44), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1065), .A2(KEYINPUT44), .A3(new_n732), .A4(new_n1066), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1064), .A2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n713), .A2(new_n726), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n729), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n713), .A2(new_n726), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1075), .B1(new_n1077), .B2(new_n1073), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n728), .A2(new_n1076), .A3(new_n729), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1080), .A2(new_n786), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1064), .A2(new_n1071), .A3(new_n728), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1074), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1054), .B1(new_n1083), .B2(new_n787), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n793), .A2(G1), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n727), .A2(new_n729), .A3(new_n1059), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1055), .B1(new_n1066), .B2(new_n685), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1087), .A2(KEYINPUT42), .B1(new_n1088), .B2(new_n720), .ZN(new_n1089));
  OR2_X1    g0889(.A1(new_n1087), .A2(KEYINPUT42), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n1089), .A2(new_n1090), .B1(KEYINPUT43), .B2(new_n1030), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1030), .A2(KEYINPUT43), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1091), .B(new_n1092), .Z(new_n1093));
  NOR2_X1   g0893(.A1(new_n728), .A2(new_n1066), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1093), .B(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1053), .B1(new_n1086), .B2(new_n1096), .ZN(G387));
  INV_X1    g0897(.A(new_n736), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1081), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1080), .A2(new_n786), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1080), .B1(G1), .B2(new_n793), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n258), .B1(new_n846), .B2(G326), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n490), .B2(new_n815), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n908), .A2(G303), .B1(new_n909), .B2(new_n1036), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n906), .A2(new_n853), .B1(new_n858), .B2(new_n912), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1106), .B1(new_n1107), .B2(KEYINPUT113), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT114), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT113), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1110), .B1(new_n858), .B2(new_n912), .C1(new_n906), .C2(new_n853), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1108), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1109), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1114));
  OAI21_X1  g0914(.A(KEYINPUT48), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1114), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT48), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(new_n1117), .A3(new_n1112), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n856), .A2(G294), .B1(G283), .B2(new_n920), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1115), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT49), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1104), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1115), .A2(new_n1118), .A3(KEYINPUT49), .A4(new_n1119), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n840), .A2(new_n412), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(G68), .B2(new_n908), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n917), .B2(new_n831), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n258), .B1(new_n844), .B2(new_n1047), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n856), .B2(G77), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(new_n444), .B2(new_n818), .C1(new_n268), .C2(new_n912), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1127), .B(new_n1130), .C1(new_n303), .C2(new_n838), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n810), .B1(new_n1124), .B2(new_n1131), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n797), .A2(new_n738), .B1(G107), .B2(new_n222), .ZN(new_n1133));
  OR2_X1    g0933(.A1(new_n240), .A2(new_n803), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n738), .ZN(new_n1135));
  AOI211_X1 g0935(.A(G45), .B(new_n1135), .C1(G68), .C2(G77), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n410), .A2(G50), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT50), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n802), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1133), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n796), .B1(new_n1140), .B2(new_n812), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n726), .B2(new_n809), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1102), .B1(new_n1132), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1101), .A2(new_n1143), .ZN(G393));
  AND2_X1   g0944(.A1(new_n1083), .A2(new_n736), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n1074), .A2(new_n1082), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1145), .B1(new_n1081), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1066), .A2(new_n809), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n811), .B1(new_n444), .B2(new_n222), .C1(new_n802), .C2(new_n250), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n796), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n256), .B1(new_n846), .B2(G143), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n897), .B(new_n1151), .C1(new_n209), .C2(new_n828), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT116), .ZN(new_n1153));
  OR2_X1    g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n822), .A2(G150), .B1(new_n909), .B2(G159), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  XOR2_X1   g0956(.A(KEYINPUT115), .B(KEYINPUT51), .Z(new_n1157));
  NOR2_X1   g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n906), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n934), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n833), .A2(new_n410), .B1(new_n840), .B2(new_n419), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1154), .A2(new_n1159), .A3(new_n1161), .A4(new_n1163), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n256), .B1(new_n844), .B2(new_n858), .C1(new_n840), .C2(new_n490), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n828), .A2(new_n903), .B1(new_n854), .B2(new_n833), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n819), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n822), .A2(G317), .B1(new_n909), .B2(G311), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT52), .Z(new_n1169));
  INV_X1    g0969(.A(G303), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1167), .B(new_n1169), .C1(new_n906), .C2(new_n1170), .ZN(new_n1171));
  OR2_X1    g0971(.A1(new_n1171), .A2(KEYINPUT117), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(KEYINPUT117), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1164), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1150), .B1(new_n1174), .B2(new_n810), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n1146), .A2(new_n1085), .B1(new_n1148), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1147), .A2(new_n1176), .ZN(G390));
  AOI21_X1  g0977(.A(new_n761), .B1(new_n782), .B2(new_n1005), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n483), .A2(new_n1178), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n939), .A2(new_n682), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1178), .A2(new_n1000), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n979), .B1(new_n784), .B2(new_n882), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n706), .B(new_n881), .C1(new_n687), .C2(new_n697), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n1182), .A2(new_n1183), .B1(new_n874), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1007), .A2(G330), .A3(new_n889), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1186), .A2(KEYINPUT118), .A3(new_n980), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n706), .B1(new_n755), .B2(new_n687), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n874), .B1(new_n1188), .B2(new_n882), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n784), .A2(new_n882), .A3(new_n979), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1187), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(KEYINPUT118), .B1(new_n1186), .B2(new_n980), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1185), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1180), .A2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n979), .B1(new_n1184), .B2(new_n874), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1195), .A2(new_n973), .B1(new_n968), .B2(new_n972), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n966), .A2(new_n973), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n720), .B1(new_n749), .B2(new_n752), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n879), .B1(new_n1198), .B2(new_n881), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1197), .B1(new_n979), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1190), .ZN(new_n1201));
  NOR3_X1   g1001(.A1(new_n1196), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n971), .A2(KEYINPUT39), .A3(new_n955), .ZN(new_n1203));
  AOI21_X1  g1003(.A(KEYINPUT39), .B1(new_n955), .B2(new_n965), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n1203), .A2(new_n1204), .B1(new_n981), .B2(new_n974), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n973), .B(new_n966), .C1(new_n1189), .C2(new_n980), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1181), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1194), .B1(new_n1202), .B2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1182), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1205), .A2(new_n1206), .A3(new_n1190), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1209), .A2(new_n1180), .A3(new_n1210), .A4(new_n1193), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1208), .A2(new_n736), .A3(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1202), .A2(new_n1207), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n807), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n796), .B1(new_n303), .B2(new_n894), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n258), .B(new_n829), .C1(G294), .C2(new_n846), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n919), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n831), .A2(new_n490), .B1(new_n840), .B2(new_n419), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G97), .B2(new_n908), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n822), .A2(G283), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1216), .A2(new_n1217), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n906), .A2(new_n540), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n906), .A2(new_n911), .ZN(new_n1223));
  OR3_X1    g1023(.A1(new_n828), .A2(KEYINPUT53), .A3(new_n1047), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n256), .B1(new_n846), .B2(G125), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n935), .B2(new_n815), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G128), .B2(new_n822), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n831), .A2(new_n916), .B1(new_n840), .B2(new_n268), .ZN(new_n1228));
  XOR2_X1   g1028(.A(KEYINPUT54), .B(G143), .Z(new_n1229));
  AOI21_X1  g1029(.A(new_n1228), .B1(new_n908), .B2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(KEYINPUT53), .B1(new_n828), .B2(new_n1047), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1224), .A2(new_n1227), .A3(new_n1230), .A4(new_n1231), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n1221), .A2(new_n1222), .B1(new_n1223), .B2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1215), .B1(new_n1233), .B2(new_n810), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1213), .A2(new_n1085), .B1(new_n1214), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1212), .A2(new_n1235), .ZN(G378));
  NAND3_X1  g1036(.A1(new_n975), .A2(new_n983), .A3(new_n984), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n401), .B1(new_n678), .B2(new_n679), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n944), .A2(new_n400), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n401), .B(new_n1239), .C1(new_n678), .C2(new_n679), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1243), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n1016), .B2(G330), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n761), .B(new_n1246), .C1(new_n1009), .C2(new_n1015), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1237), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT40), .B1(new_n971), .B2(new_n955), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1010), .A2(new_n966), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1010), .A2(new_n1251), .B1(new_n1252), .B2(KEYINPUT40), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1246), .B1(new_n1253), .B2(new_n761), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1016), .A2(new_n1247), .A3(G330), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(new_n985), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1250), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1246), .A2(new_n807), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n796), .B1(new_n934), .B2(new_n894), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n258), .A2(G41), .ZN(new_n1260));
  INV_X1    g1060(.A(G41), .ZN(new_n1261));
  AOI211_X1 g1061(.A(G50), .B(new_n1260), .C1(new_n266), .C2(new_n1261), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n831), .A2(new_n540), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1263), .B(KEYINPUT119), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n828), .A2(new_n419), .B1(new_n412), .B2(new_n833), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n1260), .B1(new_n903), .B2(new_n844), .C1(new_n815), .C2(new_n230), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n822), .A2(G116), .B1(G68), .B2(new_n920), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(new_n1268), .B(KEYINPUT120), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1267), .B(new_n1269), .C1(new_n444), .C2(new_n861), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT58), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1262), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(KEYINPUT121), .B1(new_n856), .B2(new_n1229), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(G125), .B2(new_n822), .ZN(new_n1274));
  OAI22_X1  g1074(.A1(new_n833), .A2(new_n911), .B1(new_n840), .B2(new_n1047), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(G128), .B2(new_n909), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n856), .A2(KEYINPUT121), .A3(new_n1229), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1274), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1278), .B1(G132), .B2(new_n838), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1280), .A2(KEYINPUT59), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n266), .B(new_n1261), .C1(new_n815), .C2(new_n268), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1282), .B1(G124), .B2(new_n846), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT59), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1283), .B1(new_n1279), .B2(new_n1284), .ZN(new_n1285));
  OAI221_X1 g1085(.A(new_n1272), .B1(new_n1271), .B2(new_n1270), .C1(new_n1281), .C2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1259), .B1(new_n1286), .B2(new_n810), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1257), .A2(new_n1085), .B1(new_n1258), .B2(new_n1287), .ZN(new_n1288));
  NOR3_X1   g1088(.A1(new_n1248), .A2(new_n1249), .A3(new_n1237), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n985), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1290));
  OAI21_X1  g1090(.A(KEYINPUT57), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n939), .A2(new_n682), .A3(new_n1179), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1292), .B1(new_n1213), .B2(new_n1193), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n736), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1211), .A2(new_n1180), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT57), .B1(new_n1295), .B2(new_n1257), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1288), .B1(new_n1294), .B2(new_n1296), .ZN(G375));
  NAND2_X1  g1097(.A1(new_n980), .A2(new_n807), .ZN(new_n1298));
  OAI22_X1  g1098(.A1(new_n828), .A2(new_n444), .B1(new_n903), .B2(new_n831), .ZN(new_n1299));
  AOI211_X1 g1099(.A(new_n258), .B(new_n1125), .C1(G303), .C2(new_n846), .ZN(new_n1300));
  OAI221_X1 g1100(.A(new_n1300), .B1(new_n854), .B2(new_n912), .C1(new_n818), .C2(new_n419), .ZN(new_n1301));
  AOI211_X1 g1101(.A(new_n1299), .B(new_n1301), .C1(G107), .C2(new_n908), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1160), .A2(G116), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1160), .A2(new_n1229), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n846), .A2(G128), .ZN(new_n1305));
  OAI211_X1 g1105(.A(new_n258), .B(new_n1305), .C1(new_n815), .C2(new_n230), .ZN(new_n1306));
  AOI22_X1  g1106(.A1(new_n908), .A2(G150), .B1(new_n909), .B2(G137), .ZN(new_n1307));
  OAI221_X1 g1107(.A(new_n1307), .B1(new_n917), .B2(new_n840), .C1(new_n268), .C2(new_n828), .ZN(new_n1308));
  AOI211_X1 g1108(.A(new_n1306), .B(new_n1308), .C1(G132), .C2(new_n822), .ZN(new_n1309));
  AOI22_X1  g1109(.A1(new_n1302), .A2(new_n1303), .B1(new_n1304), .B2(new_n1309), .ZN(new_n1310));
  OAI221_X1 g1110(.A(new_n796), .B1(G68), .B2(new_n894), .C1(new_n1310), .C2(new_n893), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(new_n1311), .B(KEYINPUT122), .ZN(new_n1312));
  AOI22_X1  g1112(.A1(new_n1193), .A2(new_n1085), .B1(new_n1298), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1054), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1194), .A2(new_n1314), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1180), .A2(new_n1193), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1313), .B1(new_n1315), .B2(new_n1316), .ZN(G381));
  AND3_X1   g1117(.A1(new_n1101), .A2(new_n1143), .A3(new_n868), .ZN(new_n1318));
  INV_X1    g1118(.A(G384), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  XOR2_X1   g1120(.A(new_n1320), .B(KEYINPUT123), .Z(new_n1321));
  NOR3_X1   g1121(.A1(G390), .A2(G378), .A3(G381), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(G387), .A2(G375), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1321), .A2(new_n1322), .A3(new_n1323), .ZN(G407));
  INV_X1    g1124(.A(G213), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1325), .A2(G343), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  NOR3_X1   g1127(.A1(G375), .A2(G378), .A3(new_n1327), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(new_n1328), .B(KEYINPUT124), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1329), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1130(.A(G390), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n868), .B1(new_n1101), .B2(new_n1143), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1318), .A2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT126), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1333), .B1(G387), .B2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(G393), .A2(G396), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1101), .A2(new_n1143), .A3(new_n868), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  XNOR2_X1  g1138(.A(new_n1093), .B(new_n1094), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1339), .B1(new_n1085), .B2(new_n1084), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1338), .B1(new_n1340), .B2(new_n1053), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1331), .B1(new_n1335), .B2(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(G387), .A2(new_n1333), .ZN(new_n1343));
  AOI21_X1  g1143(.A(KEYINPUT126), .B1(new_n1340), .B2(new_n1053), .ZN(new_n1344));
  OAI211_X1 g1144(.A(new_n1343), .B(G390), .C1(new_n1344), .C2(new_n1333), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1342), .A2(new_n1345), .ZN(new_n1346));
  OAI211_X1 g1146(.A(G378), .B(new_n1288), .C1(new_n1294), .C2(new_n1296), .ZN(new_n1347));
  AND2_X1   g1147(.A1(new_n1212), .A2(new_n1235), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1295), .A2(new_n1257), .A3(new_n1314), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1288), .A2(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1348), .A2(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1347), .A2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1352), .A2(new_n1327), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1326), .A2(G2897), .ZN(new_n1354));
  NOR2_X1   g1154(.A1(new_n1319), .A2(KEYINPUT125), .ZN(new_n1355));
  AND3_X1   g1155(.A1(new_n892), .A2(KEYINPUT125), .A3(new_n926), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT60), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1357), .B1(new_n1180), .B2(new_n1193), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1098), .B1(new_n1180), .B2(new_n1193), .ZN(new_n1359));
  OR2_X1    g1159(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1360));
  NAND4_X1  g1160(.A1(new_n1292), .A2(new_n1360), .A3(KEYINPUT60), .A4(new_n1185), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1358), .A2(new_n1359), .A3(new_n1361), .ZN(new_n1362));
  AOI211_X1 g1162(.A(new_n1355), .B(new_n1356), .C1(new_n1362), .C2(new_n1313), .ZN(new_n1363));
  NAND4_X1  g1163(.A1(new_n1362), .A2(KEYINPUT125), .A3(new_n1319), .A4(new_n1313), .ZN(new_n1364));
  INV_X1    g1164(.A(new_n1364), .ZN(new_n1365));
  OAI21_X1  g1165(.A(new_n1354), .B1(new_n1363), .B2(new_n1365), .ZN(new_n1366));
  AOI21_X1  g1166(.A(new_n1355), .B1(new_n1362), .B2(new_n1313), .ZN(new_n1367));
  INV_X1    g1167(.A(new_n1356), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1367), .A2(new_n1368), .ZN(new_n1369));
  INV_X1    g1169(.A(new_n1354), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1369), .A2(new_n1364), .A3(new_n1370), .ZN(new_n1371));
  AND2_X1   g1171(.A1(new_n1366), .A2(new_n1371), .ZN(new_n1372));
  AOI21_X1  g1172(.A(KEYINPUT61), .B1(new_n1353), .B2(new_n1372), .ZN(new_n1373));
  INV_X1    g1173(.A(KEYINPUT63), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1369), .A2(new_n1364), .ZN(new_n1375));
  INV_X1    g1175(.A(new_n1375), .ZN(new_n1376));
  OAI21_X1  g1176(.A(new_n1374), .B1(new_n1353), .B2(new_n1376), .ZN(new_n1377));
  AOI21_X1  g1177(.A(new_n1326), .B1(new_n1347), .B2(new_n1351), .ZN(new_n1378));
  NAND3_X1  g1178(.A1(new_n1378), .A2(KEYINPUT63), .A3(new_n1375), .ZN(new_n1379));
  NAND4_X1  g1179(.A1(new_n1346), .A2(new_n1373), .A3(new_n1377), .A4(new_n1379), .ZN(new_n1380));
  INV_X1    g1180(.A(KEYINPUT62), .ZN(new_n1381));
  AND3_X1   g1181(.A1(new_n1378), .A2(new_n1381), .A3(new_n1375), .ZN(new_n1382));
  INV_X1    g1182(.A(KEYINPUT61), .ZN(new_n1383));
  NAND2_X1  g1183(.A1(new_n1366), .A2(new_n1371), .ZN(new_n1384));
  OAI21_X1  g1184(.A(new_n1383), .B1(new_n1378), .B2(new_n1384), .ZN(new_n1385));
  AOI21_X1  g1185(.A(new_n1381), .B1(new_n1378), .B2(new_n1375), .ZN(new_n1386));
  NOR3_X1   g1186(.A1(new_n1382), .A2(new_n1385), .A3(new_n1386), .ZN(new_n1387));
  OAI21_X1  g1187(.A(new_n1380), .B1(new_n1387), .B2(new_n1346), .ZN(G405));
  NAND2_X1  g1188(.A1(new_n1375), .A2(KEYINPUT127), .ZN(new_n1389));
  NAND2_X1  g1189(.A1(G375), .A2(new_n1348), .ZN(new_n1390));
  AND3_X1   g1190(.A1(new_n1389), .A2(new_n1390), .A3(new_n1347), .ZN(new_n1391));
  AOI21_X1  g1191(.A(new_n1389), .B1(new_n1390), .B2(new_n1347), .ZN(new_n1392));
  NOR2_X1   g1192(.A1(new_n1391), .A2(new_n1392), .ZN(new_n1393));
  XNOR2_X1  g1193(.A(new_n1393), .B(new_n1346), .ZN(G402));
endmodule


