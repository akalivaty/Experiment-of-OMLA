

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U550 ( .A1(n980), .A2(n709), .ZN(n710) );
  NOR2_X1 U551 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  BUF_X2 U552 ( .A(n882), .Z(n516) );
  XOR2_X1 U553 ( .A(KEYINPUT17), .B(n526), .Z(n882) );
  NAND2_X1 U554 ( .A1(n522), .A2(n713), .ZN(n521) );
  NOR2_X1 U555 ( .A1(G164), .A2(G1384), .ZN(n787) );
  NOR2_X2 U556 ( .A1(n536), .A2(n535), .ZN(G160) );
  XNOR2_X1 U557 ( .A(n517), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U558 ( .A1(n518), .A2(n832), .ZN(n517) );
  NAND2_X1 U559 ( .A1(n519), .A2(n523), .ZN(n518) );
  XNOR2_X1 U560 ( .A(n785), .B(KEYINPUT103), .ZN(n519) );
  NAND2_X1 U561 ( .A1(n520), .A2(n719), .ZN(n724) );
  NAND2_X1 U562 ( .A1(n715), .A2(n521), .ZN(n520) );
  OR2_X2 U563 ( .A1(n714), .A2(n975), .ZN(n522) );
  NAND2_X1 U564 ( .A1(n524), .A2(n729), .ZN(n750) );
  BUF_X1 U565 ( .A(n706), .Z(n744) );
  NAND2_X1 U566 ( .A1(n703), .A2(n787), .ZN(n706) );
  AND2_X1 U567 ( .A1(n525), .A2(n820), .ZN(n523) );
  XOR2_X1 U568 ( .A(KEYINPUT29), .B(n725), .Z(n524) );
  AND2_X1 U569 ( .A1(n826), .A2(n819), .ZN(n525) );
  XOR2_X1 U570 ( .A(G651), .B(KEYINPUT68), .Z(n557) );
  NOR2_X1 U571 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U572 ( .A1(n532), .A2(G2104), .ZN(n881) );
  NOR2_X1 U573 ( .A1(G651), .A2(n657), .ZN(n669) );
  NAND2_X1 U574 ( .A1(n516), .A2(G137), .ZN(n528) );
  INV_X1 U575 ( .A(G2105), .ZN(n532) );
  AND2_X1 U576 ( .A1(G2104), .A2(G2105), .ZN(n878) );
  NAND2_X1 U577 ( .A1(G113), .A2(n878), .ZN(n527) );
  NAND2_X1 U578 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U579 ( .A(n529), .B(KEYINPUT67), .ZN(n531) );
  NOR2_X1 U580 ( .A1(G2104), .A2(n532), .ZN(n877) );
  NAND2_X1 U581 ( .A1(G125), .A2(n877), .ZN(n530) );
  NAND2_X1 U582 ( .A1(n531), .A2(n530), .ZN(n536) );
  NAND2_X1 U583 ( .A1(G101), .A2(n881), .ZN(n533) );
  XNOR2_X1 U584 ( .A(n533), .B(KEYINPUT66), .ZN(n534) );
  XNOR2_X1 U585 ( .A(n534), .B(KEYINPUT23), .ZN(n535) );
  NAND2_X1 U586 ( .A1(G102), .A2(n881), .ZN(n538) );
  NAND2_X1 U587 ( .A1(n516), .A2(G138), .ZN(n537) );
  NAND2_X1 U588 ( .A1(n538), .A2(n537), .ZN(n542) );
  NAND2_X1 U589 ( .A1(G126), .A2(n877), .ZN(n540) );
  NAND2_X1 U590 ( .A1(G114), .A2(n878), .ZN(n539) );
  NAND2_X1 U591 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U592 ( .A1(n542), .A2(n541), .ZN(G164) );
  XOR2_X1 U593 ( .A(G2443), .B(G2446), .Z(n544) );
  XNOR2_X1 U594 ( .A(G2427), .B(G2451), .ZN(n543) );
  XNOR2_X1 U595 ( .A(n544), .B(n543), .ZN(n550) );
  XOR2_X1 U596 ( .A(G2430), .B(G2454), .Z(n546) );
  XNOR2_X1 U597 ( .A(G1348), .B(G1341), .ZN(n545) );
  XNOR2_X1 U598 ( .A(n546), .B(n545), .ZN(n548) );
  XOR2_X1 U599 ( .A(G2435), .B(G2438), .Z(n547) );
  XNOR2_X1 U600 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U601 ( .A(n550), .B(n549), .Z(n551) );
  AND2_X1 U602 ( .A1(G14), .A2(n551), .ZN(G401) );
  XOR2_X1 U603 ( .A(KEYINPUT0), .B(G543), .Z(n657) );
  NAND2_X1 U604 ( .A1(G52), .A2(n669), .ZN(n552) );
  XNOR2_X1 U605 ( .A(n552), .B(KEYINPUT71), .ZN(n563) );
  NOR2_X1 U606 ( .A1(G651), .A2(G543), .ZN(n553) );
  XOR2_X1 U607 ( .A(KEYINPUT65), .B(n553), .Z(n580) );
  BUF_X1 U608 ( .A(n580), .Z(n664) );
  NAND2_X1 U609 ( .A1(G90), .A2(n664), .ZN(n555) );
  NOR2_X1 U610 ( .A1(n657), .A2(n557), .ZN(n668) );
  NAND2_X1 U611 ( .A1(G77), .A2(n668), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U613 ( .A(n556), .B(KEYINPUT9), .ZN(n561) );
  XNOR2_X1 U614 ( .A(KEYINPUT1), .B(KEYINPUT69), .ZN(n559) );
  NOR2_X1 U615 ( .A1(G543), .A2(n557), .ZN(n558) );
  XNOR2_X2 U616 ( .A(n559), .B(n558), .ZN(n665) );
  NAND2_X1 U617 ( .A1(G64), .A2(n665), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U619 ( .A1(n563), .A2(n562), .ZN(G171) );
  AND2_X1 U620 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U621 ( .A(G57), .ZN(G237) );
  INV_X1 U622 ( .A(G132), .ZN(G219) );
  INV_X1 U623 ( .A(G82), .ZN(G220) );
  NAND2_X1 U624 ( .A1(G89), .A2(n664), .ZN(n564) );
  XOR2_X1 U625 ( .A(KEYINPUT77), .B(n564), .Z(n565) );
  XNOR2_X1 U626 ( .A(n565), .B(KEYINPUT4), .ZN(n567) );
  NAND2_X1 U627 ( .A1(G76), .A2(n668), .ZN(n566) );
  NAND2_X1 U628 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U629 ( .A(KEYINPUT5), .B(n568), .ZN(n574) );
  NAND2_X1 U630 ( .A1(G63), .A2(n665), .ZN(n570) );
  NAND2_X1 U631 ( .A1(G51), .A2(n669), .ZN(n569) );
  NAND2_X1 U632 ( .A1(n570), .A2(n569), .ZN(n572) );
  XOR2_X1 U633 ( .A(KEYINPUT78), .B(KEYINPUT6), .Z(n571) );
  XNOR2_X1 U634 ( .A(n572), .B(n571), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U636 ( .A(KEYINPUT7), .B(n575), .ZN(G168) );
  XOR2_X1 U637 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U638 ( .A1(G7), .A2(G661), .ZN(n576) );
  XNOR2_X1 U639 ( .A(n576), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U640 ( .A(KEYINPUT72), .B(KEYINPUT11), .Z(n578) );
  INV_X1 U641 ( .A(G223), .ZN(n833) );
  NAND2_X1 U642 ( .A1(G567), .A2(n833), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G234) );
  NAND2_X1 U644 ( .A1(n665), .A2(G56), .ZN(n579) );
  XOR2_X1 U645 ( .A(KEYINPUT14), .B(n579), .Z(n589) );
  INV_X1 U646 ( .A(KEYINPUT13), .ZN(n587) );
  INV_X1 U647 ( .A(KEYINPUT73), .ZN(n582) );
  NAND2_X1 U648 ( .A1(G81), .A2(n580), .ZN(n581) );
  XNOR2_X1 U649 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n583), .B(KEYINPUT12), .ZN(n585) );
  NAND2_X1 U651 ( .A1(G68), .A2(n668), .ZN(n584) );
  NAND2_X1 U652 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U653 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n590), .B(KEYINPUT74), .ZN(n592) );
  NAND2_X1 U655 ( .A1(G43), .A2(n669), .ZN(n591) );
  NAND2_X1 U656 ( .A1(n592), .A2(n591), .ZN(n980) );
  INV_X1 U657 ( .A(G860), .ZN(n638) );
  OR2_X1 U658 ( .A1(n980), .A2(n638), .ZN(G153) );
  INV_X1 U659 ( .A(G171), .ZN(G301) );
  NAND2_X1 U660 ( .A1(G54), .A2(n669), .ZN(n599) );
  NAND2_X1 U661 ( .A1(G79), .A2(n668), .ZN(n594) );
  NAND2_X1 U662 ( .A1(G66), .A2(n665), .ZN(n593) );
  NAND2_X1 U663 ( .A1(n594), .A2(n593), .ZN(n597) );
  NAND2_X1 U664 ( .A1(G92), .A2(n664), .ZN(n595) );
  XNOR2_X1 U665 ( .A(KEYINPUT75), .B(n595), .ZN(n596) );
  NOR2_X1 U666 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U667 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U668 ( .A(n600), .B(KEYINPUT15), .ZN(n601) );
  XNOR2_X1 U669 ( .A(KEYINPUT76), .B(n601), .ZN(n636) );
  INV_X1 U670 ( .A(n636), .ZN(n975) );
  NOR2_X1 U671 ( .A1(n975), .A2(G868), .ZN(n603) );
  INV_X1 U672 ( .A(G868), .ZN(n686) );
  NOR2_X1 U673 ( .A1(n686), .A2(G301), .ZN(n602) );
  NOR2_X1 U674 ( .A1(n603), .A2(n602), .ZN(G284) );
  NAND2_X1 U675 ( .A1(G65), .A2(n665), .ZN(n605) );
  NAND2_X1 U676 ( .A1(G53), .A2(n669), .ZN(n604) );
  NAND2_X1 U677 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U678 ( .A1(G91), .A2(n664), .ZN(n607) );
  NAND2_X1 U679 ( .A1(G78), .A2(n668), .ZN(n606) );
  NAND2_X1 U680 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U681 ( .A1(n609), .A2(n608), .ZN(n983) );
  INV_X1 U682 ( .A(n983), .ZN(G299) );
  NOR2_X1 U683 ( .A1(G286), .A2(n686), .ZN(n611) );
  NOR2_X1 U684 ( .A1(G868), .A2(G299), .ZN(n610) );
  NOR2_X1 U685 ( .A1(n611), .A2(n610), .ZN(G297) );
  NAND2_X1 U686 ( .A1(n638), .A2(G559), .ZN(n612) );
  NAND2_X1 U687 ( .A1(n612), .A2(n636), .ZN(n613) );
  XNOR2_X1 U688 ( .A(n613), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U689 ( .A1(G868), .A2(n980), .ZN(n616) );
  NAND2_X1 U690 ( .A1(n636), .A2(G868), .ZN(n614) );
  NOR2_X1 U691 ( .A1(G559), .A2(n614), .ZN(n615) );
  NOR2_X1 U692 ( .A1(n616), .A2(n615), .ZN(G282) );
  NAND2_X1 U693 ( .A1(G123), .A2(n877), .ZN(n617) );
  XNOR2_X1 U694 ( .A(n617), .B(KEYINPUT18), .ZN(n625) );
  NAND2_X1 U695 ( .A1(n881), .A2(G99), .ZN(n618) );
  XNOR2_X1 U696 ( .A(n618), .B(KEYINPUT80), .ZN(n620) );
  NAND2_X1 U697 ( .A1(G111), .A2(n878), .ZN(n619) );
  NAND2_X1 U698 ( .A1(n620), .A2(n619), .ZN(n623) );
  NAND2_X1 U699 ( .A1(G135), .A2(n516), .ZN(n621) );
  XNOR2_X1 U700 ( .A(KEYINPUT79), .B(n621), .ZN(n622) );
  NOR2_X1 U701 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n919) );
  XNOR2_X1 U703 ( .A(n919), .B(G2096), .ZN(n626) );
  XNOR2_X1 U704 ( .A(n626), .B(KEYINPUT81), .ZN(n628) );
  INV_X1 U705 ( .A(G2100), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n628), .A2(n627), .ZN(G156) );
  NAND2_X1 U707 ( .A1(n664), .A2(G93), .ZN(n629) );
  XNOR2_X1 U708 ( .A(n629), .B(KEYINPUT82), .ZN(n631) );
  NAND2_X1 U709 ( .A1(G80), .A2(n668), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n635) );
  NAND2_X1 U711 ( .A1(G67), .A2(n665), .ZN(n633) );
  NAND2_X1 U712 ( .A1(G55), .A2(n669), .ZN(n632) );
  NAND2_X1 U713 ( .A1(n633), .A2(n632), .ZN(n634) );
  OR2_X1 U714 ( .A1(n635), .A2(n634), .ZN(n687) );
  NAND2_X1 U715 ( .A1(n636), .A2(G559), .ZN(n637) );
  XOR2_X1 U716 ( .A(n980), .B(n637), .Z(n684) );
  NAND2_X1 U717 ( .A1(n638), .A2(n684), .ZN(n639) );
  XNOR2_X1 U718 ( .A(n639), .B(KEYINPUT83), .ZN(n640) );
  XOR2_X1 U719 ( .A(n687), .B(n640), .Z(G145) );
  NAND2_X1 U720 ( .A1(G88), .A2(n664), .ZN(n642) );
  NAND2_X1 U721 ( .A1(G75), .A2(n668), .ZN(n641) );
  NAND2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U723 ( .A1(G62), .A2(n665), .ZN(n644) );
  NAND2_X1 U724 ( .A1(G50), .A2(n669), .ZN(n643) );
  NAND2_X1 U725 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U726 ( .A1(n646), .A2(n645), .ZN(G166) );
  INV_X1 U727 ( .A(G166), .ZN(G303) );
  NAND2_X1 U728 ( .A1(n664), .A2(G86), .ZN(n647) );
  XOR2_X1 U729 ( .A(KEYINPUT85), .B(n647), .Z(n649) );
  NAND2_X1 U730 ( .A1(n665), .A2(G61), .ZN(n648) );
  NAND2_X1 U731 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U732 ( .A(KEYINPUT86), .B(n650), .ZN(n654) );
  NAND2_X1 U733 ( .A1(G73), .A2(n668), .ZN(n651) );
  XNOR2_X1 U734 ( .A(n651), .B(KEYINPUT87), .ZN(n652) );
  XNOR2_X1 U735 ( .A(n652), .B(KEYINPUT2), .ZN(n653) );
  NOR2_X1 U736 ( .A1(n654), .A2(n653), .ZN(n656) );
  NAND2_X1 U737 ( .A1(n669), .A2(G48), .ZN(n655) );
  NAND2_X1 U738 ( .A1(n656), .A2(n655), .ZN(G305) );
  NAND2_X1 U739 ( .A1(G87), .A2(n657), .ZN(n658) );
  XNOR2_X1 U740 ( .A(n658), .B(KEYINPUT84), .ZN(n663) );
  NAND2_X1 U741 ( .A1(G49), .A2(n669), .ZN(n660) );
  NAND2_X1 U742 ( .A1(G74), .A2(G651), .ZN(n659) );
  NAND2_X1 U743 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U744 ( .A1(n665), .A2(n661), .ZN(n662) );
  NAND2_X1 U745 ( .A1(n663), .A2(n662), .ZN(G288) );
  NAND2_X1 U746 ( .A1(G85), .A2(n664), .ZN(n667) );
  NAND2_X1 U747 ( .A1(G60), .A2(n665), .ZN(n666) );
  NAND2_X1 U748 ( .A1(n667), .A2(n666), .ZN(n673) );
  NAND2_X1 U749 ( .A1(G72), .A2(n668), .ZN(n671) );
  NAND2_X1 U750 ( .A1(G47), .A2(n669), .ZN(n670) );
  NAND2_X1 U751 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U752 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U753 ( .A(KEYINPUT70), .B(n674), .Z(G290) );
  XNOR2_X1 U754 ( .A(n983), .B(G303), .ZN(n675) );
  XNOR2_X1 U755 ( .A(n675), .B(G305), .ZN(n681) );
  XNOR2_X1 U756 ( .A(KEYINPUT89), .B(KEYINPUT90), .ZN(n676) );
  XNOR2_X1 U757 ( .A(n676), .B(KEYINPUT88), .ZN(n677) );
  XNOR2_X1 U758 ( .A(KEYINPUT91), .B(n677), .ZN(n679) );
  XNOR2_X1 U759 ( .A(G288), .B(KEYINPUT19), .ZN(n678) );
  XNOR2_X1 U760 ( .A(n679), .B(n678), .ZN(n680) );
  XOR2_X1 U761 ( .A(n681), .B(n680), .Z(n683) );
  XOR2_X1 U762 ( .A(G290), .B(n687), .Z(n682) );
  XNOR2_X1 U763 ( .A(n683), .B(n682), .ZN(n904) );
  XOR2_X1 U764 ( .A(n904), .B(n684), .Z(n685) );
  NOR2_X1 U765 ( .A1(n686), .A2(n685), .ZN(n689) );
  NOR2_X1 U766 ( .A1(G868), .A2(n687), .ZN(n688) );
  NOR2_X1 U767 ( .A1(n689), .A2(n688), .ZN(G295) );
  NAND2_X1 U768 ( .A1(G2084), .A2(G2078), .ZN(n690) );
  XOR2_X1 U769 ( .A(KEYINPUT20), .B(n690), .Z(n691) );
  NAND2_X1 U770 ( .A1(G2090), .A2(n691), .ZN(n692) );
  XNOR2_X1 U771 ( .A(KEYINPUT21), .B(n692), .ZN(n693) );
  NAND2_X1 U772 ( .A1(n693), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U773 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U774 ( .A1(G220), .A2(G219), .ZN(n694) );
  XOR2_X1 U775 ( .A(KEYINPUT22), .B(n694), .Z(n695) );
  NOR2_X1 U776 ( .A1(G218), .A2(n695), .ZN(n696) );
  NAND2_X1 U777 ( .A1(G96), .A2(n696), .ZN(n837) );
  NAND2_X1 U778 ( .A1(n837), .A2(G2106), .ZN(n701) );
  NAND2_X1 U779 ( .A1(G120), .A2(G69), .ZN(n697) );
  NOR2_X1 U780 ( .A1(G237), .A2(n697), .ZN(n698) );
  NAND2_X1 U781 ( .A1(n698), .A2(G108), .ZN(n699) );
  XNOR2_X1 U782 ( .A(n699), .B(KEYINPUT92), .ZN(n838) );
  NAND2_X1 U783 ( .A1(n838), .A2(G567), .ZN(n700) );
  NAND2_X1 U784 ( .A1(n701), .A2(n700), .ZN(n839) );
  NAND2_X1 U785 ( .A1(G483), .A2(G661), .ZN(n702) );
  NOR2_X1 U786 ( .A1(n839), .A2(n702), .ZN(n836) );
  NAND2_X1 U787 ( .A1(n836), .A2(G36), .ZN(G176) );
  NAND2_X1 U788 ( .A1(G160), .A2(G40), .ZN(n786) );
  INV_X1 U789 ( .A(n786), .ZN(n703) );
  NAND2_X1 U790 ( .A1(G8), .A2(n706), .ZN(n782) );
  NOR2_X1 U791 ( .A1(G1966), .A2(n782), .ZN(n740) );
  INV_X1 U792 ( .A(G1996), .ZN(n704) );
  NOR2_X2 U793 ( .A1(n706), .A2(n704), .ZN(n705) );
  XOR2_X1 U794 ( .A(KEYINPUT26), .B(n705), .Z(n708) );
  NAND2_X1 U795 ( .A1(n744), .A2(G1341), .ZN(n707) );
  NAND2_X1 U796 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U797 ( .A(KEYINPUT64), .B(n710), .Z(n714) );
  INV_X1 U798 ( .A(n744), .ZN(n726) );
  NOR2_X1 U799 ( .A1(n726), .A2(G1348), .ZN(n712) );
  NOR2_X1 U800 ( .A1(G2067), .A2(n744), .ZN(n711) );
  NOR2_X1 U801 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U802 ( .A1(n975), .A2(n714), .ZN(n715) );
  NAND2_X1 U803 ( .A1(n726), .A2(G2072), .ZN(n716) );
  XNOR2_X1 U804 ( .A(n716), .B(KEYINPUT27), .ZN(n718) );
  INV_X1 U805 ( .A(G1956), .ZN(n998) );
  NOR2_X1 U806 ( .A1(n998), .A2(n726), .ZN(n717) );
  NOR2_X1 U807 ( .A1(n718), .A2(n717), .ZN(n720) );
  NAND2_X1 U808 ( .A1(n983), .A2(n720), .ZN(n719) );
  NOR2_X1 U809 ( .A1(n983), .A2(n720), .ZN(n722) );
  XNOR2_X1 U810 ( .A(KEYINPUT99), .B(KEYINPUT28), .ZN(n721) );
  XNOR2_X1 U811 ( .A(n722), .B(n721), .ZN(n723) );
  NAND2_X1 U812 ( .A1(n724), .A2(n723), .ZN(n725) );
  OR2_X1 U813 ( .A1(n726), .A2(G1961), .ZN(n728) );
  XNOR2_X1 U814 ( .A(G2078), .B(KEYINPUT25), .ZN(n945) );
  NAND2_X1 U815 ( .A1(n726), .A2(n945), .ZN(n727) );
  NAND2_X1 U816 ( .A1(n728), .A2(n727), .ZN(n730) );
  NAND2_X1 U817 ( .A1(n730), .A2(G171), .ZN(n729) );
  NOR2_X1 U818 ( .A1(G171), .A2(n730), .ZN(n736) );
  NOR2_X1 U819 ( .A1(G2084), .A2(n744), .ZN(n742) );
  NOR2_X1 U820 ( .A1(n742), .A2(n740), .ZN(n731) );
  NAND2_X1 U821 ( .A1(G8), .A2(n731), .ZN(n732) );
  XNOR2_X1 U822 ( .A(KEYINPUT100), .B(n732), .ZN(n733) );
  XNOR2_X1 U823 ( .A(KEYINPUT30), .B(n733), .ZN(n734) );
  NOR2_X1 U824 ( .A1(G168), .A2(n734), .ZN(n735) );
  NOR2_X1 U825 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X1 U826 ( .A(KEYINPUT31), .B(n737), .Z(n748) );
  NAND2_X1 U827 ( .A1(n750), .A2(n748), .ZN(n738) );
  XNOR2_X1 U828 ( .A(KEYINPUT101), .B(n738), .ZN(n739) );
  NOR2_X1 U829 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U830 ( .A(n741), .B(KEYINPUT102), .ZN(n765) );
  NAND2_X1 U831 ( .A1(n742), .A2(G8), .ZN(n743) );
  NAND2_X1 U832 ( .A1(n765), .A2(n743), .ZN(n757) );
  NOR2_X1 U833 ( .A1(G1971), .A2(n782), .ZN(n746) );
  NOR2_X1 U834 ( .A1(G2090), .A2(n744), .ZN(n745) );
  NOR2_X1 U835 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U836 ( .A1(n747), .A2(G303), .ZN(n751) );
  AND2_X1 U837 ( .A1(n748), .A2(n751), .ZN(n749) );
  NAND2_X1 U838 ( .A1(n750), .A2(n749), .ZN(n754) );
  INV_X1 U839 ( .A(n751), .ZN(n752) );
  OR2_X1 U840 ( .A1(n752), .A2(G286), .ZN(n753) );
  AND2_X1 U841 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U842 ( .A1(G8), .A2(n755), .ZN(n756) );
  XNOR2_X1 U843 ( .A(n756), .B(KEYINPUT32), .ZN(n768) );
  NAND2_X1 U844 ( .A1(n757), .A2(n768), .ZN(n760) );
  NOR2_X1 U845 ( .A1(G2090), .A2(G303), .ZN(n758) );
  NAND2_X1 U846 ( .A1(G8), .A2(n758), .ZN(n759) );
  NAND2_X1 U847 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U848 ( .A1(n761), .A2(n782), .ZN(n779) );
  NAND2_X1 U849 ( .A1(G1976), .A2(G288), .ZN(n970) );
  INV_X1 U850 ( .A(n782), .ZN(n762) );
  NAND2_X1 U851 ( .A1(n970), .A2(n762), .ZN(n766) );
  NOR2_X1 U852 ( .A1(G1976), .A2(G288), .ZN(n773) );
  NOR2_X1 U853 ( .A1(G1971), .A2(G303), .ZN(n763) );
  NOR2_X1 U854 ( .A1(n773), .A2(n763), .ZN(n971) );
  NOR2_X1 U855 ( .A1(n766), .A2(n971), .ZN(n764) );
  NOR2_X1 U856 ( .A1(n764), .A2(KEYINPUT33), .ZN(n769) );
  NAND2_X1 U857 ( .A1(n765), .A2(n769), .ZN(n772) );
  INV_X1 U858 ( .A(n766), .ZN(n767) );
  NAND2_X1 U859 ( .A1(n768), .A2(n767), .ZN(n770) );
  NAND2_X1 U860 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U861 ( .A1(n772), .A2(n771), .ZN(n776) );
  NAND2_X1 U862 ( .A1(n773), .A2(KEYINPUT33), .ZN(n774) );
  NOR2_X1 U863 ( .A1(n774), .A2(n782), .ZN(n775) );
  NOR2_X1 U864 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U865 ( .A(G1981), .B(G305), .Z(n967) );
  NAND2_X1 U866 ( .A1(n777), .A2(n967), .ZN(n778) );
  NAND2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n784) );
  NOR2_X1 U868 ( .A1(G1981), .A2(G305), .ZN(n780) );
  XOR2_X1 U869 ( .A(n780), .B(KEYINPUT24), .Z(n781) );
  NOR2_X1 U870 ( .A1(n782), .A2(n781), .ZN(n783) );
  NOR2_X2 U871 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U872 ( .A1(n787), .A2(n786), .ZN(n830) );
  NAND2_X1 U873 ( .A1(n516), .A2(G140), .ZN(n788) );
  XOR2_X1 U874 ( .A(KEYINPUT93), .B(n788), .Z(n790) );
  NAND2_X1 U875 ( .A1(n881), .A2(G104), .ZN(n789) );
  NAND2_X1 U876 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U877 ( .A(KEYINPUT34), .B(n791), .ZN(n796) );
  NAND2_X1 U878 ( .A1(G128), .A2(n877), .ZN(n793) );
  NAND2_X1 U879 ( .A1(G116), .A2(n878), .ZN(n792) );
  NAND2_X1 U880 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U881 ( .A(n794), .B(KEYINPUT35), .Z(n795) );
  NOR2_X1 U882 ( .A1(n796), .A2(n795), .ZN(n797) );
  XOR2_X1 U883 ( .A(KEYINPUT36), .B(n797), .Z(n798) );
  XOR2_X1 U884 ( .A(KEYINPUT94), .B(n798), .Z(n901) );
  XNOR2_X1 U885 ( .A(KEYINPUT37), .B(G2067), .ZN(n828) );
  OR2_X1 U886 ( .A1(n901), .A2(n828), .ZN(n799) );
  XNOR2_X1 U887 ( .A(n799), .B(KEYINPUT95), .ZN(n924) );
  NAND2_X1 U888 ( .A1(n830), .A2(n924), .ZN(n826) );
  NAND2_X1 U889 ( .A1(G95), .A2(n881), .ZN(n801) );
  NAND2_X1 U890 ( .A1(G119), .A2(n877), .ZN(n800) );
  NAND2_X1 U891 ( .A1(n801), .A2(n800), .ZN(n805) );
  NAND2_X1 U892 ( .A1(G131), .A2(n516), .ZN(n803) );
  NAND2_X1 U893 ( .A1(G107), .A2(n878), .ZN(n802) );
  NAND2_X1 U894 ( .A1(n803), .A2(n802), .ZN(n804) );
  NOR2_X1 U895 ( .A1(n805), .A2(n804), .ZN(n806) );
  XOR2_X1 U896 ( .A(KEYINPUT96), .B(n806), .Z(n898) );
  AND2_X1 U897 ( .A1(G1991), .A2(n898), .ZN(n817) );
  NAND2_X1 U898 ( .A1(G141), .A2(n516), .ZN(n807) );
  XNOR2_X1 U899 ( .A(n807), .B(KEYINPUT98), .ZN(n815) );
  NAND2_X1 U900 ( .A1(n881), .A2(G105), .ZN(n808) );
  XNOR2_X1 U901 ( .A(n808), .B(KEYINPUT38), .ZN(n810) );
  NAND2_X1 U902 ( .A1(G117), .A2(n878), .ZN(n809) );
  NAND2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n813) );
  NAND2_X1 U904 ( .A1(G129), .A2(n877), .ZN(n811) );
  XNOR2_X1 U905 ( .A(KEYINPUT97), .B(n811), .ZN(n812) );
  NOR2_X1 U906 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U907 ( .A1(n815), .A2(n814), .ZN(n891) );
  AND2_X1 U908 ( .A1(n891), .A2(G1996), .ZN(n816) );
  NOR2_X1 U909 ( .A1(n817), .A2(n816), .ZN(n920) );
  INV_X1 U910 ( .A(n830), .ZN(n818) );
  NOR2_X1 U911 ( .A1(n920), .A2(n818), .ZN(n823) );
  INV_X1 U912 ( .A(n823), .ZN(n819) );
  XNOR2_X1 U913 ( .A(G1986), .B(G290), .ZN(n987) );
  NAND2_X1 U914 ( .A1(n987), .A2(n830), .ZN(n820) );
  NOR2_X1 U915 ( .A1(G1996), .A2(n891), .ZN(n928) );
  NOR2_X1 U916 ( .A1(G1986), .A2(G290), .ZN(n821) );
  NOR2_X1 U917 ( .A1(G1991), .A2(n898), .ZN(n922) );
  NOR2_X1 U918 ( .A1(n821), .A2(n922), .ZN(n822) );
  NOR2_X1 U919 ( .A1(n823), .A2(n822), .ZN(n824) );
  NOR2_X1 U920 ( .A1(n928), .A2(n824), .ZN(n825) );
  XNOR2_X1 U921 ( .A(n825), .B(KEYINPUT39), .ZN(n827) );
  NAND2_X1 U922 ( .A1(n827), .A2(n826), .ZN(n829) );
  NAND2_X1 U923 ( .A1(n901), .A2(n828), .ZN(n936) );
  NAND2_X1 U924 ( .A1(n829), .A2(n936), .ZN(n831) );
  NAND2_X1 U925 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U926 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U928 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U930 ( .A1(n836), .A2(n835), .ZN(G188) );
  XOR2_X1 U931 ( .A(G69), .B(KEYINPUT104), .Z(G235) );
  INV_X1 U933 ( .A(G120), .ZN(G236) );
  INV_X1 U934 ( .A(G96), .ZN(G221) );
  NOR2_X1 U935 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U936 ( .A(G325), .ZN(G261) );
  INV_X1 U937 ( .A(n839), .ZN(G319) );
  XOR2_X1 U938 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n841) );
  XNOR2_X1 U939 ( .A(KEYINPUT105), .B(G2678), .ZN(n840) );
  XNOR2_X1 U940 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U941 ( .A(KEYINPUT42), .B(G2090), .Z(n843) );
  XNOR2_X1 U942 ( .A(G2067), .B(G2072), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U944 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U945 ( .A(G2096), .B(G2100), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(n849) );
  XOR2_X1 U947 ( .A(G2084), .B(G2078), .Z(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(G227) );
  XOR2_X1 U949 ( .A(G1956), .B(G1961), .Z(n851) );
  XNOR2_X1 U950 ( .A(G1996), .B(G1986), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U952 ( .A(G1976), .B(G1981), .Z(n853) );
  XNOR2_X1 U953 ( .A(G1966), .B(G1971), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U955 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U956 ( .A(KEYINPUT41), .B(G2474), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U958 ( .A(KEYINPUT107), .B(n858), .ZN(n859) );
  XOR2_X1 U959 ( .A(n859), .B(G1991), .Z(G229) );
  NAND2_X1 U960 ( .A1(G124), .A2(n877), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n860), .B(KEYINPUT44), .ZN(n863) );
  NAND2_X1 U962 ( .A1(G100), .A2(n881), .ZN(n861) );
  XOR2_X1 U963 ( .A(KEYINPUT109), .B(n861), .Z(n862) );
  NAND2_X1 U964 ( .A1(n863), .A2(n862), .ZN(n868) );
  NAND2_X1 U965 ( .A1(n516), .A2(G136), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n864), .B(KEYINPUT108), .ZN(n866) );
  NAND2_X1 U967 ( .A1(G112), .A2(n878), .ZN(n865) );
  NAND2_X1 U968 ( .A1(n866), .A2(n865), .ZN(n867) );
  NOR2_X1 U969 ( .A1(n868), .A2(n867), .ZN(G162) );
  NAND2_X1 U970 ( .A1(G103), .A2(n881), .ZN(n870) );
  NAND2_X1 U971 ( .A1(G139), .A2(n516), .ZN(n869) );
  NAND2_X1 U972 ( .A1(n870), .A2(n869), .ZN(n875) );
  NAND2_X1 U973 ( .A1(G127), .A2(n877), .ZN(n872) );
  NAND2_X1 U974 ( .A1(G115), .A2(n878), .ZN(n871) );
  NAND2_X1 U975 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U976 ( .A(KEYINPUT47), .B(n873), .Z(n874) );
  NOR2_X1 U977 ( .A1(n875), .A2(n874), .ZN(n915) );
  XOR2_X1 U978 ( .A(n915), .B(G162), .Z(n876) );
  XNOR2_X1 U979 ( .A(n919), .B(n876), .ZN(n890) );
  NAND2_X1 U980 ( .A1(G130), .A2(n877), .ZN(n880) );
  NAND2_X1 U981 ( .A1(G118), .A2(n878), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n888) );
  NAND2_X1 U983 ( .A1(G106), .A2(n881), .ZN(n884) );
  NAND2_X1 U984 ( .A1(G142), .A2(n516), .ZN(n883) );
  NAND2_X1 U985 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U986 ( .A(KEYINPUT45), .B(n885), .Z(n886) );
  XNOR2_X1 U987 ( .A(KEYINPUT110), .B(n886), .ZN(n887) );
  NOR2_X1 U988 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U989 ( .A(n890), .B(n889), .Z(n893) );
  XOR2_X1 U990 ( .A(G160), .B(n891), .Z(n892) );
  XNOR2_X1 U991 ( .A(n893), .B(n892), .ZN(n897) );
  XOR2_X1 U992 ( .A(KEYINPUT46), .B(KEYINPUT111), .Z(n895) );
  XNOR2_X1 U993 ( .A(KEYINPUT112), .B(KEYINPUT48), .ZN(n894) );
  XNOR2_X1 U994 ( .A(n895), .B(n894), .ZN(n896) );
  XOR2_X1 U995 ( .A(n897), .B(n896), .Z(n900) );
  XNOR2_X1 U996 ( .A(G164), .B(n898), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n902) );
  XOR2_X1 U998 ( .A(n902), .B(n901), .Z(n903) );
  NOR2_X1 U999 ( .A1(G37), .A2(n903), .ZN(G395) );
  XOR2_X1 U1000 ( .A(n904), .B(G286), .Z(n906) );
  XNOR2_X1 U1001 ( .A(G171), .B(n975), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1003 ( .A(n907), .B(n980), .Z(n908) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n908), .ZN(G397) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n909) );
  XOR2_X1 U1006 ( .A(KEYINPUT49), .B(n909), .Z(n910) );
  NAND2_X1 U1007 ( .A1(G319), .A2(n910), .ZN(n911) );
  NOR2_X1 U1008 ( .A1(G401), .A2(n911), .ZN(n914) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n912) );
  XOR2_X1 U1010 ( .A(KEYINPUT113), .B(n912), .Z(n913) );
  NAND2_X1 U1011 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G108), .ZN(G238) );
  INV_X1 U1014 ( .A(KEYINPUT55), .ZN(n962) );
  XOR2_X1 U1015 ( .A(KEYINPUT116), .B(KEYINPUT52), .Z(n939) );
  XOR2_X1 U1016 ( .A(G2072), .B(n915), .Z(n917) );
  XOR2_X1 U1017 ( .A(G164), .B(G2078), .Z(n916) );
  NOR2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n918) );
  XOR2_X1 U1019 ( .A(KEYINPUT50), .B(n918), .Z(n935) );
  NAND2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n926) );
  XOR2_X1 U1022 ( .A(G160), .B(G2084), .Z(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n932) );
  XOR2_X1 U1025 ( .A(G2090), .B(G162), .Z(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1027 ( .A(KEYINPUT114), .B(n929), .Z(n930) );
  XOR2_X1 U1028 ( .A(KEYINPUT51), .B(n930), .Z(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1030 ( .A(KEYINPUT115), .B(n933), .ZN(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n937) );
  NAND2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1033 ( .A(n939), .B(n938), .ZN(n940) );
  NAND2_X1 U1034 ( .A1(n962), .A2(n940), .ZN(n941) );
  NAND2_X1 U1035 ( .A1(n941), .A2(G29), .ZN(n1025) );
  XNOR2_X1 U1036 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n942) );
  XNOR2_X1 U1037 ( .A(n942), .B(G34), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(G2084), .B(n943), .ZN(n960) );
  XNOR2_X1 U1039 ( .A(G2090), .B(G35), .ZN(n958) );
  XOR2_X1 U1040 ( .A(G25), .B(G1991), .Z(n944) );
  NAND2_X1 U1041 ( .A1(n944), .A2(G28), .ZN(n955) );
  XNOR2_X1 U1042 ( .A(G27), .B(KEYINPUT117), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(n946), .B(n945), .ZN(n948) );
  XNOR2_X1 U1044 ( .A(G32), .B(G1996), .ZN(n947) );
  NOR2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1046 ( .A(KEYINPUT118), .B(n949), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(G2067), .B(G26), .ZN(n951) );
  XNOR2_X1 U1048 ( .A(G33), .B(G2072), .ZN(n950) );
  NOR2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(KEYINPUT53), .B(n956), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(n962), .B(n961), .ZN(n964) );
  INV_X1 U1056 ( .A(G29), .ZN(n963) );
  NAND2_X1 U1057 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1058 ( .A1(G11), .A2(n965), .ZN(n1023) );
  XNOR2_X1 U1059 ( .A(G16), .B(KEYINPUT56), .ZN(n992) );
  XNOR2_X1 U1060 ( .A(G1966), .B(G168), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(n966), .B(KEYINPUT120), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(n969), .B(KEYINPUT57), .ZN(n979) );
  NAND2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n973) );
  AND2_X1 U1065 ( .A1(G303), .A2(G1971), .ZN(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(n974), .B(KEYINPUT121), .ZN(n977) );
  XNOR2_X1 U1068 ( .A(n975), .B(G1348), .ZN(n976) );
  NOR2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n982) );
  XNOR2_X1 U1071 ( .A(G1341), .B(n980), .ZN(n981) );
  NOR2_X1 U1072 ( .A1(n982), .A2(n981), .ZN(n989) );
  XNOR2_X1 U1073 ( .A(n983), .B(G1956), .ZN(n985) );
  XNOR2_X1 U1074 ( .A(G171), .B(G1961), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1078 ( .A(KEYINPUT122), .B(n990), .ZN(n991) );
  NAND2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n1021) );
  INV_X1 U1080 ( .A(G16), .ZN(n1019) );
  XOR2_X1 U1081 ( .A(G1976), .B(G23), .Z(n994) );
  XOR2_X1 U1082 ( .A(G1971), .B(G22), .Z(n993) );
  NAND2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n996) );
  XNOR2_X1 U1084 ( .A(G24), .B(G1986), .ZN(n995) );
  NOR2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1086 ( .A(KEYINPUT58), .B(n997), .Z(n1015) );
  XOR2_X1 U1087 ( .A(G1341), .B(G19), .Z(n1000) );
  XNOR2_X1 U1088 ( .A(n998), .B(G20), .ZN(n999) );
  NAND2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1006) );
  XOR2_X1 U1090 ( .A(G1981), .B(G6), .Z(n1004) );
  XOR2_X1 U1091 ( .A(G1348), .B(G4), .Z(n1001) );
  XNOR2_X1 U1092 ( .A(KEYINPUT123), .B(n1001), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(n1002), .B(KEYINPUT59), .ZN(n1003) );
  NAND2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(KEYINPUT60), .B(n1007), .ZN(n1009) );
  XOR2_X1 U1097 ( .A(G1961), .B(G5), .Z(n1008) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(G21), .B(G1966), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(KEYINPUT124), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(KEYINPUT125), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1104 ( .A(n1016), .B(KEYINPUT61), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(n1017), .B(KEYINPUT126), .ZN(n1018) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1026), .Z(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

