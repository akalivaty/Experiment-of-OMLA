//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 0 1 0 0 1 1 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986;
  INV_X1    g000(.A(KEYINPUT15), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G478), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT89), .ZN(new_n189));
  XOR2_X1   g003(.A(KEYINPUT9), .B(G234), .Z(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(G217), .A3(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT87), .ZN(new_n194));
  INV_X1    g008(.A(G122), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G116), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT14), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n194), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(G116), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n196), .A2(new_n197), .ZN(new_n200));
  OAI211_X1 g014(.A(KEYINPUT87), .B(KEYINPUT14), .C1(new_n195), .C2(G116), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n198), .A2(new_n199), .A3(new_n200), .A4(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G107), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT88), .ZN(new_n204));
  INV_X1    g018(.A(new_n196), .ZN(new_n205));
  AND2_X1   g019(.A1(new_n205), .A2(new_n199), .ZN(new_n206));
  INV_X1    g020(.A(G107), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(G128), .B(G143), .ZN(new_n209));
  INV_X1    g023(.A(G134), .ZN(new_n210));
  XNOR2_X1  g024(.A(new_n209), .B(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT88), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n202), .A2(new_n212), .A3(G107), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n204), .A2(new_n208), .A3(new_n211), .A4(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n206), .B(new_n207), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n209), .A2(new_n210), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n210), .B1(new_n209), .B2(KEYINPUT13), .ZN(new_n217));
  INV_X1    g031(.A(G143), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G128), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n217), .B1(KEYINPUT13), .B2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n215), .A2(new_n216), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n193), .B1(new_n214), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n214), .A2(new_n221), .A3(new_n193), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G902), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n189), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n224), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n189), .B(new_n226), .C1(new_n228), .C2(new_n222), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n188), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n229), .A2(new_n187), .A3(G478), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(G214), .B1(G237), .B2(G902), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  XOR2_X1   g049(.A(G110), .B(G122), .Z(new_n236));
  INV_X1    g050(.A(G104), .ZN(new_n237));
  NOR3_X1   g051(.A1(new_n237), .A2(KEYINPUT3), .A3(G107), .ZN(new_n238));
  OR2_X1    g052(.A1(KEYINPUT75), .A2(G104), .ZN(new_n239));
  NAND2_X1  g053(.A1(KEYINPUT75), .A2(G104), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n238), .B1(new_n241), .B2(G107), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(new_n207), .A3(new_n240), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT76), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n243), .A2(new_n244), .A3(KEYINPUT3), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n244), .B1(new_n243), .B2(KEYINPUT3), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n242), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G101), .ZN(new_n248));
  INV_X1    g062(.A(G101), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n249), .B(new_n242), .C1(new_n245), .C2(new_n246), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n248), .A2(KEYINPUT4), .A3(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(G116), .B(G119), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT2), .B(G113), .ZN(new_n254));
  OR2_X1    g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n254), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n247), .A2(new_n258), .A3(G101), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n251), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n261));
  INV_X1    g075(.A(G119), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(new_n262), .A3(G116), .ZN(new_n263));
  OAI211_X1 g077(.A(G113), .B(new_n263), .C1(new_n253), .C2(new_n261), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n255), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n243), .B1(G104), .B2(new_n207), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G101), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n250), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT79), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT79), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n250), .A2(new_n270), .A3(new_n267), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n265), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n236), .B1(new_n260), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n251), .A2(new_n257), .A3(new_n259), .ZN(new_n274));
  INV_X1    g088(.A(new_n236), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n250), .A2(new_n270), .A3(new_n267), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n270), .B1(new_n250), .B2(new_n267), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n274), .B(new_n275), .C1(new_n278), .C2(new_n265), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n273), .A2(KEYINPUT6), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n281), .B(new_n236), .C1(new_n260), .C2(new_n272), .ZN(new_n282));
  XNOR2_X1  g096(.A(G143), .B(G146), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(KEYINPUT0), .A3(G128), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT0), .B(G128), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n284), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G125), .ZN(new_n287));
  INV_X1    g101(.A(G128), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n218), .B(G146), .C1(new_n288), .C2(KEYINPUT1), .ZN(new_n289));
  INV_X1    g103(.A(G146), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(new_n290), .A3(G143), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT1), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n283), .A2(new_n294), .A3(G128), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n287), .B1(G125), .B2(new_n296), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n191), .A2(G224), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n297), .B(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n280), .A2(new_n282), .A3(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n265), .B1(KEYINPUT79), .B2(KEYINPUT81), .ZN(new_n301));
  OR2_X1    g115(.A1(new_n301), .A2(new_n268), .ZN(new_n302));
  XOR2_X1   g116(.A(new_n236), .B(KEYINPUT8), .Z(new_n303));
  INV_X1    g117(.A(KEYINPUT81), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n278), .A2(new_n304), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n302), .B(new_n303), .C1(new_n305), .C2(new_n265), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT7), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n298), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n297), .B(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n306), .A2(new_n279), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n300), .A2(new_n226), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(G210), .B1(G237), .B2(G902), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n300), .A2(new_n226), .A3(new_n312), .A4(new_n310), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n235), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G952), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n317), .A2(KEYINPUT90), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(KEYINPUT90), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n191), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n320), .B1(G234), .B2(G237), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  XOR2_X1   g136(.A(KEYINPUT21), .B(G898), .Z(new_n323));
  XNOR2_X1  g137(.A(new_n323), .B(KEYINPUT91), .ZN(new_n324));
  AOI211_X1 g138(.A(new_n226), .B(new_n191), .C1(G234), .C2(G237), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n322), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G475), .ZN(new_n328));
  XNOR2_X1  g142(.A(G113), .B(G122), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT85), .B(G104), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n329), .B(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G237), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(new_n191), .A3(G214), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n218), .ZN(new_n335));
  NOR2_X1   g149(.A1(G237), .A2(G953), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(G143), .A3(G214), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(KEYINPUT18), .A2(G131), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  AND2_X1   g155(.A1(G125), .A2(G140), .ZN(new_n342));
  NOR2_X1   g156(.A1(G125), .A2(G140), .ZN(new_n343));
  OR2_X1    g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(new_n290), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT83), .ZN(new_n346));
  INV_X1    g160(.A(new_n337), .ZN(new_n347));
  AOI21_X1  g161(.A(G143), .B1(new_n336), .B2(G214), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n346), .B1(new_n349), .B2(new_n339), .ZN(new_n350));
  NOR3_X1   g164(.A1(new_n338), .A2(KEYINPUT83), .A3(new_n340), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n341), .B(new_n345), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT84), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n349), .A2(new_n346), .A3(new_n339), .ZN(new_n354));
  OAI21_X1  g168(.A(KEYINPUT83), .B1(new_n338), .B2(new_n340), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT84), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n356), .A2(new_n357), .A3(new_n341), .A4(new_n345), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT16), .B1(new_n342), .B2(new_n343), .ZN(new_n360));
  INV_X1    g174(.A(G125), .ZN(new_n361));
  OR3_X1    g175(.A1(new_n361), .A2(KEYINPUT16), .A3(G140), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n360), .A2(new_n362), .A3(G146), .ZN(new_n363));
  XOR2_X1   g177(.A(new_n344), .B(KEYINPUT19), .Z(new_n364));
  OAI21_X1  g178(.A(new_n363), .B1(new_n364), .B2(G146), .ZN(new_n365));
  OAI21_X1  g179(.A(G131), .B1(new_n347), .B2(new_n348), .ZN(new_n366));
  INV_X1    g180(.A(G131), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n335), .A2(new_n367), .A3(new_n337), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  OR2_X1    g183(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n332), .B1(new_n359), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n331), .B(KEYINPUT86), .ZN(new_n372));
  INV_X1    g186(.A(new_n363), .ZN(new_n373));
  AOI21_X1  g187(.A(G146), .B1(new_n360), .B2(new_n362), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT17), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n366), .A2(new_n376), .A3(new_n368), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n338), .A2(KEYINPUT17), .A3(G131), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n375), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  AOI211_X1 g193(.A(new_n372), .B(new_n379), .C1(new_n353), .C2(new_n358), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n328), .B(new_n226), .C1(new_n371), .C2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT82), .B(KEYINPUT20), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n379), .ZN(new_n384));
  INV_X1    g198(.A(new_n372), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n359), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n365), .A2(new_n369), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n387), .B1(new_n353), .B2(new_n358), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n386), .B1(new_n388), .B2(new_n332), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT20), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n389), .A2(new_n390), .A3(new_n328), .A4(new_n226), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n379), .B1(new_n353), .B2(new_n358), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n392), .A2(new_n332), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n226), .B1(new_n393), .B2(new_n380), .ZN(new_n394));
  AOI22_X1  g208(.A1(new_n383), .A2(new_n391), .B1(G475), .B2(new_n394), .ZN(new_n395));
  AND4_X1   g209(.A1(new_n233), .A2(new_n316), .A3(new_n327), .A4(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(KEYINPUT22), .B(G137), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n398));
  XOR2_X1   g212(.A(new_n397), .B(new_n398), .Z(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n262), .A2(G128), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n401), .B1(KEYINPUT69), .B2(KEYINPUT23), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT23), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n403), .B1(new_n262), .B2(G128), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT69), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n405), .B1(new_n262), .B2(G128), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n402), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(G119), .B(G128), .ZN(new_n408));
  XOR2_X1   g222(.A(KEYINPUT24), .B(G110), .Z(new_n409));
  OAI22_X1  g223(.A1(new_n407), .A2(G110), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n344), .A2(new_n290), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n363), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT70), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n407), .A2(G110), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n409), .A2(new_n408), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n414), .B(new_n415), .C1(new_n373), .C2(new_n374), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n412), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n413), .B1(new_n412), .B2(new_n416), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n400), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n412), .A2(new_n416), .A3(new_n399), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(new_n226), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT25), .ZN(new_n422));
  INV_X1    g236(.A(G217), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n423), .B1(G234), .B2(new_n226), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT25), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n419), .A2(new_n425), .A3(new_n226), .A4(new_n420), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n422), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT71), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n424), .A2(G902), .ZN(new_n430));
  XOR2_X1   g244(.A(KEYINPUT72), .B(KEYINPUT73), .Z(new_n431));
  XNOR2_X1  g245(.A(new_n430), .B(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n419), .A2(new_n420), .A3(new_n432), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n433), .B(KEYINPUT74), .Z(new_n434));
  NAND4_X1  g248(.A1(new_n422), .A2(KEYINPUT71), .A3(new_n424), .A4(new_n426), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n429), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT32), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT31), .ZN(new_n438));
  INV_X1    g252(.A(new_n286), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT64), .ZN(new_n440));
  INV_X1    g254(.A(G137), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n440), .B1(new_n441), .B2(G134), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n210), .A2(KEYINPUT64), .A3(G137), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n441), .A2(G134), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT11), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n441), .A2(KEYINPUT11), .A3(G134), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n444), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n449), .A2(G131), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n444), .A2(new_n367), .A3(new_n447), .A4(new_n448), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n439), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n257), .ZN(new_n454));
  INV_X1    g268(.A(new_n445), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n441), .A2(G134), .ZN(new_n456));
  OAI21_X1  g270(.A(G131), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n296), .A2(new_n451), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n453), .A2(new_n454), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n451), .A2(new_n457), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT65), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n451), .A2(KEYINPUT65), .A3(new_n457), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n296), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT30), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n466), .A3(new_n453), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n449), .A2(G131), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n286), .B1(new_n468), .B2(new_n451), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n296), .A2(new_n451), .A3(new_n457), .ZN(new_n470));
  OAI21_X1  g284(.A(KEYINPUT30), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n460), .B1(new_n472), .B2(new_n257), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n336), .A2(G210), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n474), .B(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT26), .B(G101), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n476), .B(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n438), .B1(new_n473), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n454), .B1(new_n467), .B2(new_n471), .ZN(new_n480));
  INV_X1    g294(.A(new_n478), .ZN(new_n481));
  NOR4_X1   g295(.A1(new_n480), .A2(KEYINPUT31), .A3(new_n460), .A4(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n469), .A2(new_n470), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT28), .B1(new_n483), .B2(new_n454), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT28), .ZN(new_n485));
  NOR4_X1   g299(.A1(new_n469), .A2(new_n470), .A3(new_n485), .A4(new_n257), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n465), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n257), .B1(new_n488), .B2(new_n469), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n478), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n479), .A2(new_n482), .A3(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(G472), .A2(G902), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n437), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n472), .A2(new_n257), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(new_n459), .A3(new_n478), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT31), .ZN(new_n497));
  INV_X1    g311(.A(new_n490), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n473), .A2(new_n438), .A3(new_n478), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(KEYINPUT32), .A3(new_n492), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n494), .A2(KEYINPUT68), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT68), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n500), .A2(new_n503), .A3(KEYINPUT32), .A4(new_n492), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n459), .A2(new_n485), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n483), .A2(KEYINPUT28), .A3(new_n454), .ZN(new_n507));
  AND4_X1   g321(.A1(new_n489), .A2(new_n506), .A3(new_n507), .A4(new_n478), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n481), .B1(new_n480), .B2(new_n460), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n508), .B1(KEYINPUT67), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n489), .A2(new_n506), .A3(new_n507), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT67), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n511), .A2(new_n512), .A3(new_n481), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n510), .A2(KEYINPUT29), .A3(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n257), .B1(new_n469), .B2(new_n470), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n506), .A2(new_n507), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n478), .A2(KEYINPUT29), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n226), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(G472), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n436), .B1(new_n505), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(G221), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n521), .B1(new_n190), .B2(new_n226), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n296), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n293), .A2(KEYINPUT77), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT77), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n292), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(new_n295), .A3(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT78), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n250), .A2(new_n528), .A3(new_n529), .A4(new_n267), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n250), .A2(new_n267), .A3(new_n528), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT78), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n278), .A2(new_n524), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n450), .A2(new_n452), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT12), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n532), .A2(new_n530), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT10), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n251), .A2(new_n439), .A3(new_n259), .ZN(new_n539));
  OAI211_X1 g353(.A(KEYINPUT10), .B(new_n296), .C1(new_n276), .C2(new_n277), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n538), .A2(new_n534), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n269), .A2(new_n524), .A3(new_n271), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT12), .ZN(new_n544));
  INV_X1    g358(.A(new_n534), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n535), .A2(new_n541), .A3(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(G110), .B(G140), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n191), .A2(G227), .ZN(new_n549));
  XOR2_X1   g363(.A(new_n548), .B(new_n549), .Z(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n545), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n554), .A2(new_n541), .A3(new_n550), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n226), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT80), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n557), .A2(new_n558), .A3(G469), .ZN(new_n559));
  AOI21_X1  g373(.A(G902), .B1(new_n552), .B2(new_n555), .ZN(new_n560));
  INV_X1    g374(.A(G469), .ZN(new_n561));
  OAI21_X1  g375(.A(KEYINPUT80), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n535), .A2(new_n546), .A3(new_n541), .A4(new_n550), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n550), .B1(new_n554), .B2(new_n541), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n561), .B(new_n226), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n559), .A2(new_n562), .A3(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n396), .A2(new_n520), .A3(new_n523), .A4(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT92), .B(G101), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n568), .B(new_n569), .ZN(G3));
  INV_X1    g384(.A(new_n436), .ZN(new_n571));
  OAI21_X1  g385(.A(G472), .B1(new_n491), .B2(G902), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n500), .A2(new_n492), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n567), .A2(new_n571), .A3(new_n523), .A4(new_n574), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n316), .A2(new_n327), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n383), .A2(new_n391), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n394), .A2(G475), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n225), .A2(KEYINPUT33), .ZN(new_n580));
  OR3_X1    g394(.A1(new_n228), .A2(new_n222), .A3(KEYINPUT33), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(new_n581), .A3(G478), .ZN(new_n582));
  INV_X1    g396(.A(G478), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n225), .A2(new_n583), .A3(new_n226), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n583), .A2(new_n226), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n582), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n579), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(KEYINPUT93), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n576), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n575), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(new_n237), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT94), .B(KEYINPUT34), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(G6));
  NAND2_X1  g408(.A1(new_n314), .A2(new_n315), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n231), .A2(new_n232), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT95), .ZN(new_n597));
  INV_X1    g411(.A(new_n382), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n389), .A2(new_n328), .A3(new_n226), .A4(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n383), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  OR3_X1    g414(.A1(new_n381), .A2(new_n597), .A3(new_n382), .ZN(new_n601));
  AND4_X1   g415(.A1(new_n596), .A2(new_n600), .A3(new_n601), .A4(new_n578), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n595), .A2(new_n602), .A3(new_n327), .A4(new_n234), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(KEYINPUT96), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n604), .A2(new_n575), .ZN(new_n605));
  XNOR2_X1  g419(.A(KEYINPUT35), .B(G107), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G9));
  NOR2_X1   g421(.A1(new_n417), .A2(new_n418), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n400), .A2(KEYINPUT36), .ZN(new_n609));
  XOR2_X1   g423(.A(new_n608), .B(new_n609), .Z(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n432), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n429), .A2(new_n435), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(new_n572), .A3(new_n573), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT97), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n612), .A2(new_n572), .A3(KEYINPUT97), .A4(new_n573), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n396), .A2(new_n523), .A3(new_n617), .A4(new_n567), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G110), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT98), .B(KEYINPUT37), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G12));
  AND2_X1   g435(.A1(new_n567), .A2(new_n523), .ZN(new_n622));
  INV_X1    g436(.A(G900), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n321), .B1(new_n623), .B2(new_n325), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n602), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n612), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n505), .B2(new_n519), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n622), .A2(new_n316), .A3(new_n627), .A4(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G128), .ZN(G30));
  XOR2_X1   g445(.A(new_n624), .B(KEYINPUT39), .Z(new_n632));
  NAND2_X1  g446(.A1(new_n622), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(KEYINPUT40), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n460), .A2(new_n478), .ZN(new_n635));
  AOI21_X1  g449(.A(G902), .B1(new_n635), .B2(new_n515), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n478), .B1(new_n480), .B2(new_n460), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI22_X1  g452(.A1(new_n502), .A2(new_n504), .B1(G472), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n579), .A2(new_n596), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT40), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n622), .A2(new_n642), .A3(new_n632), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n595), .B(new_n644), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n645), .A2(new_n235), .A3(new_n612), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n634), .A2(new_n641), .A3(new_n643), .A4(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT100), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT101), .B(G143), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G45));
  INV_X1    g464(.A(KEYINPUT103), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n579), .A2(new_n587), .A3(new_n625), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT102), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n316), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n654), .B1(new_n316), .B2(new_n653), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n629), .A2(new_n523), .A3(new_n567), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n651), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n595), .A2(new_n234), .ZN(new_n661));
  OAI21_X1  g475(.A(KEYINPUT102), .B1(new_n661), .B2(new_n652), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n655), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n663), .A2(new_n622), .A3(KEYINPUT103), .A4(new_n629), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G146), .ZN(G48));
  OAI21_X1  g480(.A(new_n226), .B1(new_n564), .B2(new_n565), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT104), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI211_X1 g483(.A(KEYINPUT104), .B(new_n226), .C1(new_n564), .C2(new_n565), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n669), .A2(G469), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n566), .A2(KEYINPUT105), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n669), .A2(KEYINPUT105), .A3(G469), .A4(new_n670), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n520), .A2(new_n673), .A3(new_n523), .A4(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n590), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT41), .B(G113), .Z(new_n677));
  XOR2_X1   g491(.A(new_n677), .B(KEYINPUT106), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n676), .B(new_n678), .ZN(G15));
  NOR2_X1   g493(.A1(new_n604), .A2(new_n675), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n680), .B(G116), .Z(G18));
  NAND4_X1  g495(.A1(new_n629), .A2(new_n673), .A3(new_n523), .A4(new_n674), .ZN(new_n682));
  INV_X1    g496(.A(new_n396), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n262), .ZN(G21));
  AOI21_X1  g499(.A(KEYINPUT107), .B1(new_n487), .B2(new_n515), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n481), .B1(new_n516), .B2(new_n687), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n497), .B(new_n499), .C1(new_n686), .C2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n492), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT108), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n689), .A2(new_n692), .A3(new_n492), .ZN(new_n693));
  AND4_X1   g507(.A1(new_n571), .A2(new_n691), .A3(new_n572), .A4(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n673), .A2(new_n523), .A3(new_n674), .A4(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n316), .A2(new_n596), .A3(new_n327), .A4(new_n579), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(new_n195), .ZN(G24));
  NAND4_X1  g512(.A1(new_n673), .A2(new_n523), .A3(new_n316), .A4(new_n674), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n691), .A2(new_n693), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n700), .A2(new_n572), .A3(new_n653), .A4(new_n612), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n361), .ZN(G27));
  NAND2_X1  g517(.A1(new_n556), .A2(KEYINPUT109), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT109), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n555), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n704), .A2(G469), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(G469), .A2(G902), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n708), .A2(new_n566), .A3(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n314), .A2(new_n523), .A3(new_n234), .A4(new_n315), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n520), .A2(new_n653), .A3(new_n710), .A4(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT42), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n652), .A2(new_n714), .ZN(new_n717));
  AOI21_X1  g531(.A(KEYINPUT111), .B1(new_n573), .B2(new_n437), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n719));
  AOI211_X1 g533(.A(new_n719), .B(KEYINPUT32), .C1(new_n500), .C2(new_n492), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT110), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n501), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n500), .A2(KEYINPUT110), .A3(KEYINPUT32), .A4(new_n492), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n519), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n571), .B(new_n717), .C1(new_n721), .C2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n710), .A2(new_n712), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n716), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n566), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n706), .B1(KEYINPUT109), .B2(new_n556), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n729), .B1(new_n730), .B2(G469), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n711), .B1(new_n731), .B2(new_n709), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n519), .A2(new_n723), .A3(new_n724), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n718), .A2(new_n720), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n436), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n732), .A2(KEYINPUT112), .A3(new_n735), .A4(new_n717), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n715), .A2(new_n728), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT113), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT113), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n715), .A2(new_n728), .A3(new_n736), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G131), .ZN(G33));
  NAND3_X1  g556(.A1(new_n732), .A2(new_n520), .A3(new_n627), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G134), .ZN(G36));
  NAND2_X1  g558(.A1(new_n730), .A2(KEYINPUT45), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT45), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n556), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n745), .A2(G469), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n709), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT46), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n748), .A2(KEYINPUT46), .A3(new_n709), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(new_n566), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n523), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n595), .A2(new_n235), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n395), .A2(new_n587), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(KEYINPUT43), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n759), .A2(new_n574), .A3(new_n628), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n757), .B1(new_n760), .B2(KEYINPUT44), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n760), .A2(KEYINPUT44), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n755), .A2(new_n632), .A3(new_n761), .A4(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G137), .ZN(G39));
  INV_X1    g578(.A(KEYINPUT47), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n754), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n753), .A2(KEYINPUT47), .A3(new_n523), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n505), .A2(new_n519), .A3(new_n436), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n757), .A2(new_n652), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(KEYINPUT114), .B(G140), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(G42));
  NOR2_X1   g587(.A1(KEYINPUT119), .A2(KEYINPUT51), .ZN(new_n774));
  INV_X1    g588(.A(new_n694), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n759), .A2(new_n322), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT118), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(KEYINPUT118), .B1(new_n759), .B2(new_n322), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n775), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n673), .A2(new_n674), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n781), .A2(new_n523), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n645), .A2(new_n235), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n780), .A2(new_n782), .A3(KEYINPUT50), .A4(new_n783), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n774), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n781), .A2(new_n712), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n639), .A2(new_n571), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n790), .A2(new_n322), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n582), .A2(new_n584), .A3(new_n586), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(new_n395), .A3(new_n793), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n788), .A2(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n781), .A2(new_n522), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n756), .B(new_n780), .C1(new_n768), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n778), .A2(new_n779), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n789), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(new_n572), .A3(new_n612), .A4(new_n700), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n795), .A2(new_n797), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(KEYINPUT119), .A2(KEYINPUT51), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n803), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n795), .A2(new_n797), .A3(new_n805), .A4(new_n801), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n738), .A2(new_n740), .ZN(new_n808));
  OAI22_X1  g622(.A1(new_n675), .A2(new_n590), .B1(new_n695), .B2(new_n696), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n233), .A2(new_n579), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT116), .B1(new_n579), .B2(new_n587), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n812), .B1(new_n813), .B2(new_n810), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n576), .ZN(new_n815));
  OAI22_X1  g629(.A1(new_n682), .A2(new_n683), .B1(new_n575), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n809), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n568), .B(new_n618), .C1(new_n604), .C2(new_n675), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n732), .A2(new_n520), .A3(new_n627), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n595), .A2(new_n235), .A3(new_n624), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n629), .A2(new_n523), .A3(new_n567), .A4(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n596), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n600), .A2(new_n601), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n578), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n820), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n727), .A2(new_n701), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n817), .A2(new_n819), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n808), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n629), .A2(new_n523), .A3(new_n567), .A4(new_n316), .ZN(new_n831));
  OAI22_X1  g645(.A1(new_n831), .A2(new_n626), .B1(new_n699), .B2(new_n701), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n612), .B1(new_n731), .B2(new_n709), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n316), .A2(new_n596), .A3(new_n579), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n835), .A2(new_n639), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n834), .A2(new_n836), .A3(new_n523), .A4(new_n625), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n665), .A2(new_n833), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n630), .B(KEYINPUT117), .C1(new_n699), .C2(new_n701), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n832), .A2(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n837), .A2(KEYINPUT52), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n841), .A2(new_n843), .A3(new_n665), .A4(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n830), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n818), .A2(new_n809), .A3(new_n816), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n622), .A2(new_n233), .A3(new_n629), .A4(new_n821), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n743), .B(new_n828), .C1(new_n850), .C2(new_n825), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n741), .A2(new_n849), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n832), .B1(new_n660), .B2(new_n664), .ZN(new_n854));
  AOI22_X1  g668(.A1(new_n838), .A2(new_n839), .B1(new_n854), .B2(new_n844), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT53), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n848), .A2(new_n856), .A3(KEYINPUT54), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n800), .A2(new_n735), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT48), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n780), .A2(new_n782), .A3(new_n316), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n320), .B1(new_n792), .B2(new_n589), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n847), .B1(new_n853), .B2(new_n855), .ZN(new_n863));
  INV_X1    g677(.A(new_n829), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n737), .A2(KEYINPUT53), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n846), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n863), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n857), .A2(new_n862), .A3(new_n868), .ZN(new_n869));
  OAI22_X1  g683(.A1(new_n807), .A2(new_n869), .B1(G952), .B2(G953), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n781), .B(KEYINPUT49), .ZN(new_n871));
  NOR4_X1   g685(.A1(new_n791), .A2(new_n522), .A3(new_n235), .A4(new_n758), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n645), .A3(new_n872), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n873), .B(KEYINPUT115), .Z(new_n874));
  NAND2_X1  g688(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT120), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n870), .A2(KEYINPUT120), .A3(new_n874), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(G75));
  AOI21_X1  g693(.A(new_n226), .B1(new_n863), .B2(new_n866), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT56), .B1(new_n880), .B2(G210), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n280), .A2(new_n282), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(new_n299), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT55), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n317), .A2(G953), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n881), .A2(new_n884), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(G51));
  XOR2_X1   g702(.A(new_n709), .B(KEYINPUT57), .Z(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n854), .A2(new_n844), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n840), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT53), .B1(new_n830), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n865), .A2(new_n849), .A3(new_n852), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n894), .B1(new_n840), .B2(new_n845), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT54), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n890), .B1(new_n896), .B2(new_n868), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n564), .A2(new_n565), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT121), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n880), .A2(G469), .A3(new_n747), .A4(new_n745), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n863), .A2(new_n866), .A3(new_n867), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n867), .B1(new_n863), .B2(new_n866), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n889), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT121), .ZN(new_n904));
  INV_X1    g718(.A(new_n898), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n899), .A2(new_n900), .A3(new_n906), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n907), .A2(new_n886), .ZN(G54));
  NAND3_X1  g722(.A1(new_n880), .A2(KEYINPUT58), .A3(G475), .ZN(new_n909));
  INV_X1    g723(.A(new_n389), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n880), .A2(KEYINPUT58), .A3(G475), .A4(new_n389), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n911), .A2(new_n886), .A3(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT122), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n913), .B(new_n914), .ZN(G60));
  XNOR2_X1  g729(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n586), .B(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n917), .B1(new_n857), .B2(new_n868), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n580), .A2(new_n581), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT123), .Z(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT125), .ZN(new_n923));
  INV_X1    g737(.A(new_n917), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n921), .B(new_n924), .C1(new_n901), .C2(new_n902), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n922), .A2(new_n923), .A3(new_n886), .A4(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n886), .B1(new_n918), .B2(new_n921), .ZN(new_n927));
  INV_X1    g741(.A(new_n925), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT125), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n926), .A2(new_n929), .ZN(G63));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT126), .Z(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT60), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n863), .B2(new_n866), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n419), .A2(new_n420), .ZN(new_n935));
  OR2_X1    g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n934), .A2(new_n610), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n936), .A2(new_n886), .A3(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT61), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(G66));
  AOI21_X1  g754(.A(new_n191), .B1(new_n324), .B2(G224), .ZN(new_n941));
  INV_X1    g755(.A(new_n849), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n941), .B1(new_n942), .B2(new_n191), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n882), .B1(G898), .B2(new_n191), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n943), .B(new_n944), .Z(G69));
  NAND4_X1  g759(.A1(new_n753), .A2(new_n523), .A3(new_n632), .A4(new_n735), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n743), .B1(new_n946), .B2(new_n835), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n841), .A2(new_n843), .A3(new_n665), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n771), .A2(new_n949), .A3(new_n741), .A4(new_n763), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n191), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n191), .A2(G900), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(KEYINPUT127), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n951), .A2(new_n956), .A3(new_n953), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n472), .B(new_n364), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n771), .A2(new_n763), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n520), .A2(new_n814), .ZN(new_n963));
  OR3_X1    g777(.A1(new_n633), .A2(new_n757), .A3(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n648), .A2(new_n948), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n965), .A2(KEYINPUT62), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n648), .A2(new_n948), .A3(new_n967), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n962), .B(new_n964), .C1(new_n966), .C2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n960), .B1(new_n969), .B2(new_n191), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n191), .B1(G227), .B2(G900), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n961), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n959), .B1(new_n955), .B2(new_n957), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n972), .B1(new_n975), .B2(new_n970), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n974), .A2(new_n976), .ZN(G72));
  OR2_X1    g791(.A1(new_n969), .A2(new_n942), .ZN(new_n978));
  NAND2_X1  g792(.A1(G472), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT63), .Z(new_n980));
  AOI21_X1  g794(.A(new_n637), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n980), .B1(new_n950), .B2(new_n942), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n982), .A2(new_n495), .A3(new_n635), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n496), .A2(new_n509), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n848), .A2(new_n856), .A3(new_n980), .A4(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n983), .A2(new_n886), .A3(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n981), .A2(new_n986), .ZN(G57));
endmodule


