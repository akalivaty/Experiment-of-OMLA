

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724;

  AND2_X1 U365 ( .A1(n459), .A2(n537), .ZN(n462) );
  OR2_X1 U366 ( .A1(n530), .A2(n529), .ZN(n641) );
  NOR2_X1 U367 ( .A1(n572), .A2(n565), .ZN(n499) );
  XNOR2_X1 U368 ( .A(n440), .B(n439), .ZN(n353) );
  NAND2_X1 U369 ( .A1(n438), .A2(n374), .ZN(n440) );
  OR2_X1 U370 ( .A1(n626), .A2(G902), .ZN(n417) );
  NAND2_X2 U371 ( .A1(n343), .A2(n701), .ZN(n654) );
  XNOR2_X2 U372 ( .A(n379), .B(KEYINPUT83), .ZN(n343) );
  XNOR2_X2 U373 ( .A(n710), .B(G146), .ZN(n446) );
  INV_X2 U374 ( .A(G953), .ZN(n718) );
  AND2_X4 U375 ( .A1(n594), .A2(n654), .ZN(n624) );
  OR2_X2 U376 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X2 U377 ( .A(n501), .B(KEYINPUT35), .ZN(n570) );
  NOR2_X1 U378 ( .A1(n520), .A2(n722), .ZN(n521) );
  NAND2_X1 U379 ( .A1(n576), .A2(n564), .ZN(n390) );
  OR2_X1 U380 ( .A1(n522), .A2(n566), .ZN(n514) );
  NOR2_X1 U381 ( .A1(n507), .A2(n506), .ZN(n508) );
  XNOR2_X1 U382 ( .A(n449), .B(n448), .ZN(n566) );
  AND2_X1 U383 ( .A1(n380), .A2(n381), .ZN(n717) );
  XNOR2_X1 U384 ( .A(n559), .B(n382), .ZN(n380) );
  NAND2_X1 U385 ( .A1(n354), .A2(n558), .ZN(n559) );
  AND2_X1 U386 ( .A1(n363), .A2(n583), .ZN(n362) );
  XNOR2_X1 U387 ( .A(n356), .B(n355), .ZN(n354) );
  AND2_X1 U388 ( .A1(n549), .A2(n548), .ZN(n357) );
  NOR2_X1 U389 ( .A1(n692), .A2(n517), .ZN(n519) );
  OR2_X1 U390 ( .A1(n541), .A2(n540), .ZN(n640) );
  OR2_X1 U391 ( .A1(n565), .A2(n522), .ZN(n378) );
  OR2_X1 U392 ( .A1(n566), .A2(n678), .ZN(n452) );
  XNOR2_X1 U393 ( .A(n566), .B(n496), .ZN(n565) );
  XNOR2_X1 U394 ( .A(n386), .B(n385), .ZN(n442) );
  XNOR2_X1 U395 ( .A(n424), .B(n423), .ZN(n711) );
  XOR2_X1 U396 ( .A(G125), .B(G146), .Z(n423) );
  XNOR2_X2 U397 ( .A(n484), .B(n409), .ZN(n710) );
  NOR2_X1 U398 ( .A1(n571), .A2(KEYINPUT44), .ZN(n364) );
  NAND2_X1 U399 ( .A1(n493), .A2(n345), .ZN(n391) );
  XNOR2_X1 U400 ( .A(n584), .B(KEYINPUT45), .ZN(n592) );
  NAND2_X1 U401 ( .A1(n362), .A2(n359), .ZN(n584) );
  AND2_X1 U402 ( .A1(n361), .A2(n360), .ZN(n359) );
  INV_X1 U403 ( .A(n560), .ZN(n381) );
  INV_X1 U404 ( .A(n723), .ZN(n558) );
  AND2_X1 U405 ( .A1(n353), .A2(n673), .ZN(n459) );
  XNOR2_X1 U406 ( .A(n499), .B(n498), .ZN(n672) );
  XNOR2_X1 U407 ( .A(n495), .B(KEYINPUT1), .ZN(n377) );
  XNOR2_X1 U408 ( .A(n393), .B(KEYINPUT3), .ZN(n385) );
  XNOR2_X1 U409 ( .A(n388), .B(n387), .ZN(n386) );
  INV_X1 U410 ( .A(KEYINPUT66), .ZN(n393) );
  XNOR2_X1 U411 ( .A(G110), .B(G107), .ZN(n394) );
  XNOR2_X1 U412 ( .A(n700), .B(n366), .ZN(n610) );
  XNOR2_X1 U413 ( .A(n368), .B(n367), .ZN(n366) );
  XNOR2_X1 U414 ( .A(n405), .B(n399), .ZN(n367) );
  XNOR2_X1 U415 ( .A(n401), .B(n400), .ZN(n368) );
  BUF_X1 U416 ( .A(n592), .Z(n701) );
  INV_X1 U417 ( .A(n661), .ZN(n375) );
  INV_X1 U418 ( .A(n565), .ZN(n372) );
  INV_X1 U419 ( .A(KEYINPUT22), .ZN(n389) );
  BUF_X1 U420 ( .A(n377), .Z(n373) );
  NAND2_X1 U421 ( .A1(n542), .A2(n640), .ZN(n543) );
  XNOR2_X1 U422 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n408) );
  INV_X1 U423 ( .A(KEYINPUT48), .ZN(n355) );
  XNOR2_X1 U424 ( .A(G101), .B(G113), .ZN(n387) );
  XNOR2_X1 U425 ( .A(G116), .B(G119), .ZN(n388) );
  XNOR2_X1 U426 ( .A(n350), .B(KEYINPUT71), .ZN(n572) );
  XNOR2_X1 U427 ( .A(G128), .B(G119), .ZN(n425) );
  XNOR2_X1 U428 ( .A(G116), .B(G122), .ZN(n475) );
  XNOR2_X1 U429 ( .A(KEYINPUT105), .B(KEYINPUT104), .ZN(n477) );
  XNOR2_X1 U430 ( .A(n378), .B(KEYINPUT112), .ZN(n523) );
  XNOR2_X1 U431 ( .A(n524), .B(n348), .ZN(n493) );
  INV_X1 U432 ( .A(KEYINPUT115), .ZN(n515) );
  XNOR2_X1 U433 ( .A(n514), .B(KEYINPUT28), .ZN(n516) );
  XNOR2_X1 U434 ( .A(n369), .B(n344), .ZN(n700) );
  XNOR2_X1 U435 ( .A(n442), .B(n384), .ZN(n369) );
  INV_X1 U436 ( .A(KEYINPUT16), .ZN(n384) );
  NAND2_X1 U437 ( .A1(n591), .A2(n590), .ZN(n594) );
  XNOR2_X1 U438 ( .A(n446), .B(n415), .ZN(n626) );
  OR2_X1 U439 ( .A1(n718), .A2(G952), .ZN(n622) );
  NAND2_X1 U440 ( .A1(n351), .A2(n539), .ZN(n501) );
  XNOR2_X1 U441 ( .A(n352), .B(n500), .ZN(n351) );
  XNOR2_X1 U442 ( .A(n370), .B(KEYINPUT32), .ZN(n724) );
  NOR2_X1 U443 ( .A1(n346), .A2(n372), .ZN(n371) );
  AND2_X1 U444 ( .A1(n567), .A2(n565), .ZN(n579) );
  XOR2_X1 U445 ( .A(G122), .B(n414), .Z(n344) );
  OR2_X1 U446 ( .A1(n492), .A2(n491), .ZN(n345) );
  INV_X1 U447 ( .A(n659), .ZN(n374) );
  NAND2_X1 U448 ( .A1(n376), .A2(n375), .ZN(n346) );
  AND2_X1 U449 ( .A1(n381), .A2(KEYINPUT2), .ZN(n347) );
  XNOR2_X1 U450 ( .A(KEYINPUT72), .B(KEYINPUT19), .ZN(n348) );
  XNOR2_X1 U451 ( .A(KEYINPUT86), .B(KEYINPUT46), .ZN(n349) );
  NOR2_X1 U452 ( .A1(n377), .A2(n659), .ZN(n350) );
  XNOR2_X2 U453 ( .A(n417), .B(n416), .ZN(n495) );
  NAND2_X1 U454 ( .A1(n672), .A2(n576), .ZN(n352) );
  NAND2_X1 U455 ( .A1(n537), .A2(n353), .ZN(n541) );
  AND2_X1 U456 ( .A1(n353), .A2(n665), .ZN(n575) );
  NAND2_X1 U457 ( .A1(n358), .A2(n357), .ZN(n356) );
  XNOR2_X1 U458 ( .A(n521), .B(n349), .ZN(n358) );
  INV_X1 U459 ( .A(n377), .ZN(n376) );
  NAND2_X1 U460 ( .A1(n571), .A2(KEYINPUT44), .ZN(n360) );
  NAND2_X1 U461 ( .A1(n570), .A2(KEYINPUT44), .ZN(n361) );
  NAND2_X1 U462 ( .A1(n365), .A2(n364), .ZN(n363) );
  INV_X1 U463 ( .A(n570), .ZN(n365) );
  NAND2_X1 U464 ( .A1(n493), .A2(n438), .ZN(n529) );
  NAND2_X1 U465 ( .A1(n567), .A2(n371), .ZN(n370) );
  XNOR2_X2 U466 ( .A(n390), .B(n389), .ZN(n567) );
  AND2_X1 U467 ( .A1(n373), .A2(n661), .ZN(n580) );
  NAND2_X1 U468 ( .A1(n373), .A2(n659), .ZN(n660) );
  NAND2_X1 U469 ( .A1(n551), .A2(n373), .ZN(n553) );
  NOR2_X1 U470 ( .A1(n528), .A2(n373), .ZN(n650) );
  NAND2_X1 U471 ( .A1(n569), .A2(n373), .ZN(n637) );
  XNOR2_X2 U472 ( .A(n405), .B(G134), .ZN(n484) );
  NAND2_X1 U473 ( .A1(n380), .A2(n347), .ZN(n379) );
  INV_X1 U474 ( .A(KEYINPUT84), .ZN(n382) );
  XNOR2_X2 U475 ( .A(n383), .B(G143), .ZN(n405) );
  XNOR2_X2 U476 ( .A(G128), .B(KEYINPUT64), .ZN(n383) );
  XNOR2_X2 U477 ( .A(n391), .B(n494), .ZN(n576) );
  BUF_X1 U478 ( .A(n566), .Z(n665) );
  XOR2_X1 U479 ( .A(n468), .B(n467), .Z(n392) );
  INV_X1 U480 ( .A(KEYINPUT5), .ZN(n441) );
  XNOR2_X1 U481 ( .A(n442), .B(n441), .ZN(n444) );
  OR2_X1 U482 ( .A1(n678), .A2(n676), .ZN(n509) );
  XNOR2_X1 U483 ( .A(n447), .B(G472), .ZN(n448) );
  XNOR2_X1 U484 ( .A(n472), .B(G475), .ZN(n473) );
  XNOR2_X1 U485 ( .A(n474), .B(n473), .ZN(n506) );
  XNOR2_X1 U486 ( .A(n394), .B(G104), .ZN(n414) );
  XOR2_X1 U487 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n396) );
  XNOR2_X1 U488 ( .A(KEYINPUT74), .B(KEYINPUT91), .ZN(n395) );
  XNOR2_X1 U489 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U490 ( .A(n397), .B(n408), .ZN(n401) );
  INV_X1 U491 ( .A(n423), .ZN(n398) );
  XNOR2_X1 U492 ( .A(KEYINPUT75), .B(n398), .ZN(n400) );
  NAND2_X1 U493 ( .A1(G224), .A2(n718), .ZN(n399) );
  XNOR2_X1 U494 ( .A(G902), .B(KEYINPUT15), .ZN(n585) );
  NAND2_X1 U495 ( .A1(n610), .A2(n585), .ZN(n403) );
  OR2_X1 U496 ( .A1(G902), .A2(G237), .ZN(n450) );
  AND2_X1 U497 ( .A1(G210), .A2(n450), .ZN(n402) );
  XNOR2_X2 U498 ( .A(n403), .B(n402), .ZN(n538) );
  XNOR2_X1 U499 ( .A(KEYINPUT70), .B(KEYINPUT38), .ZN(n404) );
  XNOR2_X1 U500 ( .A(n538), .B(n404), .ZN(n677) );
  INV_X1 U501 ( .A(G137), .ZN(n406) );
  XNOR2_X1 U502 ( .A(n406), .B(G131), .ZN(n407) );
  XNOR2_X1 U503 ( .A(n408), .B(n407), .ZN(n409) );
  NAND2_X1 U504 ( .A1(n718), .A2(G227), .ZN(n410) );
  XNOR2_X1 U505 ( .A(n410), .B(G101), .ZN(n412) );
  XNOR2_X1 U506 ( .A(KEYINPUT73), .B(G140), .ZN(n411) );
  XNOR2_X1 U507 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U508 ( .A(n414), .B(n413), .ZN(n415) );
  INV_X1 U509 ( .A(G469), .ZN(n416) );
  INV_X1 U510 ( .A(n495), .ZN(n438) );
  XOR2_X1 U511 ( .A(KEYINPUT96), .B(KEYINPUT21), .Z(n421) );
  XOR2_X1 U512 ( .A(KEYINPUT95), .B(KEYINPUT20), .Z(n419) );
  NAND2_X1 U513 ( .A1(G234), .A2(n585), .ZN(n418) );
  XNOR2_X1 U514 ( .A(n419), .B(n418), .ZN(n433) );
  NAND2_X1 U515 ( .A1(n433), .A2(G221), .ZN(n420) );
  XNOR2_X1 U516 ( .A(n421), .B(n420), .ZN(n662) );
  INV_X1 U517 ( .A(KEYINPUT97), .ZN(n422) );
  XNOR2_X1 U518 ( .A(n662), .B(n422), .ZN(n562) );
  XNOR2_X1 U519 ( .A(G140), .B(KEYINPUT10), .ZN(n424) );
  XOR2_X1 U520 ( .A(G137), .B(G110), .Z(n426) );
  XNOR2_X1 U521 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U522 ( .A(n711), .B(n427), .ZN(n432) );
  NAND2_X1 U523 ( .A1(G234), .A2(n718), .ZN(n428) );
  XOR2_X1 U524 ( .A(KEYINPUT8), .B(n428), .Z(n481) );
  NAND2_X1 U525 ( .A1(G221), .A2(n481), .ZN(n430) );
  XOR2_X1 U526 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n429) );
  XNOR2_X1 U527 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U528 ( .A(n432), .B(n431), .ZN(n621) );
  INV_X1 U529 ( .A(G902), .ZN(n486) );
  NAND2_X1 U530 ( .A1(n621), .A2(n486), .ZN(n437) );
  XOR2_X1 U531 ( .A(KEYINPUT25), .B(KEYINPUT94), .Z(n435) );
  NAND2_X1 U532 ( .A1(n433), .A2(G217), .ZN(n434) );
  XNOR2_X1 U533 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X2 U534 ( .A(n437), .B(n436), .ZN(n661) );
  NAND2_X1 U535 ( .A1(n562), .A2(n661), .ZN(n659) );
  INV_X1 U536 ( .A(KEYINPUT98), .ZN(n439) );
  NOR2_X1 U537 ( .A1(G953), .A2(G237), .ZN(n463) );
  NAND2_X1 U538 ( .A1(n463), .A2(G210), .ZN(n443) );
  XNOR2_X1 U539 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U540 ( .A(n446), .B(n445), .ZN(n602) );
  NOR2_X1 U541 ( .A1(n602), .A2(G902), .ZN(n449) );
  INV_X1 U542 ( .A(KEYINPUT99), .ZN(n447) );
  NAND2_X1 U543 ( .A1(G214), .A2(n450), .ZN(n674) );
  INV_X1 U544 ( .A(n674), .ZN(n678) );
  INV_X1 U545 ( .A(KEYINPUT30), .ZN(n451) );
  XNOR2_X1 U546 ( .A(n452), .B(n451), .ZN(n458) );
  XOR2_X1 U547 ( .A(KEYINPUT69), .B(KEYINPUT14), .Z(n454) );
  NAND2_X1 U548 ( .A1(G237), .A2(G234), .ZN(n453) );
  XNOR2_X1 U549 ( .A(n454), .B(n453), .ZN(n455) );
  NAND2_X1 U550 ( .A1(G952), .A2(n455), .ZN(n690) );
  NOR2_X1 U551 ( .A1(G953), .A2(n690), .ZN(n492) );
  NAND2_X1 U552 ( .A1(G902), .A2(n455), .ZN(n489) );
  OR2_X1 U553 ( .A1(n718), .A2(n489), .ZN(n456) );
  NOR2_X1 U554 ( .A1(G900), .A2(n456), .ZN(n457) );
  OR2_X1 U555 ( .A1(n492), .A2(n457), .ZN(n511) );
  AND2_X1 U556 ( .A1(n458), .A2(n511), .ZN(n537) );
  XOR2_X1 U557 ( .A(KEYINPUT87), .B(KEYINPUT39), .Z(n460) );
  XNOR2_X1 U558 ( .A(n460), .B(KEYINPUT68), .ZN(n461) );
  XNOR2_X1 U559 ( .A(n462), .B(n461), .ZN(n504) );
  NAND2_X1 U560 ( .A1(G214), .A2(n463), .ZN(n464) );
  XNOR2_X1 U561 ( .A(n711), .B(n464), .ZN(n471) );
  XOR2_X1 U562 ( .A(G113), .B(G131), .Z(n466) );
  XNOR2_X1 U563 ( .A(G122), .B(G104), .ZN(n465) );
  XNOR2_X1 U564 ( .A(n466), .B(n465), .ZN(n469) );
  XOR2_X1 U565 ( .A(KEYINPUT101), .B(KEYINPUT11), .Z(n468) );
  XNOR2_X1 U566 ( .A(G143), .B(KEYINPUT12), .ZN(n467) );
  XNOR2_X1 U567 ( .A(n469), .B(n392), .ZN(n470) );
  XNOR2_X1 U568 ( .A(n471), .B(n470), .ZN(n596) );
  NOR2_X1 U569 ( .A1(G902), .A2(n596), .ZN(n474) );
  XNOR2_X1 U570 ( .A(KEYINPUT102), .B(KEYINPUT13), .ZN(n472) );
  XOR2_X1 U571 ( .A(KEYINPUT103), .B(G107), .Z(n476) );
  XNOR2_X1 U572 ( .A(n476), .B(n475), .ZN(n480) );
  XOR2_X1 U573 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n478) );
  XNOR2_X1 U574 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U575 ( .A(n480), .B(n479), .Z(n483) );
  NAND2_X1 U576 ( .A1(G217), .A2(n481), .ZN(n482) );
  XNOR2_X1 U577 ( .A(n483), .B(n482), .ZN(n485) );
  XNOR2_X1 U578 ( .A(n485), .B(n484), .ZN(n616) );
  NAND2_X1 U579 ( .A1(n616), .A2(n486), .ZN(n487) );
  XNOR2_X1 U580 ( .A(n487), .B(G478), .ZN(n507) );
  INV_X1 U581 ( .A(n507), .ZN(n502) );
  OR2_X1 U582 ( .A1(n506), .A2(n502), .ZN(n646) );
  NOR2_X1 U583 ( .A1(n504), .A2(n646), .ZN(n560) );
  XOR2_X1 U584 ( .A(G134), .B(n560), .Z(G36) );
  NAND2_X1 U585 ( .A1(n538), .A2(n674), .ZN(n524) );
  NOR2_X1 U586 ( .A1(G898), .A2(n718), .ZN(n488) );
  XOR2_X1 U587 ( .A(KEYINPUT92), .B(n488), .Z(n699) );
  NOR2_X1 U588 ( .A1(n699), .A2(n489), .ZN(n490) );
  XOR2_X1 U589 ( .A(KEYINPUT93), .B(n490), .Z(n491) );
  INV_X1 U590 ( .A(KEYINPUT0), .ZN(n494) );
  XNOR2_X1 U591 ( .A(KEYINPUT107), .B(KEYINPUT6), .ZN(n496) );
  XNOR2_X1 U592 ( .A(KEYINPUT110), .B(KEYINPUT33), .ZN(n497) );
  XNOR2_X1 U593 ( .A(n497), .B(KEYINPUT67), .ZN(n498) );
  INV_X1 U594 ( .A(KEYINPUT34), .ZN(n500) );
  AND2_X1 U595 ( .A1(n506), .A2(n507), .ZN(n539) );
  XOR2_X1 U596 ( .A(n570), .B(G122), .Z(G24) );
  NAND2_X1 U597 ( .A1(n506), .A2(n502), .ZN(n503) );
  XNOR2_X1 U598 ( .A(n503), .B(KEYINPUT106), .ZN(n531) );
  NOR2_X1 U599 ( .A1(n504), .A2(n531), .ZN(n505) );
  XNOR2_X1 U600 ( .A(n505), .B(KEYINPUT40), .ZN(n520) );
  XOR2_X1 U601 ( .A(n520), .B(G131), .Z(G33) );
  XOR2_X1 U602 ( .A(n508), .B(KEYINPUT108), .Z(n676) );
  NOR2_X1 U603 ( .A1(n509), .A2(n677), .ZN(n510) );
  XNOR2_X1 U604 ( .A(n510), .B(KEYINPUT41), .ZN(n692) );
  INV_X1 U605 ( .A(n511), .ZN(n512) );
  NOR2_X1 U606 ( .A1(n661), .A2(n512), .ZN(n513) );
  NAND2_X1 U607 ( .A1(n662), .A2(n513), .ZN(n522) );
  XNOR2_X1 U608 ( .A(n516), .B(n515), .ZN(n530) );
  OR2_X1 U609 ( .A1(n530), .A2(n495), .ZN(n517) );
  XNOR2_X1 U610 ( .A(KEYINPUT116), .B(KEYINPUT42), .ZN(n518) );
  XNOR2_X1 U611 ( .A(n519), .B(n518), .ZN(n722) );
  XOR2_X1 U612 ( .A(KEYINPUT111), .B(n531), .Z(n643) );
  NOR2_X1 U613 ( .A1(n643), .A2(n523), .ZN(n550) );
  INV_X1 U614 ( .A(n524), .ZN(n525) );
  AND2_X1 U615 ( .A1(n550), .A2(n525), .ZN(n527) );
  INV_X1 U616 ( .A(KEYINPUT36), .ZN(n526) );
  XNOR2_X1 U617 ( .A(n527), .B(n526), .ZN(n528) );
  AND2_X1 U618 ( .A1(n531), .A2(n646), .ZN(n680) );
  XNOR2_X1 U619 ( .A(n680), .B(KEYINPUT79), .ZN(n577) );
  INV_X1 U620 ( .A(KEYINPUT47), .ZN(n532) );
  NAND2_X1 U621 ( .A1(n577), .A2(n532), .ZN(n533) );
  NOR2_X1 U622 ( .A1(n641), .A2(n533), .ZN(n534) );
  NOR2_X1 U623 ( .A1(n650), .A2(n534), .ZN(n549) );
  INV_X1 U624 ( .A(KEYINPUT77), .ZN(n547) );
  INV_X1 U625 ( .A(KEYINPUT78), .ZN(n536) );
  NAND2_X1 U626 ( .A1(KEYINPUT47), .A2(n641), .ZN(n535) );
  XNOR2_X1 U627 ( .A(n536), .B(n535), .ZN(n545) );
  NAND2_X1 U628 ( .A1(n680), .A2(KEYINPUT47), .ZN(n542) );
  NAND2_X1 U629 ( .A1(n538), .A2(n539), .ZN(n540) );
  XNOR2_X1 U630 ( .A(KEYINPUT76), .B(n543), .ZN(n544) );
  NOR2_X1 U631 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U632 ( .A(n547), .B(n546), .ZN(n548) );
  AND2_X1 U633 ( .A1(n550), .A2(n674), .ZN(n551) );
  XOR2_X1 U634 ( .A(KEYINPUT43), .B(KEYINPUT113), .Z(n552) );
  XNOR2_X1 U635 ( .A(n553), .B(n552), .ZN(n555) );
  INV_X1 U636 ( .A(n538), .ZN(n554) );
  NAND2_X1 U637 ( .A1(n555), .A2(n554), .ZN(n557) );
  INV_X1 U638 ( .A(KEYINPUT114), .ZN(n556) );
  XNOR2_X1 U639 ( .A(n557), .B(n556), .ZN(n723) );
  INV_X1 U640 ( .A(n676), .ZN(n561) );
  NAND2_X1 U641 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U642 ( .A(n563), .B(KEYINPUT109), .ZN(n564) );
  NAND2_X1 U643 ( .A1(n665), .A2(n567), .ZN(n568) );
  NOR2_X1 U644 ( .A1(n661), .A2(n568), .ZN(n569) );
  NAND2_X1 U645 ( .A1(n724), .A2(n637), .ZN(n571) );
  NOR2_X1 U646 ( .A1(n572), .A2(n665), .ZN(n669) );
  NAND2_X1 U647 ( .A1(n576), .A2(n669), .ZN(n574) );
  XOR2_X1 U648 ( .A(KEYINPUT100), .B(KEYINPUT31), .Z(n573) );
  XNOR2_X1 U649 ( .A(n574), .B(n573), .ZN(n647) );
  NAND2_X1 U650 ( .A1(n576), .A2(n575), .ZN(n633) );
  NAND2_X1 U651 ( .A1(n647), .A2(n633), .ZN(n578) );
  AND2_X1 U652 ( .A1(n578), .A2(n577), .ZN(n582) );
  XNOR2_X1 U653 ( .A(n579), .B(KEYINPUT88), .ZN(n581) );
  AND2_X1 U654 ( .A1(n581), .A2(n580), .ZN(n631) );
  NOR2_X1 U655 ( .A1(n582), .A2(n631), .ZN(n583) );
  INV_X1 U656 ( .A(n585), .ZN(n589) );
  NAND2_X1 U657 ( .A1(n592), .A2(n589), .ZN(n587) );
  INV_X1 U658 ( .A(KEYINPUT82), .ZN(n586) );
  XNOR2_X1 U659 ( .A(n587), .B(n586), .ZN(n588) );
  NAND2_X1 U660 ( .A1(n717), .A2(n588), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n589), .A2(KEYINPUT2), .ZN(n590) );
  NAND2_X1 U662 ( .A1(n624), .A2(G475), .ZN(n598) );
  XNOR2_X1 U663 ( .A(KEYINPUT90), .B(KEYINPUT59), .ZN(n595) );
  XNOR2_X1 U664 ( .A(n596), .B(n595), .ZN(n597) );
  XNOR2_X1 U665 ( .A(n598), .B(n597), .ZN(n599) );
  NAND2_X1 U666 ( .A1(n599), .A2(n622), .ZN(n601) );
  INV_X1 U667 ( .A(KEYINPUT60), .ZN(n600) );
  XNOR2_X1 U668 ( .A(n601), .B(n600), .ZN(G60) );
  NAND2_X1 U669 ( .A1(n624), .A2(G472), .ZN(n605) );
  XNOR2_X1 U670 ( .A(KEYINPUT117), .B(KEYINPUT62), .ZN(n603) );
  XNOR2_X1 U671 ( .A(n602), .B(n603), .ZN(n604) );
  XNOR2_X1 U672 ( .A(n605), .B(n604), .ZN(n606) );
  NAND2_X1 U673 ( .A1(n606), .A2(n622), .ZN(n607) );
  XNOR2_X1 U674 ( .A(n607), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U675 ( .A1(n624), .A2(G210), .ZN(n612) );
  XNOR2_X1 U676 ( .A(KEYINPUT89), .B(KEYINPUT54), .ZN(n608) );
  XNOR2_X1 U677 ( .A(n608), .B(KEYINPUT55), .ZN(n609) );
  XNOR2_X1 U678 ( .A(n610), .B(n609), .ZN(n611) );
  XNOR2_X1 U679 ( .A(n612), .B(n611), .ZN(n613) );
  NAND2_X1 U680 ( .A1(n613), .A2(n622), .ZN(n615) );
  XNOR2_X1 U681 ( .A(KEYINPUT85), .B(KEYINPUT56), .ZN(n614) );
  XNOR2_X1 U682 ( .A(n615), .B(n614), .ZN(G51) );
  NAND2_X1 U683 ( .A1(n624), .A2(G478), .ZN(n617) );
  XNOR2_X1 U684 ( .A(n617), .B(n616), .ZN(n618) );
  NAND2_X1 U685 ( .A1(n618), .A2(n622), .ZN(n619) );
  XNOR2_X1 U686 ( .A(n619), .B(KEYINPUT123), .ZN(G63) );
  AND2_X1 U687 ( .A1(n624), .A2(G217), .ZN(n620) );
  XNOR2_X1 U688 ( .A(n621), .B(n620), .ZN(n623) );
  INV_X1 U689 ( .A(n622), .ZN(n629) );
  NOR2_X1 U690 ( .A1(n623), .A2(n629), .ZN(G66) );
  NAND2_X1 U691 ( .A1(n624), .A2(G469), .ZN(n628) );
  XOR2_X1 U692 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n625) );
  XNOR2_X1 U693 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X1 U694 ( .A(n628), .B(n627), .ZN(n630) );
  NOR2_X1 U695 ( .A1(n630), .A2(n629), .ZN(G54) );
  XOR2_X1 U696 ( .A(G101), .B(n631), .Z(G3) );
  NOR2_X1 U697 ( .A1(n643), .A2(n633), .ZN(n632) );
  XOR2_X1 U698 ( .A(G104), .B(n632), .Z(G6) );
  NOR2_X1 U699 ( .A1(n646), .A2(n633), .ZN(n635) );
  XNOR2_X1 U700 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n634) );
  XNOR2_X1 U701 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U702 ( .A(G107), .B(n636), .ZN(G9) );
  XNOR2_X1 U703 ( .A(G110), .B(n637), .ZN(G12) );
  XOR2_X1 U704 ( .A(G128), .B(KEYINPUT29), .Z(n639) );
  OR2_X1 U705 ( .A1(n641), .A2(n646), .ZN(n638) );
  XNOR2_X1 U706 ( .A(n639), .B(n638), .ZN(G30) );
  XNOR2_X1 U707 ( .A(G143), .B(n640), .ZN(G45) );
  NOR2_X1 U708 ( .A1(n643), .A2(n641), .ZN(n642) );
  XOR2_X1 U709 ( .A(G146), .B(n642), .Z(G48) );
  NOR2_X1 U710 ( .A1(n647), .A2(n643), .ZN(n644) );
  XOR2_X1 U711 ( .A(KEYINPUT118), .B(n644), .Z(n645) );
  XNOR2_X1 U712 ( .A(G113), .B(n645), .ZN(G15) );
  NOR2_X1 U713 ( .A1(n647), .A2(n646), .ZN(n649) );
  XNOR2_X1 U714 ( .A(G116), .B(KEYINPUT119), .ZN(n648) );
  XNOR2_X1 U715 ( .A(n649), .B(n648), .ZN(G18) );
  XNOR2_X1 U716 ( .A(n650), .B(G125), .ZN(n651) );
  XNOR2_X1 U717 ( .A(n651), .B(KEYINPUT37), .ZN(G27) );
  NOR2_X1 U718 ( .A1(n717), .A2(KEYINPUT2), .ZN(n652) );
  XNOR2_X1 U719 ( .A(n652), .B(KEYINPUT81), .ZN(n653) );
  NAND2_X1 U720 ( .A1(n654), .A2(n653), .ZN(n657) );
  NOR2_X1 U721 ( .A1(n701), .A2(KEYINPUT2), .ZN(n655) );
  XNOR2_X1 U722 ( .A(n655), .B(KEYINPUT80), .ZN(n656) );
  NAND2_X1 U723 ( .A1(n658), .A2(n718), .ZN(n697) );
  XNOR2_X1 U724 ( .A(KEYINPUT121), .B(KEYINPUT52), .ZN(n688) );
  XOR2_X1 U725 ( .A(KEYINPUT50), .B(n660), .Z(n667) );
  NOR2_X1 U726 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U727 ( .A(n663), .B(KEYINPUT49), .ZN(n664) );
  NAND2_X1 U728 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U729 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U730 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U731 ( .A(KEYINPUT51), .B(n670), .Z(n671) );
  NOR2_X1 U732 ( .A1(n692), .A2(n671), .ZN(n686) );
  INV_X1 U733 ( .A(n672), .ZN(n691) );
  INV_X1 U734 ( .A(n677), .ZN(n673) );
  NOR2_X1 U735 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U736 ( .A1(n676), .A2(n675), .ZN(n682) );
  OR2_X1 U737 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U738 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U739 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U740 ( .A(n683), .B(KEYINPUT120), .ZN(n684) );
  NOR2_X1 U741 ( .A1(n691), .A2(n684), .ZN(n685) );
  NOR2_X1 U742 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U743 ( .A(n688), .B(n687), .Z(n689) );
  NOR2_X1 U744 ( .A1(n690), .A2(n689), .ZN(n694) );
  NOR2_X1 U745 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U746 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U747 ( .A(KEYINPUT122), .B(n695), .Z(n696) );
  NOR2_X1 U748 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U749 ( .A(KEYINPUT53), .B(n698), .ZN(G75) );
  NAND2_X1 U750 ( .A1(n700), .A2(n699), .ZN(n709) );
  NAND2_X1 U751 ( .A1(n701), .A2(n718), .ZN(n706) );
  NAND2_X1 U752 ( .A1(G224), .A2(G953), .ZN(n702) );
  XNOR2_X1 U753 ( .A(n702), .B(KEYINPUT61), .ZN(n703) );
  XNOR2_X1 U754 ( .A(KEYINPUT124), .B(n703), .ZN(n704) );
  NAND2_X1 U755 ( .A1(n704), .A2(G898), .ZN(n705) );
  NAND2_X1 U756 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U757 ( .A(n707), .B(KEYINPUT125), .ZN(n708) );
  XNOR2_X1 U758 ( .A(n709), .B(n708), .ZN(G69) );
  XOR2_X1 U759 ( .A(n710), .B(n711), .Z(n716) );
  XOR2_X1 U760 ( .A(G227), .B(n716), .Z(n712) );
  NAND2_X1 U761 ( .A1(n712), .A2(G900), .ZN(n713) );
  XOR2_X1 U762 ( .A(KEYINPUT126), .B(n713), .Z(n714) );
  NOR2_X1 U763 ( .A1(n718), .A2(n714), .ZN(n715) );
  XNOR2_X1 U764 ( .A(n715), .B(KEYINPUT127), .ZN(n721) );
  XNOR2_X1 U765 ( .A(n717), .B(n716), .ZN(n719) );
  NAND2_X1 U766 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U767 ( .A1(n721), .A2(n720), .ZN(G72) );
  XOR2_X1 U768 ( .A(G137), .B(n722), .Z(G39) );
  XOR2_X1 U769 ( .A(G140), .B(n723), .Z(G42) );
  XNOR2_X1 U770 ( .A(n724), .B(G119), .ZN(G21) );
endmodule

