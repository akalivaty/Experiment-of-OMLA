//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G125), .ZN(new_n191));
  INV_X1    g005(.A(G125), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G140), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT16), .ZN(new_n194));
  OR3_X1    g008(.A1(new_n192), .A2(KEYINPUT16), .A3(G140), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n194), .A2(new_n195), .A3(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(G119), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT68), .B(G128), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(G119), .ZN(new_n204));
  XOR2_X1   g018(.A(KEYINPUT24), .B(G110), .Z(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT74), .ZN(new_n207));
  AOI21_X1  g021(.A(KEYINPUT23), .B1(new_n201), .B2(G119), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(new_n202), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n201), .A2(KEYINPUT68), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT68), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G128), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n210), .A2(new_n212), .A3(KEYINPUT23), .A4(G119), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n209), .A2(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n207), .B1(new_n214), .B2(G110), .ZN(new_n215));
  INV_X1    g029(.A(G110), .ZN(new_n216));
  AOI211_X1 g030(.A(KEYINPUT74), .B(new_n216), .C1(new_n209), .C2(new_n213), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n200), .B(new_n206), .C1(new_n215), .C2(new_n217), .ZN(new_n218));
  OAI22_X1  g032(.A1(new_n214), .A2(G110), .B1(new_n204), .B2(new_n205), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n191), .A2(new_n193), .ZN(new_n220));
  AND2_X1   g034(.A1(KEYINPUT64), .A2(G146), .ZN(new_n221));
  NOR2_X1   g035(.A1(KEYINPUT64), .A2(G146), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT75), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n199), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n194), .A2(new_n195), .A3(KEYINPUT75), .A4(G146), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n219), .A2(new_n224), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G953), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(G221), .A3(G234), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n230), .B(KEYINPUT76), .ZN(new_n231));
  XNOR2_X1  g045(.A(KEYINPUT22), .B(G137), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n231), .B(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n218), .A2(new_n228), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n233), .B1(new_n218), .B2(new_n228), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n188), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT25), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n218), .A2(new_n228), .ZN(new_n240));
  INV_X1    g054(.A(new_n233), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n234), .ZN(new_n243));
  AOI21_X1  g057(.A(KEYINPUT25), .B1(new_n243), .B2(new_n188), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n189), .B1(new_n239), .B2(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n189), .A2(G902), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT64), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(new_n197), .ZN(new_n250));
  NAND2_X1  g064(.A1(KEYINPUT64), .A2(G146), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(G143), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G143), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT65), .A3(G146), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT65), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n255), .B1(new_n197), .B2(G143), .ZN(new_n256));
  AND2_X1   g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n252), .A2(new_n254), .A3(new_n256), .A4(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n197), .A2(G143), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n250), .A2(new_n251), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n260), .B1(new_n261), .B2(new_n253), .ZN(new_n262));
  NOR2_X1   g076(.A1(KEYINPUT0), .A2(G128), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n258), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT11), .ZN(new_n267));
  INV_X1    g081(.A(G134), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n267), .B1(new_n268), .B2(G137), .ZN(new_n269));
  INV_X1    g083(.A(G137), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT11), .A3(G134), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n268), .A2(G137), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G131), .ZN(new_n274));
  AND2_X1   g088(.A1(KEYINPUT66), .A2(G131), .ZN(new_n275));
  NOR2_X1   g089(.A1(KEYINPUT66), .A2(G131), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n277), .A2(new_n269), .A3(new_n271), .A4(new_n272), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT69), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n274), .A2(new_n278), .A3(KEYINPUT69), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n266), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n252), .A2(new_n254), .A3(new_n256), .A4(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n203), .B1(new_n252), .B2(KEYINPUT1), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n285), .B1(new_n286), .B2(new_n262), .ZN(new_n287));
  INV_X1    g101(.A(new_n273), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT67), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n289), .B1(new_n268), .B2(G137), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n270), .A2(KEYINPUT67), .A3(G134), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(new_n272), .A3(new_n291), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n288), .A2(new_n277), .B1(new_n292), .B2(G131), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n287), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT71), .B1(new_n283), .B2(new_n294), .ZN(new_n295));
  XOR2_X1   g109(.A(KEYINPUT2), .B(G113), .Z(new_n296));
  XNOR2_X1  g110(.A(G116), .B(G119), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n296), .B(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n252), .A2(new_n254), .A3(new_n256), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n259), .B1(new_n223), .B2(G143), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n300), .A2(new_n257), .B1(new_n301), .B2(new_n264), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n274), .A2(new_n278), .A3(KEYINPUT69), .ZN(new_n303));
  AOI21_X1  g117(.A(KEYINPUT69), .B1(new_n274), .B2(new_n278), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT71), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n287), .A2(new_n293), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n295), .A2(new_n299), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT28), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n305), .A2(new_n299), .A3(new_n307), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n301), .A2(new_n264), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n279), .A2(new_n313), .A3(new_n258), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n307), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n298), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n310), .B1(new_n312), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n311), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT26), .B(G101), .ZN(new_n320));
  NOR2_X1   g134(.A1(G237), .A2(G953), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G210), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n320), .B(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n323), .B(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT30), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n315), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n326), .B1(new_n287), .B2(new_n293), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n305), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n329), .A3(new_n298), .ZN(new_n330));
  INV_X1    g144(.A(new_n325), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n312), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT31), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n330), .A2(KEYINPUT31), .A3(new_n312), .A4(new_n331), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n319), .A2(new_n325), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(G472), .A2(G902), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT32), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n334), .A2(new_n335), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n305), .A2(new_n307), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n298), .B1(new_n341), .B2(KEYINPUT71), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT28), .B1(new_n342), .B2(new_n308), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n325), .B1(new_n343), .B2(new_n317), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT32), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n346), .A3(new_n337), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n339), .A2(new_n347), .ZN(new_n348));
  NOR3_X1   g162(.A1(new_n283), .A2(new_n294), .A3(new_n298), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n299), .B1(new_n305), .B2(new_n307), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT28), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT29), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n325), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n188), .B1(new_n354), .B2(new_n343), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT73), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n311), .A2(new_n318), .A3(new_n331), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n315), .A2(new_n326), .B1(new_n305), .B2(new_n328), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n349), .B1(new_n358), .B2(new_n298), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT72), .B1(new_n359), .B2(new_n331), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n330), .A2(new_n312), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT72), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n362), .A3(new_n325), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n357), .A2(new_n360), .A3(new_n352), .A4(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT73), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n365), .B(new_n188), .C1(new_n354), .C2(new_n343), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n356), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G472), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n248), .B1(new_n348), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(G113), .B(G122), .ZN(new_n370));
  INV_X1    g184(.A(G104), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n370), .B(new_n371), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n220), .A2(KEYINPUT19), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n220), .A2(KEYINPUT19), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n223), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OR2_X1    g189(.A1(new_n275), .A2(new_n276), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n321), .A2(G143), .A3(G214), .ZN(new_n377));
  AOI21_X1  g191(.A(G143), .B1(new_n321), .B2(G214), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G237), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(new_n229), .A3(G214), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n253), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n321), .A2(G143), .A3(G214), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n277), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n375), .A2(new_n385), .A3(new_n226), .A4(new_n227), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n224), .B1(new_n197), .B2(new_n220), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n382), .A2(new_n383), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(KEYINPUT18), .A3(G131), .ZN(new_n389));
  NAND2_X1  g203(.A1(KEYINPUT18), .A2(G131), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n382), .A2(new_n383), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n387), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n372), .B1(new_n386), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n392), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT17), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n379), .A2(new_n395), .A3(new_n384), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT89), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n397), .B1(new_n379), .B2(new_n395), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n388), .A2(KEYINPUT89), .A3(KEYINPUT17), .A4(new_n376), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n396), .A2(KEYINPUT90), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT90), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n379), .A2(new_n395), .A3(new_n384), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n200), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n394), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n372), .B(KEYINPUT88), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n393), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(G475), .A2(G902), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT20), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT20), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n398), .A2(new_n399), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n402), .A2(new_n401), .ZN(new_n412));
  INV_X1    g226(.A(new_n200), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n379), .A2(new_n384), .A3(KEYINPUT90), .A4(new_n395), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n411), .A2(new_n412), .A3(new_n413), .A4(new_n414), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n415), .A2(new_n392), .A3(new_n405), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n410), .B(new_n407), .C1(new_n416), .C2(new_n393), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n409), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n415), .A2(new_n392), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT91), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n372), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n415), .A2(KEYINPUT91), .A3(new_n392), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n416), .ZN(new_n425));
  AOI21_X1  g239(.A(G902), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G475), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n418), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n229), .A2(G952), .ZN(new_n430));
  NAND2_X1  g244(.A1(G234), .A2(G237), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(KEYINPUT96), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n431), .A2(G902), .A3(G953), .ZN(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(G898), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G122), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT92), .B1(new_n439), .B2(G116), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT92), .ZN(new_n441));
  INV_X1    g255(.A(G116), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n441), .A2(new_n442), .A3(G122), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n444), .A2(KEYINPUT14), .B1(G116), .B2(new_n439), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n445), .B1(KEYINPUT14), .B2(new_n444), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G107), .ZN(new_n447));
  INV_X1    g261(.A(G107), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT93), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n439), .A2(G116), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n444), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n449), .B1(new_n444), .B2(new_n450), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n448), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n201), .A2(G143), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n210), .A2(new_n212), .A3(G143), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT94), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n203), .A2(KEYINPUT94), .A3(G143), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n455), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(new_n268), .ZN(new_n461));
  AOI211_X1 g275(.A(G134), .B(new_n455), .C1(new_n458), .C2(new_n459), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n447), .B(new_n454), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n455), .A2(KEYINPUT13), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n455), .A2(KEYINPUT13), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(KEYINPUT94), .B1(new_n203), .B2(G143), .ZN(new_n468));
  AND4_X1   g282(.A1(KEYINPUT94), .A2(new_n210), .A3(new_n212), .A4(G143), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n465), .B1(new_n470), .B2(KEYINPUT95), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n466), .B1(new_n458), .B2(new_n459), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT95), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n268), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n460), .A2(new_n268), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n452), .A2(new_n453), .A3(new_n448), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n444), .A2(new_n450), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT93), .ZN(new_n479));
  AOI21_X1  g293(.A(G107), .B1(new_n479), .B2(new_n451), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n476), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n463), .B1(new_n475), .B2(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(KEYINPUT9), .B(G234), .ZN(new_n483));
  NOR3_X1   g297(.A1(new_n483), .A2(new_n187), .A3(G953), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n463), .B(new_n484), .C1(new_n475), .C2(new_n481), .ZN(new_n487));
  AOI21_X1  g301(.A(G902), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G478), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n489), .A2(KEYINPUT15), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n488), .B(new_n490), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n429), .A2(KEYINPUT97), .A3(new_n438), .A4(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT97), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n488), .B1(KEYINPUT15), .B2(new_n489), .ZN(new_n494));
  INV_X1    g308(.A(new_n487), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n464), .B1(new_n472), .B2(new_n473), .ZN(new_n496));
  AOI211_X1 g310(.A(KEYINPUT95), .B(new_n466), .C1(new_n458), .C2(new_n459), .ZN(new_n497));
  OAI21_X1  g311(.A(G134), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n479), .A2(G107), .A3(new_n451), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n462), .B1(new_n454), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n484), .B1(new_n501), .B2(new_n463), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n188), .B1(new_n495), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n490), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n494), .A2(new_n504), .A3(new_n438), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n493), .B1(new_n505), .B2(new_n428), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n492), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(G221), .B1(new_n483), .B2(G902), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(KEYINPUT77), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n303), .A2(new_n304), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT78), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n448), .B2(G104), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n371), .A2(KEYINPUT78), .A3(G107), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n448), .A2(KEYINPUT3), .A3(G104), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT3), .B1(new_n448), .B2(G104), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n512), .B(new_n513), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT4), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n517), .A3(G101), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n518), .A2(new_n258), .A3(new_n313), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n516), .A2(G101), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT3), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n521), .B1(new_n371), .B2(G107), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n448), .A2(KEYINPUT3), .A3(G104), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(G101), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n524), .A2(new_n525), .A3(new_n512), .A4(new_n513), .ZN(new_n526));
  AND4_X1   g340(.A1(KEYINPUT79), .A2(new_n520), .A3(KEYINPUT4), .A4(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n517), .B1(new_n516), .B2(G101), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT79), .B1(new_n528), .B2(new_n526), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n519), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT80), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n531), .B1(new_n371), .B2(G107), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n371), .A2(G107), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n448), .A2(KEYINPUT80), .A3(G104), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(G101), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n256), .A2(new_n254), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n259), .A2(KEYINPUT1), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n537), .A2(new_n252), .B1(G128), .B2(new_n538), .ZN(new_n539));
  AND4_X1   g353(.A1(new_n252), .A2(new_n254), .A3(new_n256), .A4(new_n284), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n526), .B(new_n536), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  XOR2_X1   g355(.A(KEYINPUT81), .B(KEYINPUT10), .Z(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n526), .A2(KEYINPUT10), .A3(new_n536), .ZN(new_n544));
  AOI22_X1  g358(.A1(new_n541), .A2(new_n543), .B1(new_n287), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n510), .B1(new_n530), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n530), .A2(new_n545), .A3(new_n510), .ZN(new_n547));
  XNOR2_X1  g361(.A(G110), .B(G140), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n229), .A2(G227), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n548), .B(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT83), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n546), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n547), .A2(KEYINPUT83), .A3(new_n551), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n526), .A2(new_n536), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n541), .B(KEYINPUT82), .C1(new_n287), .C2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n510), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n557), .A2(new_n287), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n537), .A2(new_n252), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n538), .A2(G128), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n556), .B1(new_n285), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT82), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(KEYINPUT12), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n558), .B(new_n559), .C1(new_n565), .C2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n279), .B1(new_n560), .B2(new_n564), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT12), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n568), .A2(new_n547), .A3(new_n570), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n554), .A2(new_n555), .B1(new_n571), .B2(new_n550), .ZN(new_n572));
  OAI21_X1  g386(.A(G469), .B1(new_n572), .B2(G902), .ZN(new_n573));
  INV_X1    g387(.A(G469), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n530), .A2(new_n510), .A3(new_n545), .ZN(new_n575));
  OAI211_X1 g389(.A(KEYINPUT84), .B(new_n550), .C1(new_n575), .C2(new_n546), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n568), .A2(new_n551), .A3(new_n547), .A4(new_n570), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n302), .A2(new_n518), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n528), .A2(new_n526), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT79), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n528), .A2(KEYINPUT79), .A3(new_n526), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n579), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n544), .A2(new_n287), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n585), .B1(new_n564), .B2(new_n542), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n559), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n547), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT84), .B1(new_n588), .B2(new_n550), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n574), .B(new_n188), .C1(new_n578), .C2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n509), .B1(new_n573), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(G214), .B1(G237), .B2(G902), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(G110), .B(G122), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n298), .A2(new_n518), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n596), .B1(new_n582), .B2(new_n583), .ZN(new_n597));
  INV_X1    g411(.A(G119), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(G116), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n442), .A2(G119), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(new_n600), .A3(KEYINPUT5), .ZN(new_n601));
  OR3_X1    g415(.A1(new_n442), .A2(KEYINPUT5), .A3(G119), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n602), .A3(G113), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n296), .A2(new_n297), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n526), .A2(new_n536), .A3(new_n603), .A4(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n595), .B1(new_n597), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n596), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n608), .B1(new_n527), .B2(new_n529), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(new_n605), .A3(new_n594), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n607), .A2(KEYINPUT6), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT6), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n612), .B(new_n595), .C1(new_n597), .C2(new_n606), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n192), .B(new_n285), .C1(new_n286), .C2(new_n262), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n192), .B1(new_n313), .B2(new_n258), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n229), .A2(G224), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n611), .A2(new_n613), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT87), .ZN(new_n621));
  OAI211_X1 g435(.A(KEYINPUT7), .B(new_n618), .C1(new_n615), .C2(new_n616), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n266), .A2(G125), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n618), .A2(KEYINPUT7), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n614), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n603), .A2(new_n604), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n556), .A2(KEYINPUT86), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT85), .B(KEYINPUT8), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n594), .B(new_n628), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n556), .A2(new_n626), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT86), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n631), .A2(new_n632), .A3(new_n605), .ZN(new_n633));
  AOI22_X1  g447(.A1(new_n622), .A2(new_n625), .B1(new_n630), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n610), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n621), .B1(new_n635), .B2(new_n188), .ZN(new_n636));
  AOI211_X1 g450(.A(KEYINPUT87), .B(G902), .C1(new_n634), .C2(new_n610), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n620), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(G210), .B1(G237), .B2(G902), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n620), .B(new_n639), .C1(new_n636), .C2(new_n637), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n593), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n369), .A2(new_n507), .A3(new_n591), .A4(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G101), .ZN(G3));
  INV_X1    g459(.A(new_n610), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n633), .A2(new_n627), .A3(new_n629), .ZN(new_n647));
  INV_X1    g461(.A(new_n625), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n624), .B1(new_n623), .B2(new_n614), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n188), .B1(new_n646), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(KEYINPUT87), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n635), .A2(new_n621), .A3(new_n188), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n639), .B1(new_n654), .B2(new_n620), .ZN(new_n655));
  INV_X1    g469(.A(new_n642), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n592), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(new_n437), .ZN(new_n658));
  INV_X1    g472(.A(new_n248), .ZN(new_n659));
  AOI21_X1  g473(.A(G902), .B1(new_n340), .B2(new_n344), .ZN(new_n660));
  INV_X1    g474(.A(G472), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n662), .B1(new_n337), .B2(new_n345), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n658), .A2(new_n659), .A3(new_n591), .A4(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n489), .A2(G902), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(KEYINPUT98), .B1(new_n495), .B2(new_n502), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT33), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n668), .B1(new_n501), .B2(new_n463), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(KEYINPUT33), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n486), .A2(new_n487), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n482), .A2(KEYINPUT33), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n668), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n672), .A2(new_n674), .A3(KEYINPUT98), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n666), .B1(new_n671), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n488), .A2(G478), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n428), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n664), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT99), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT34), .B(G104), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G6));
  NOR3_X1   g496(.A1(new_n491), .A2(new_n428), .A3(new_n437), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n643), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT100), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT100), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n643), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n663), .A2(new_n659), .A3(new_n591), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT35), .B(G107), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G9));
  NOR2_X1   g506(.A1(new_n233), .A2(KEYINPUT36), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n240), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n246), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n245), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n657), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n698), .A2(new_n507), .A3(new_n591), .A4(new_n663), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT37), .B(G110), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G12));
  NOR2_X1   g515(.A1(new_n491), .A2(new_n428), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(G900), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n434), .A2(new_n704), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n433), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n348), .A2(new_n368), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n698), .A2(new_n707), .A3(new_n708), .A4(new_n591), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G128), .ZN(G30));
  XOR2_X1   g524(.A(new_n706), .B(KEYINPUT39), .Z(new_n711));
  NAND2_X1  g525(.A1(new_n591), .A2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT102), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT40), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n712), .B(KEYINPUT102), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(KEYINPUT40), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n641), .A2(new_n642), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(KEYINPUT38), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n359), .A2(new_n325), .ZN(new_n721));
  INV_X1    g535(.A(new_n350), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(new_n312), .A3(new_n325), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n188), .ZN(new_n724));
  OAI21_X1  g538(.A(G472), .B1(new_n721), .B2(new_n724), .ZN(new_n725));
  XOR2_X1   g539(.A(new_n725), .B(KEYINPUT101), .Z(new_n726));
  AOI21_X1  g540(.A(new_n696), .B1(new_n726), .B2(new_n348), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n372), .B1(new_n419), .B2(new_n420), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n416), .B1(new_n728), .B2(new_n423), .ZN(new_n729));
  OAI21_X1  g543(.A(G475), .B1(new_n729), .B2(G902), .ZN(new_n730));
  AOI22_X1  g544(.A1(new_n730), .A2(new_n418), .B1(new_n494), .B2(new_n504), .ZN(new_n731));
  AND4_X1   g545(.A1(new_n592), .A2(new_n720), .A3(new_n727), .A4(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n716), .A2(new_n718), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(KEYINPUT103), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G143), .ZN(G45));
  INV_X1    g549(.A(new_n706), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n428), .B(new_n736), .C1(new_n676), .C2(new_n677), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n698), .A2(new_n708), .A3(new_n591), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G146), .ZN(G48));
  NOR3_X1   g554(.A1(new_n657), .A2(new_n437), .A3(new_n678), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n188), .B1(new_n578), .B2(new_n589), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(G469), .ZN(new_n743));
  INV_X1    g557(.A(new_n509), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(new_n744), .A3(new_n590), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n741), .A2(new_n369), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(KEYINPUT41), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G113), .ZN(G15));
  AND3_X1   g563(.A1(new_n643), .A2(new_n683), .A3(new_n686), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n686), .B1(new_n643), .B2(new_n683), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n369), .B(new_n746), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G116), .ZN(G18));
  NOR2_X1   g567(.A1(new_n657), .A2(new_n745), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n754), .A2(new_n708), .A3(new_n507), .A4(new_n696), .ZN(new_n755));
  XOR2_X1   g569(.A(KEYINPUT104), .B(G119), .Z(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(G21));
  INV_X1    g571(.A(KEYINPUT105), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n245), .A2(new_n758), .A3(new_n247), .ZN(new_n759));
  INV_X1    g573(.A(new_n189), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n237), .A2(new_n238), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n243), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n247), .ZN(new_n764));
  OAI21_X1  g578(.A(KEYINPUT105), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n759), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(G472), .B1(new_n336), .B2(G902), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n334), .A2(new_n335), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n331), .B1(new_n311), .B2(new_n351), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n337), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n766), .A2(new_n767), .A3(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n743), .A2(new_n438), .A3(new_n744), .A4(new_n590), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n643), .A2(KEYINPUT106), .A3(new_n731), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT106), .B1(new_n643), .B2(new_n731), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G122), .ZN(G24));
  OAI211_X1 g591(.A(new_n770), .B(new_n696), .C1(new_n661), .C2(new_n660), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(new_n737), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n754), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT107), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n754), .A2(new_n779), .A3(KEYINPUT107), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G125), .ZN(G27));
  INV_X1    g599(.A(KEYINPUT42), .ZN(new_n786));
  INV_X1    g600(.A(new_n590), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n554), .A2(new_n555), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n571), .A2(new_n550), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(G469), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(G469), .A2(G902), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n744), .B1(new_n787), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n641), .A2(new_n592), .A3(new_n642), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n793), .A2(new_n737), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n766), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(new_n348), .B2(new_n368), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n786), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n794), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n737), .A2(KEYINPUT42), .ZN(new_n800));
  AND4_X1   g614(.A1(new_n369), .A2(new_n591), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G131), .ZN(G33));
  NOR2_X1   g617(.A1(new_n793), .A2(new_n794), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n369), .A3(new_n707), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G134), .ZN(G36));
  OAI21_X1  g620(.A(new_n429), .B1(new_n676), .B2(new_n677), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n807), .B(KEYINPUT43), .Z(new_n808));
  NOR2_X1   g622(.A1(new_n663), .A2(new_n697), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT44), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n572), .A2(KEYINPUT45), .ZN(new_n812));
  OAI21_X1  g626(.A(G469), .B1(new_n572), .B2(KEYINPUT45), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n791), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT46), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n590), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n815), .A2(new_n816), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n744), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n711), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XOR2_X1   g636(.A(new_n794), .B(KEYINPUT108), .Z(new_n823));
  NAND3_X1  g637(.A1(new_n811), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G137), .ZN(G39));
  XNOR2_X1  g639(.A(new_n820), .B(KEYINPUT47), .ZN(new_n826));
  OR4_X1    g640(.A1(new_n708), .A2(new_n659), .A3(new_n737), .A4(new_n794), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(G140), .ZN(G42));
  NAND2_X1  g643(.A1(new_n726), .A2(new_n348), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n796), .A2(new_n807), .A3(new_n509), .A4(new_n593), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT109), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n743), .A2(new_n590), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT49), .ZN(new_n834));
  OR4_X1    g648(.A1(new_n830), .A2(new_n832), .A3(new_n720), .A4(new_n834), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n754), .A2(KEYINPUT107), .A3(new_n779), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT107), .B1(new_n754), .B2(new_n779), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n709), .B(new_n739), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n643), .A2(new_n731), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT106), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n643), .A2(KEYINPUT106), .A3(new_n731), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n793), .A2(new_n706), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n843), .A2(new_n727), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT52), .B1(new_n838), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n708), .A2(new_n591), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n643), .A2(new_n702), .A3(new_n696), .A4(new_n736), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n849), .B1(new_n782), .B2(new_n783), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT52), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n843), .A2(new_n727), .A3(new_n844), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n850), .A2(new_n851), .A3(new_n739), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n846), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT111), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n776), .A2(new_n755), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n699), .A2(new_n644), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n369), .A2(new_n746), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n858), .B1(new_n688), .B2(new_n741), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n678), .A2(KEYINPUT110), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT110), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n861), .B(new_n428), .C1(new_n676), .C2(new_n677), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n860), .A2(new_n703), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n689), .A2(new_n658), .A3(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n856), .A2(new_n857), .A3(new_n859), .A4(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n778), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n866), .A2(new_n738), .A3(new_n591), .A4(new_n799), .ZN(new_n867));
  AND4_X1   g681(.A1(new_n429), .A2(new_n491), .A3(new_n696), .A4(new_n736), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n708), .A2(new_n868), .A3(new_n591), .A4(new_n799), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n805), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n802), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n855), .B1(new_n865), .B2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n752), .A2(new_n776), .A3(new_n747), .A4(new_n755), .ZN(new_n873));
  INV_X1    g687(.A(new_n863), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n644), .B(new_n699), .C1(new_n664), .C2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n805), .A2(new_n867), .A3(new_n869), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n877), .A2(new_n798), .A3(new_n801), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n876), .A2(KEYINPUT111), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n854), .B1(new_n872), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT112), .B1(new_n880), .B2(KEYINPUT53), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n846), .A2(new_n853), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n865), .A2(new_n871), .A3(new_n855), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT111), .B1(new_n876), .B2(new_n878), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT112), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT53), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n865), .A2(new_n871), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n709), .B1(new_n836), .B2(new_n837), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n887), .B1(new_n890), .B2(KEYINPUT52), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n882), .A2(KEYINPUT113), .A3(new_n889), .A4(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT113), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n891), .A2(new_n876), .A3(new_n878), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n893), .B1(new_n894), .B2(new_n854), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT54), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n881), .A2(new_n888), .A3(new_n896), .A4(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT53), .B1(new_n890), .B2(KEYINPUT52), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n885), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n880), .A2(KEYINPUT53), .ZN(new_n901));
  OAI21_X1  g715(.A(KEYINPUT54), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n433), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n808), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n771), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n754), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n430), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n745), .A2(new_n794), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n905), .A2(new_n797), .A3(new_n910), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT48), .Z(new_n912));
  INV_X1    g726(.A(new_n678), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n830), .A2(new_n248), .A3(new_n433), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n910), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT116), .Z(new_n916));
  AOI211_X1 g730(.A(new_n909), .B(new_n912), .C1(new_n913), .C2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n826), .B1(new_n744), .B2(new_n833), .ZN(new_n918));
  INV_X1    g732(.A(new_n907), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n918), .A2(new_n823), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n905), .A2(new_n910), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n921), .A2(new_n778), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n676), .A2(new_n428), .A3(new_n677), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n922), .B1(new_n916), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n907), .A2(new_n720), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n746), .A2(new_n593), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT114), .Z(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AOI211_X1 g742(.A(KEYINPUT115), .B(KEYINPUT50), .C1(new_n925), .C2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(KEYINPUT115), .A2(KEYINPUT50), .ZN(new_n930));
  NOR4_X1   g744(.A1(new_n907), .A2(new_n927), .A3(new_n720), .A4(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n924), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n920), .A2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT51), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n917), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n934), .B1(new_n920), .B2(new_n932), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n936), .A2(KEYINPUT117), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(KEYINPUT117), .ZN(new_n938));
  AOI211_X1 g752(.A(new_n903), .B(new_n935), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(G952), .A2(G953), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n835), .B1(new_n939), .B2(new_n940), .ZN(G75));
  INV_X1    g755(.A(KEYINPUT118), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n881), .A2(new_n888), .A3(new_n896), .ZN(new_n943));
  AND2_X1   g757(.A1(G210), .A2(G902), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT56), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n611), .A2(new_n613), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(new_n619), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT55), .Z(new_n950));
  AOI21_X1  g764(.A(new_n942), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT56), .B1(new_n943), .B2(new_n944), .ZN(new_n952));
  INV_X1    g766(.A(new_n950), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n952), .A2(KEYINPUT118), .A3(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n229), .A2(G952), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n943), .A2(KEYINPUT119), .A3(new_n944), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n950), .A2(KEYINPUT56), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT119), .B1(new_n943), .B2(new_n944), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(KEYINPUT120), .B1(new_n955), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n962), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT120), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n947), .A2(new_n942), .A3(new_n950), .ZN(new_n966));
  OAI21_X1  g780(.A(KEYINPUT118), .B1(new_n952), .B2(new_n953), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n964), .A2(new_n965), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n963), .A2(new_n969), .ZN(G51));
  NAND2_X1  g784(.A1(new_n943), .A2(KEYINPUT54), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n898), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n791), .B(KEYINPUT57), .Z(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(KEYINPUT121), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT121), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n972), .A2(new_n976), .A3(new_n973), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n975), .B(new_n977), .C1(new_n589), .C2(new_n578), .ZN(new_n978));
  INV_X1    g792(.A(new_n814), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n943), .A2(G902), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n956), .B1(new_n978), .B2(new_n980), .ZN(G54));
  NAND4_X1  g795(.A1(new_n943), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n982), .A2(new_n406), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n982), .A2(new_n406), .ZN(new_n984));
  NOR3_X1   g798(.A1(new_n983), .A2(new_n984), .A3(new_n956), .ZN(G60));
  NAND2_X1  g799(.A1(new_n671), .A2(new_n675), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT122), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(G478), .A2(G902), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT59), .Z(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n988), .B1(new_n903), .B2(new_n991), .ZN(new_n992));
  OR2_X1    g806(.A1(new_n992), .A2(KEYINPUT123), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(KEYINPUT123), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n987), .A2(new_n990), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n956), .B1(new_n972), .B2(new_n995), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n993), .A2(new_n994), .A3(new_n996), .ZN(G63));
  NAND2_X1  g811(.A1(G217), .A2(G902), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT60), .Z(new_n999));
  AOI21_X1  g813(.A(new_n243), .B1(new_n943), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n1000), .A2(new_n956), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n943), .A2(new_n694), .A3(new_n999), .ZN(new_n1002));
  AOI22_X1  g816(.A1(new_n1001), .A2(new_n1002), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n1003));
  NOR2_X1   g817(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1003), .B(new_n1004), .ZN(G66));
  INV_X1    g819(.A(G224), .ZN(new_n1006));
  OAI21_X1  g820(.A(G953), .B1(new_n435), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1007), .B1(new_n876), .B2(G953), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n948), .B1(G898), .B2(new_n229), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1008), .B(new_n1009), .ZN(G69));
  NOR2_X1   g824(.A1(new_n373), .A2(new_n374), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n358), .B(new_n1011), .Z(new_n1012));
  INV_X1    g826(.A(new_n838), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n734), .A2(new_n1013), .ZN(new_n1014));
  OR2_X1    g828(.A1(new_n1014), .A2(KEYINPUT62), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n714), .A2(new_n369), .A3(new_n799), .A4(new_n863), .ZN(new_n1016));
  AND3_X1   g830(.A1(new_n828), .A2(new_n824), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1014), .A2(KEYINPUT62), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1015), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1012), .B1(new_n1019), .B2(new_n229), .ZN(new_n1020));
  OR2_X1    g834(.A1(new_n1020), .A2(KEYINPUT125), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1020), .A2(KEYINPUT125), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n802), .A2(new_n805), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(KEYINPUT126), .Z(new_n1024));
  AND2_X1   g838(.A1(new_n843), .A2(new_n797), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n838), .B1(new_n822), .B2(new_n1025), .ZN(new_n1026));
  AND4_X1   g840(.A1(new_n824), .A2(new_n828), .A3(new_n1024), .A4(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1027), .A2(new_n229), .ZN(new_n1028));
  OAI211_X1 g842(.A(new_n1028), .B(new_n1012), .C1(new_n704), .C2(new_n229), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1021), .A2(new_n1022), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n229), .B1(G227), .B2(G900), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1031), .ZN(new_n1033));
  NAND4_X1  g847(.A1(new_n1021), .A2(new_n1033), .A3(new_n1022), .A4(new_n1029), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1032), .A2(new_n1034), .ZN(G72));
  XNOR2_X1  g849(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1036));
  NAND2_X1  g850(.A1(G472), .A2(G902), .ZN(new_n1037));
  XNOR2_X1  g851(.A(new_n1036), .B(new_n1037), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n360), .A2(new_n332), .A3(new_n363), .ZN(new_n1039));
  OAI211_X1 g853(.A(new_n1038), .B(new_n1039), .C1(new_n900), .C2(new_n901), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1040), .A2(new_n957), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1027), .A2(new_n876), .ZN(new_n1042));
  AOI211_X1 g856(.A(new_n331), .B(new_n361), .C1(new_n1042), .C2(new_n1038), .ZN(new_n1043));
  OAI21_X1  g857(.A(new_n1038), .B1(new_n1019), .B2(new_n865), .ZN(new_n1044));
  AOI211_X1 g858(.A(new_n1041), .B(new_n1043), .C1(new_n721), .C2(new_n1044), .ZN(G57));
endmodule


