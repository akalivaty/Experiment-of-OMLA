//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 0 0 1 1 1 0 1 0 1 0 0 0 1 1 1 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND3_X1   g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n187), .B(new_n189), .Z(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G125), .ZN(new_n193));
  INV_X1    g007(.A(G125), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G140), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n193), .A2(new_n195), .A3(KEYINPUT16), .ZN(new_n196));
  OR3_X1    g010(.A1(new_n194), .A2(KEYINPUT16), .A3(G140), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(G146), .ZN(new_n198));
  XNOR2_X1  g012(.A(G125), .B(G140), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n198), .A2(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT65), .B(G128), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(KEYINPUT23), .A3(G119), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  AOI21_X1  g019(.A(KEYINPUT23), .B1(new_n205), .B2(G119), .ZN(new_n206));
  INV_X1    g020(.A(G119), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n204), .A2(new_n208), .ZN(new_n209));
  OR2_X1    g023(.A1(new_n209), .A2(G110), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n203), .A2(G119), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n211), .B1(G119), .B2(new_n205), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT24), .B(G110), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT75), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT75), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n210), .A2(new_n217), .A3(new_n214), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n202), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n209), .A2(G110), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n220), .B(KEYINPUT73), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n196), .A2(new_n197), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n200), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT74), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n224), .A3(new_n198), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n222), .A2(KEYINPUT74), .A3(new_n200), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n225), .B(new_n226), .C1(new_n212), .C2(new_n213), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n221), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n191), .B1(new_n219), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n202), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n210), .A2(new_n217), .A3(new_n214), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n217), .B1(new_n210), .B2(new_n214), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n233), .B(new_n190), .C1(new_n221), .C2(new_n227), .ZN(new_n234));
  INV_X1    g048(.A(G902), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n229), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT25), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n229), .A2(new_n234), .A3(KEYINPUT25), .A4(new_n235), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G217), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n241), .B1(G234), .B2(new_n235), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n229), .A2(new_n234), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n242), .A2(G902), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G137), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(KEYINPUT11), .A3(G134), .ZN(new_n249));
  INV_X1    g063(.A(G134), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G137), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT11), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n253), .B1(new_n250), .B2(G137), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT64), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n248), .A2(G134), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT64), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(new_n257), .A3(new_n253), .ZN(new_n258));
  AOI211_X1 g072(.A(G131), .B(new_n252), .C1(new_n255), .C2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G131), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n255), .A2(new_n258), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n249), .A2(new_n251), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n200), .A2(G143), .ZN(new_n265));
  INV_X1    g079(.A(G143), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G146), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n265), .A2(new_n267), .A3(KEYINPUT0), .A4(G128), .ZN(new_n268));
  XNOR2_X1  g082(.A(G143), .B(G146), .ZN(new_n269));
  OR2_X1    g083(.A1(KEYINPUT0), .A2(G128), .ZN(new_n270));
  NAND2_X1  g084(.A1(KEYINPUT0), .A2(G128), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n268), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT66), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT66), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n268), .B(new_n275), .C1(new_n269), .C2(new_n272), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT67), .B1(new_n264), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n261), .A2(new_n262), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G131), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n257), .B1(new_n256), .B2(new_n253), .ZN(new_n281));
  AOI211_X1 g095(.A(KEYINPUT64), .B(KEYINPUT11), .C1(new_n248), .C2(G134), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n262), .B(new_n260), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n276), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n265), .A2(new_n267), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(new_n271), .A3(new_n270), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n275), .B1(new_n287), .B2(new_n268), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT67), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n284), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT1), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n292), .B1(G143), .B2(new_n200), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n286), .B1(new_n203), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n269), .A2(new_n292), .A3(G128), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n256), .A2(new_n251), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G131), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n296), .A2(new_n283), .A3(new_n298), .ZN(new_n299));
  XOR2_X1   g113(.A(G116), .B(G119), .Z(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT2), .B(G113), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n300), .B(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n278), .A2(new_n291), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n273), .B1(new_n280), .B2(new_n283), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(new_n299), .ZN(new_n307));
  INV_X1    g121(.A(new_n302), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT28), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n303), .B1(new_n264), .B2(new_n277), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT28), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  XOR2_X1   g129(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n316));
  NOR2_X1   g130(.A1(G237), .A2(G953), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G210), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n316), .B(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT26), .B(G101), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n319), .B(new_n320), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n315), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT30), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n299), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n278), .A2(new_n291), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT68), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT68), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n278), .A2(new_n291), .A3(new_n325), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n324), .B1(new_n306), .B2(new_n299), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n302), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT69), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT69), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n330), .A2(new_n336), .A3(new_n333), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n321), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n305), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT31), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n336), .B1(new_n330), .B2(new_n333), .ZN(new_n342));
  AOI211_X1 g156(.A(KEYINPUT69), .B(new_n332), .C1(new_n327), .C2(new_n329), .ZN(new_n343));
  OAI211_X1 g157(.A(KEYINPUT31), .B(new_n340), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n323), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT71), .ZN(new_n347));
  NOR2_X1   g161(.A1(G472), .A2(G902), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n340), .B1(new_n342), .B2(new_n343), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT31), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n322), .B1(new_n352), .B2(new_n344), .ZN(new_n353));
  INV_X1    g167(.A(new_n348), .ZN(new_n354));
  OAI21_X1  g168(.A(KEYINPUT71), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT32), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n349), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n352), .A2(new_n344), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n354), .B1(new_n358), .B2(new_n323), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT29), .B1(new_n315), .B2(new_n321), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n305), .B1(new_n335), .B2(new_n337), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n360), .B1(new_n361), .B2(new_n321), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n278), .A2(new_n291), .ZN(new_n363));
  INV_X1    g177(.A(new_n299), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n305), .B1(new_n365), .B2(new_n302), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n366), .A2(new_n312), .ZN(new_n367));
  XOR2_X1   g181(.A(new_n313), .B(KEYINPUT72), .Z(new_n368));
  NOR2_X1   g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n321), .A2(KEYINPUT29), .ZN(new_n370));
  AOI21_X1  g184(.A(G902), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n362), .A2(new_n371), .ZN(new_n372));
  AOI22_X1  g186(.A1(new_n359), .A2(KEYINPUT32), .B1(new_n372), .B2(G472), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n247), .B1(new_n357), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT9), .B(G234), .ZN(new_n375));
  OAI21_X1  g189(.A(G221), .B1(new_n375), .B2(G902), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT12), .ZN(new_n378));
  INV_X1    g192(.A(G104), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT3), .B1(new_n379), .B2(G107), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT3), .ZN(new_n381));
  INV_X1    g195(.A(G107), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(G104), .ZN(new_n383));
  INV_X1    g197(.A(G101), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n379), .A2(G107), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n380), .A2(new_n383), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n379), .A2(G107), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n382), .A2(G104), .ZN(new_n388));
  OAI21_X1  g202(.A(G101), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n265), .A2(KEYINPUT1), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n269), .B1(G128), .B2(new_n390), .ZN(new_n391));
  AND4_X1   g205(.A1(new_n292), .A2(new_n265), .A3(new_n267), .A4(G128), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n386), .B(new_n389), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n386), .A2(new_n389), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n393), .B1(new_n296), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n378), .B1(new_n395), .B2(new_n284), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n380), .A2(new_n383), .A3(new_n385), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G101), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(KEYINPUT4), .A3(new_n386), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n398), .A2(new_n401), .A3(G101), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n400), .A2(new_n274), .A3(new_n276), .A4(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT10), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n393), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n394), .A2(new_n296), .A3(KEYINPUT10), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n403), .A2(new_n405), .A3(new_n264), .A4(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n395), .A2(new_n378), .A3(new_n284), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n397), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(G110), .B(G140), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n188), .A2(G227), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n410), .B(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n403), .A2(new_n405), .A3(new_n406), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n284), .ZN(new_n415));
  INV_X1    g229(.A(new_n412), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n407), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n235), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G469), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT76), .B(G469), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n415), .A2(new_n407), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n412), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(KEYINPUT77), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n397), .A2(new_n407), .A3(new_n408), .A4(new_n416), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n416), .B1(new_n415), .B2(new_n407), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT77), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n235), .B(new_n421), .C1(new_n424), .C2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n377), .B1(new_n420), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(G214), .B1(G237), .B2(G902), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n273), .A2(G125), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n433), .B1(G125), .B2(new_n296), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT7), .ZN(new_n435));
  INV_X1    g249(.A(G224), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n436), .A2(G953), .ZN(new_n437));
  OR3_X1    g251(.A1(new_n434), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(G110), .B(G122), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(KEYINPUT8), .ZN(new_n440));
  OR2_X1    g254(.A1(new_n300), .A2(new_n301), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT5), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n442), .A2(new_n207), .A3(G116), .ZN(new_n443));
  OAI211_X1 g257(.A(G113), .B(new_n443), .C1(new_n300), .C2(new_n442), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n394), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n394), .B1(new_n441), .B2(new_n444), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n440), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n302), .A2(new_n402), .ZN(new_n449));
  INV_X1    g263(.A(new_n400), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n439), .B(new_n445), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n434), .B1(new_n435), .B2(new_n437), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n438), .A2(new_n448), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n235), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT78), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n445), .B1(new_n449), .B2(new_n450), .ZN(new_n457));
  INV_X1    g271(.A(new_n439), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(KEYINPUT6), .A3(new_n451), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n434), .B(new_n437), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT6), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n457), .A2(new_n462), .A3(new_n458), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n460), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n453), .A2(KEYINPUT78), .A3(new_n235), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n456), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(G210), .B1(G237), .B2(G902), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(KEYINPUT79), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n468), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n456), .A2(new_n470), .A3(new_n464), .A4(new_n465), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n432), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n430), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(G122), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(G116), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n382), .B1(new_n475), .B2(KEYINPUT14), .ZN(new_n476));
  XNOR2_X1  g290(.A(G116), .B(G122), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n476), .B(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n203), .A2(G143), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n205), .A2(G143), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n479), .A2(new_n250), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n250), .B1(new_n479), .B2(new_n481), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n478), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  XOR2_X1   g299(.A(G116), .B(G122), .Z(new_n486));
  INV_X1    g300(.A(KEYINPUT84), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n477), .A2(KEYINPUT84), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G107), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n488), .A2(new_n489), .A3(new_n382), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(new_n482), .A3(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n480), .A2(KEYINPUT13), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n494), .B(KEYINPUT85), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n203), .A2(G143), .B1(KEYINPUT13), .B2(new_n480), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n250), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n485), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  NOR3_X1   g312(.A1(new_n375), .A2(new_n241), .A3(G953), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n485), .B(new_n499), .C1(new_n493), .C2(new_n497), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(KEYINPUT86), .B1(new_n503), .B2(new_n235), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT86), .ZN(new_n505));
  AOI211_X1 g319(.A(new_n505), .B(G902), .C1(new_n501), .C2(new_n502), .ZN(new_n506));
  INV_X1    g320(.A(G478), .ZN(new_n507));
  OAI22_X1  g321(.A1(new_n504), .A2(new_n506), .B1(KEYINPUT15), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n507), .A2(KEYINPUT15), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n503), .A2(new_n235), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n509), .B1(new_n510), .B2(new_n505), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(G113), .B(G122), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(new_n379), .ZN(new_n514));
  INV_X1    g328(.A(G237), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n515), .A2(new_n188), .A3(G214), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n266), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n317), .A2(G143), .A3(G214), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g333(.A1(KEYINPUT18), .A2(G131), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT80), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT80), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n519), .A2(new_n523), .A3(new_n520), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n199), .B(new_n200), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n525), .B(new_n526), .C1(new_n519), .C2(new_n520), .ZN(new_n527));
  INV_X1    g341(.A(new_n518), .ZN(new_n528));
  AOI21_X1  g342(.A(G143), .B1(new_n317), .B2(G214), .ZN(new_n529));
  OAI21_X1  g343(.A(G131), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n517), .A2(new_n260), .A3(new_n518), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n519), .A2(KEYINPUT17), .A3(G131), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT81), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n225), .A2(new_n536), .A3(new_n226), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n536), .B1(new_n225), .B2(new_n226), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n514), .B(new_n527), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n514), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT19), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n199), .B(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n198), .B1(new_n543), .B2(G146), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n544), .B1(new_n530), .B2(new_n532), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n526), .B1(new_n519), .B2(new_n520), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n524), .B2(new_n522), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n541), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n540), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT82), .ZN(new_n550));
  AOI21_X1  g364(.A(KEYINPUT20), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(G475), .A2(G902), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n553), .B1(new_n540), .B2(new_n548), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n551), .B(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n527), .B1(new_n538), .B2(new_n539), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT83), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n556), .A2(new_n557), .A3(new_n541), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n557), .B1(new_n556), .B2(new_n541), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n540), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n235), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(G475), .ZN(new_n562));
  INV_X1    g376(.A(G952), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(G953), .ZN(new_n564));
  NAND2_X1  g378(.A1(G234), .A2(G237), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(G902), .A3(G953), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT21), .B(G898), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n567), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n512), .A2(new_n555), .A3(new_n562), .A4(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT87), .B1(new_n473), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n508), .A2(new_n572), .A3(new_n511), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n551), .A2(new_n554), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT20), .ZN(new_n577));
  AND4_X1   g391(.A1(KEYINPUT82), .A2(new_n549), .A3(new_n577), .A4(new_n552), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(G475), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n580), .B1(new_n560), .B2(new_n235), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n575), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT87), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n582), .A2(new_n583), .A3(new_n472), .A4(new_n430), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n574), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n374), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(G101), .ZN(G3));
  OAI21_X1  g401(.A(G472), .B1(new_n353), .B2(G902), .ZN(new_n588));
  INV_X1    g402(.A(new_n430), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n589), .A2(new_n247), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n349), .A2(new_n355), .A3(new_n588), .A4(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n555), .A2(new_n562), .ZN(new_n593));
  AOI211_X1 g407(.A(KEYINPUT88), .B(G478), .C1(new_n503), .C2(new_n235), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT88), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n595), .B1(new_n510), .B2(new_n507), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT33), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n503), .B(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n507), .A2(G902), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  OAI22_X1  g414(.A1(new_n594), .A2(new_n596), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n593), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(KEYINPUT89), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n472), .A2(new_n572), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n592), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT34), .B(G104), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G6));
  XOR2_X1   g422(.A(new_n571), .B(KEYINPUT91), .Z(new_n609));
  NAND2_X1  g423(.A1(new_n472), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n549), .ZN(new_n612));
  AOI211_X1 g426(.A(new_n553), .B(new_n612), .C1(KEYINPUT90), .C2(KEYINPUT20), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n614));
  NOR2_X1   g428(.A1(new_n554), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n562), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(new_n512), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n592), .A2(new_n611), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT35), .B(G107), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT92), .B(KEYINPUT93), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G9));
  NOR2_X1   g436(.A1(new_n219), .A2(new_n228), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n191), .A2(KEYINPUT36), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n623), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n245), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n243), .A2(KEYINPUT94), .A3(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT94), .ZN(new_n629));
  INV_X1    g443(.A(new_n242), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n630), .B1(new_n238), .B2(new_n239), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n626), .A2(new_n245), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n574), .A2(new_n634), .A3(new_n584), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n349), .A2(new_n355), .A3(new_n588), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT37), .B(G110), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT95), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n637), .B(new_n639), .ZN(G12));
  NAND3_X1  g454(.A1(new_n634), .A2(new_n472), .A3(new_n430), .ZN(new_n641));
  OR2_X1    g455(.A1(new_n568), .A2(G900), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n566), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n617), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n357), .A2(new_n373), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G128), .ZN(G30));
  INV_X1    g462(.A(new_n361), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n321), .ZN(new_n650));
  AOI21_X1  g464(.A(G902), .B1(new_n366), .B2(new_n339), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI22_X1  g466(.A1(new_n359), .A2(KEYINPUT32), .B1(new_n652), .B2(G472), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n357), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n643), .B(KEYINPUT39), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n430), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT96), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(KEYINPUT40), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT40), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n469), .A2(new_n471), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n662), .B(KEYINPUT38), .Z(new_n663));
  NOR2_X1   g477(.A1(new_n579), .A2(new_n581), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n631), .A2(new_n632), .ZN(new_n665));
  INV_X1    g479(.A(new_n512), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n665), .A2(new_n666), .A3(new_n431), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n663), .A2(new_n664), .A3(new_n667), .ZN(new_n668));
  AND4_X1   g482(.A1(new_n654), .A2(new_n659), .A3(new_n661), .A4(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT97), .B(G143), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G45));
  OAI211_X1 g485(.A(new_n601), .B(new_n643), .C1(new_n579), .C2(new_n581), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n641), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n646), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G146), .ZN(G48));
  NOR2_X1   g489(.A1(new_n424), .A2(new_n428), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(G902), .ZN(new_n677));
  INV_X1    g491(.A(G469), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n376), .B(new_n429), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n247), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n646), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n605), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT41), .B(G113), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G15));
  NOR3_X1   g498(.A1(new_n610), .A2(new_n512), .A3(new_n616), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G116), .ZN(G18));
  NAND3_X1  g501(.A1(new_n582), .A2(new_n628), .A3(new_n633), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n662), .A2(new_n431), .ZN(new_n689));
  OR3_X1    g503(.A1(new_n679), .A2(new_n689), .A3(KEYINPUT98), .ZN(new_n690));
  OAI21_X1  g504(.A(KEYINPUT98), .B1(new_n679), .B2(new_n689), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n688), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n646), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G119), .ZN(G21));
  OAI21_X1  g508(.A(new_n339), .B1(new_n367), .B2(new_n368), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n695), .B1(new_n341), .B2(new_n345), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n348), .ZN(new_n697));
  INV_X1    g511(.A(new_n247), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n588), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT99), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT99), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n588), .A2(new_n697), .A3(new_n701), .A4(new_n698), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n689), .A2(new_n664), .A3(new_n512), .ZN(new_n704));
  INV_X1    g518(.A(new_n679), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n704), .A2(new_n609), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G122), .ZN(G24));
  AOI21_X1  g522(.A(new_n672), .B1(new_n690), .B2(new_n691), .ZN(new_n709));
  INV_X1    g523(.A(new_n665), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n588), .A2(new_n697), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G125), .ZN(G27));
  NAND2_X1  g527(.A1(new_n359), .A2(KEYINPUT32), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n372), .A2(G472), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n356), .B1(new_n353), .B2(new_n354), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(G469), .A2(G902), .ZN(new_n718));
  XOR2_X1   g532(.A(new_n718), .B(KEYINPUT100), .Z(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n429), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n408), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n722), .A2(new_n396), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n416), .B1(new_n723), .B2(new_n407), .ZN(new_n724));
  INV_X1    g538(.A(new_n417), .ZN(new_n725));
  OAI21_X1  g539(.A(KEYINPUT101), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT101), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n413), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n726), .A2(G469), .A3(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT102), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n726), .A2(KEYINPUT102), .A3(G469), .A4(new_n728), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n721), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n469), .A2(new_n431), .A3(new_n471), .A4(new_n376), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n733), .A2(new_n672), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n717), .A2(new_n698), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(KEYINPUT42), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n733), .A2(new_n734), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n672), .A2(KEYINPUT42), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n646), .A2(new_n698), .A3(new_n738), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(new_n260), .ZN(G33));
  INV_X1    g556(.A(new_n644), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n646), .A2(new_n698), .A3(new_n743), .A4(new_n738), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT103), .B(G134), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G36));
  NAND2_X1  g560(.A1(new_n664), .A2(new_n601), .ZN(new_n747));
  XOR2_X1   g561(.A(new_n747), .B(KEYINPUT43), .Z(new_n748));
  NAND2_X1  g562(.A1(new_n636), .A2(new_n710), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n749), .A2(KEYINPUT104), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n749), .A2(KEYINPUT104), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n748), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n662), .A2(new_n432), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n752), .A2(new_n753), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT105), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n726), .A2(KEYINPUT45), .A3(new_n728), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n724), .A2(new_n725), .ZN(new_n761));
  OAI21_X1  g575(.A(G469), .B1(new_n761), .B2(KEYINPUT45), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n720), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT46), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI22_X1  g579(.A1(new_n763), .A2(new_n764), .B1(new_n677), .B2(new_n421), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n377), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n767), .A2(new_n655), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n754), .A2(KEYINPUT105), .A3(new_n755), .A4(new_n756), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n759), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  XOR2_X1   g584(.A(KEYINPUT106), .B(G137), .Z(new_n771));
  XNOR2_X1  g585(.A(new_n770), .B(new_n771), .ZN(G39));
  OR2_X1    g586(.A1(new_n767), .A2(KEYINPUT47), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n767), .A2(KEYINPUT47), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n755), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n776), .A2(new_n698), .A3(new_n672), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n775), .A2(new_n357), .A3(new_n373), .A4(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G140), .ZN(G42));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n780));
  AOI22_X1  g594(.A1(new_n374), .A2(new_n585), .B1(new_n646), .B2(new_n692), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n646), .B(new_n680), .C1(new_n605), .C2(new_n685), .ZN(new_n782));
  XOR2_X1   g596(.A(new_n602), .B(KEYINPUT108), .Z(new_n783));
  NAND3_X1  g597(.A1(new_n592), .A2(new_n611), .A3(new_n783), .ZN(new_n784));
  AND4_X1   g598(.A1(new_n707), .A2(new_n781), .A3(new_n782), .A4(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n593), .A2(new_n512), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n591), .A2(new_n610), .A3(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT109), .B1(new_n788), .B2(new_n637), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n349), .A2(new_n355), .A3(new_n588), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n790), .A2(new_n590), .A3(new_n611), .A4(new_n786), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT109), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n790), .A2(new_n585), .A3(new_n634), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n789), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n354), .B1(new_n358), .B2(new_n695), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n346), .A2(new_n235), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n796), .B1(new_n797), .B2(G472), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n798), .A2(KEYINPUT110), .A3(new_n710), .A4(new_n735), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n735), .A2(new_n588), .A3(new_n697), .A4(new_n710), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT110), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n628), .A2(new_n633), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n755), .A2(new_n512), .A3(new_n643), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n804), .A2(new_n805), .A3(new_n589), .A4(new_n616), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n646), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n744), .A2(new_n803), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n741), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n785), .A2(new_n795), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n704), .ZN(new_n811));
  INV_X1    g625(.A(new_n733), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n643), .A2(new_n376), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n812), .A2(KEYINPUT111), .A3(new_n665), .A4(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT111), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n665), .A2(new_n813), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n815), .B1(new_n816), .B2(new_n733), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n811), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n654), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n647), .A2(new_n674), .A3(new_n819), .A4(new_n712), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT52), .ZN(new_n821));
  AOI22_X1  g635(.A1(new_n645), .A2(new_n646), .B1(new_n709), .B2(new_n711), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n822), .A2(new_n823), .A3(new_n674), .A4(new_n819), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n780), .B1(new_n810), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT114), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n781), .A2(new_n707), .A3(new_n782), .A4(new_n784), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n789), .A2(new_n794), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n809), .A3(new_n824), .A4(new_n821), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(KEYINPUT114), .A3(new_n780), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n822), .A2(KEYINPUT112), .A3(new_n674), .A4(new_n819), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n821), .A2(new_n824), .A3(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(KEYINPUT112), .B(KEYINPUT113), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n836), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n821), .A2(new_n824), .A3(new_n834), .A4(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n810), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n828), .A2(new_n833), .B1(new_n840), .B2(KEYINPUT53), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n748), .A2(new_n567), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n844), .A2(new_n705), .A3(new_n755), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n247), .B1(new_n373), .B2(new_n716), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n848), .A2(KEYINPUT48), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n848), .A2(KEYINPUT48), .ZN(new_n850));
  OR3_X1    g664(.A1(new_n847), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n844), .A2(new_n703), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n690), .A2(new_n691), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n603), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n698), .A2(new_n705), .A3(new_n567), .A4(new_n755), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n654), .A2(new_n856), .ZN(new_n857));
  AOI22_X1  g671(.A1(new_n847), .A2(new_n850), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n851), .A2(new_n564), .A3(new_n854), .A4(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n852), .A2(new_n755), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT115), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n429), .B1(new_n677), .B2(new_n678), .ZN(new_n862));
  OAI22_X1  g676(.A1(new_n775), .A2(new_n861), .B1(new_n376), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT115), .B1(new_n773), .B2(new_n774), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n860), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n663), .A2(new_n705), .A3(new_n432), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n844), .A2(new_n703), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT50), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n867), .A2(new_n868), .ZN(new_n870));
  OAI22_X1  g684(.A1(new_n869), .A2(new_n870), .B1(KEYINPUT116), .B2(KEYINPUT51), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n867), .B(new_n868), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n865), .B(new_n871), .C1(KEYINPUT116), .C2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT117), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT51), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n593), .A2(new_n601), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n845), .A2(new_n711), .B1(new_n857), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n862), .A2(new_n376), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n860), .B1(new_n775), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n881), .B1(new_n878), .B2(new_n874), .ZN(new_n882));
  INV_X1    g696(.A(new_n872), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT51), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n859), .B1(new_n879), .B2(new_n884), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n832), .A2(new_n780), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n886), .B1(new_n840), .B2(KEYINPUT53), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT54), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n843), .A2(new_n885), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n563), .A2(new_n188), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR4_X1   g705(.A1(new_n747), .A2(new_n247), .A3(new_n432), .A4(new_n377), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n862), .A2(KEYINPUT49), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT107), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n663), .B1(KEYINPUT49), .B2(new_n862), .ZN(new_n896));
  OR3_X1    g710(.A1(new_n895), .A2(new_n654), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n891), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT119), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT119), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n891), .A2(new_n900), .A3(new_n897), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n901), .ZN(G75));
  NOR2_X1   g716(.A1(new_n841), .A2(new_n235), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n468), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT56), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n460), .A2(new_n463), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(new_n461), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT55), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n904), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n908), .B1(new_n904), .B2(new_n905), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n188), .A2(G952), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(G51));
  XNOR2_X1  g726(.A(new_n841), .B(KEYINPUT54), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n719), .B(KEYINPUT57), .Z(new_n914));
  OAI22_X1  g728(.A1(new_n913), .A2(new_n914), .B1(new_n424), .B2(new_n428), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n760), .A2(new_n762), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n903), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n911), .B1(new_n915), .B2(new_n917), .ZN(G54));
  NAND3_X1  g732(.A1(new_n903), .A2(KEYINPUT58), .A3(G475), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n919), .A2(new_n612), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n919), .A2(new_n612), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n920), .A2(new_n921), .A3(new_n911), .ZN(G60));
  INV_X1    g736(.A(new_n911), .ZN(new_n923));
  INV_X1    g737(.A(new_n598), .ZN(new_n924));
  NAND2_X1  g738(.A1(G478), .A2(G902), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT59), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n923), .B1(new_n913), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n843), .A2(new_n888), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n924), .B1(new_n929), .B2(new_n926), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n928), .A2(new_n930), .ZN(G63));
  NAND2_X1  g745(.A1(new_n837), .A2(new_n839), .ZN(new_n932));
  INV_X1    g746(.A(new_n810), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n932), .A2(KEYINPUT53), .A3(new_n933), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n832), .A2(KEYINPUT114), .A3(new_n780), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT114), .B1(new_n832), .B2(new_n780), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(G217), .A2(G902), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT60), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n937), .A2(new_n626), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(KEYINPUT120), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT61), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT121), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n828), .A2(new_n833), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n939), .B1(new_n946), .B2(new_n934), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n911), .B1(new_n947), .B2(new_n626), .ZN(new_n948));
  INV_X1    g762(.A(new_n244), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(new_n841), .B2(new_n939), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n945), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  AND4_X1   g765(.A1(new_n945), .A2(new_n950), .A3(new_n923), .A4(new_n941), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n944), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n950), .A2(new_n941), .A3(new_n923), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(KEYINPUT121), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n948), .A2(new_n945), .A3(new_n950), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n955), .A2(new_n956), .A3(new_n943), .A4(new_n942), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n953), .A2(new_n957), .ZN(G66));
  NOR2_X1   g772(.A1(new_n831), .A2(G953), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT122), .ZN(new_n960));
  OAI21_X1  g774(.A(G953), .B1(new_n570), .B2(new_n436), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n906), .B1(G898), .B2(new_n188), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT123), .Z(new_n964));
  XNOR2_X1  g778(.A(new_n962), .B(new_n964), .ZN(G69));
  AOI21_X1  g779(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(KEYINPUT126), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n658), .A2(new_n776), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n968), .B(new_n374), .C1(new_n783), .C2(new_n786), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT124), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n822), .A2(new_n674), .ZN(new_n971));
  OAI21_X1  g785(.A(KEYINPUT62), .B1(new_n971), .B2(new_n669), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n970), .A2(new_n778), .A3(new_n972), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n971), .A2(new_n669), .A3(KEYINPUT62), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(G953), .B1(new_n770), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n330), .A2(new_n331), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(new_n543), .Z(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n967), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n768), .A2(new_n704), .A3(new_n846), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n778), .A2(new_n744), .A3(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n982), .A2(new_n741), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT125), .ZN(new_n984));
  INV_X1    g798(.A(new_n971), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n770), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n984), .B1(new_n770), .B2(new_n985), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n188), .B(new_n983), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n978), .B1(G900), .B2(G953), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n980), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n966), .A2(KEYINPUT126), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  AOI211_X1 g808(.A(new_n992), .B(new_n980), .C1(new_n989), .C2(new_n990), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n994), .A2(new_n995), .ZN(G72));
  OAI211_X1 g810(.A(new_n831), .B(new_n983), .C1(new_n987), .C2(new_n988), .ZN(new_n997));
  NAND2_X1  g811(.A1(G472), .A2(G902), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT63), .Z(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT127), .Z(new_n1000));
  AOI211_X1 g814(.A(new_n321), .B(new_n649), .C1(new_n997), .C2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n350), .B1(new_n361), .B2(new_n321), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n887), .A2(new_n999), .A3(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n770), .A2(new_n831), .A3(new_n975), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n1004), .A2(new_n1000), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n923), .B(new_n1003), .C1(new_n1005), .C2(new_n650), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n1001), .A2(new_n1006), .ZN(G57));
endmodule


