//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0 1 0 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n988,
    new_n989, new_n990;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT25), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT65), .ZN(new_n205));
  OAI211_X1 g004(.A(G183gat), .B(G190gat), .C1(new_n205), .C2(KEYINPUT24), .ZN(new_n206));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT24), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n207), .A2(KEYINPUT65), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT67), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G190gat), .ZN(new_n213));
  INV_X1    g012(.A(G183gat), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G190gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT66), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G190gat), .ZN(new_n219));
  AND4_X1   g018(.A1(new_n212), .A2(new_n217), .A3(new_n219), .A4(new_n214), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n211), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT23), .ZN(new_n223));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G169gat), .B2(G176gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n223), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n204), .B1(new_n221), .B2(new_n228), .ZN(new_n229));
  AND4_X1   g028(.A1(new_n204), .A2(new_n223), .A3(new_n226), .A4(new_n224), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n207), .A2(new_n208), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT64), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n207), .A2(new_n233), .A3(new_n208), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n214), .A2(new_n216), .ZN(new_n235));
  NAND3_X1  g034(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n232), .A2(new_n234), .A3(new_n235), .A4(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n230), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT28), .ZN(new_n239));
  NAND2_X1  g038(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT27), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT27), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(KEYINPUT68), .A3(G183gat), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n241), .A2(new_n243), .A3(new_n217), .A4(new_n219), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n217), .A2(new_n219), .A3(KEYINPUT28), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT27), .B(G183gat), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n239), .A2(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n222), .A2(KEYINPUT26), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n207), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT26), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n224), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n251), .A2(new_n222), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n238), .B1(new_n247), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n229), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n203), .B1(new_n256), .B2(KEYINPUT29), .ZN(new_n257));
  XNOR2_X1  g056(.A(G197gat), .B(G204gat), .ZN(new_n258));
  INV_X1    g057(.A(G211gat), .ZN(new_n259));
  INV_X1    g058(.A(G218gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n258), .B1(KEYINPUT22), .B2(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(G211gat), .B(G218gat), .Z(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  NOR3_X1   g063(.A1(new_n256), .A2(KEYINPUT74), .A3(new_n203), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n244), .A2(new_n239), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n213), .A2(new_n246), .A3(KEYINPUT28), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI22_X1  g067(.A1(new_n268), .A2(new_n253), .B1(new_n237), .B2(new_n230), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n217), .A2(new_n219), .A3(new_n214), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT67), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n213), .A2(new_n212), .A3(new_n214), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n210), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT25), .B1(new_n273), .B2(new_n227), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n203), .B1(new_n269), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT74), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n257), .B(new_n264), .C1(new_n265), .C2(new_n277), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n262), .A2(new_n263), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n262), .A2(new_n263), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n269), .A2(new_n274), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT73), .B(KEYINPUT29), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n282), .A2(new_n283), .B1(G226gat), .B2(G233gat), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n281), .B1(new_n284), .B2(new_n275), .ZN(new_n285));
  XNOR2_X1  g084(.A(G8gat), .B(G36gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(G64gat), .B(G92gat), .ZN(new_n287));
  XOR2_X1   g086(.A(new_n286), .B(new_n287), .Z(new_n288));
  AND3_X1   g087(.A1(new_n278), .A2(new_n285), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n288), .B1(new_n278), .B2(new_n285), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT30), .ZN(new_n291));
  OR3_X1    g090(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n278), .A2(new_n285), .ZN(new_n293));
  INV_X1    g092(.A(new_n288), .ZN(new_n294));
  NOR3_X1   g093(.A1(new_n293), .A2(KEYINPUT30), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G1gat), .B(G29gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n298), .B(KEYINPUT0), .ZN(new_n299));
  XNOR2_X1  g098(.A(G57gat), .B(G85gat), .ZN(new_n300));
  XOR2_X1   g099(.A(new_n299), .B(new_n300), .Z(new_n301));
  INV_X1    g100(.A(G113gat), .ZN(new_n302));
  INV_X1    g101(.A(G120gat), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT1), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G113gat), .A2(G120gat), .ZN(new_n305));
  INV_X1    g104(.A(G134gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G127gat), .ZN(new_n307));
  INV_X1    g106(.A(G127gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G134gat), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n304), .A2(new_n305), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n302), .A2(new_n303), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT70), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT1), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n311), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n307), .A2(new_n309), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT69), .B(G113gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G120gat), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n310), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G141gat), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT78), .B1(new_n322), .B2(G148gat), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT78), .ZN(new_n324));
  INV_X1    g123(.A(G148gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(new_n325), .A3(G141gat), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n322), .A2(KEYINPUT77), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT77), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G141gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(new_n330), .A3(G148gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(G162gat), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT2), .B1(new_n333), .B2(KEYINPUT79), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(G155gat), .ZN(new_n335));
  INV_X1    g134(.A(G155gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G162gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n334), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n332), .A2(new_n339), .ZN(new_n340));
  OR2_X1    g139(.A1(KEYINPUT75), .A2(KEYINPUT2), .ZN(new_n341));
  NAND2_X1  g140(.A1(KEYINPUT75), .A2(KEYINPUT2), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n322), .A2(G148gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n325), .A2(G141gat), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n341), .B(new_n342), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n335), .A2(new_n337), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT76), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G141gat), .B(G148gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT75), .B(KEYINPUT2), .ZN(new_n349));
  OAI211_X1 g148(.A(KEYINPUT76), .B(new_n346), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n321), .B(new_n340), .C1(new_n347), .C2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT4), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n338), .B1(new_n327), .B2(new_n331), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n346), .B1(new_n348), .B2(new_n349), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT76), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n355), .B1(new_n358), .B2(new_n350), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n359), .A2(KEYINPUT4), .A3(new_n321), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n354), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT5), .ZN(new_n362));
  NAND2_X1  g161(.A1(G225gat), .A2(G233gat), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n340), .B1(new_n351), .B2(new_n347), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT3), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT3), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n359), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n321), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n365), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n361), .A2(new_n362), .A3(new_n363), .A4(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n363), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n358), .A2(new_n350), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n372), .A2(new_n340), .A3(new_n321), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n321), .B1(new_n372), .B2(new_n340), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n371), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT81), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT82), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT81), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n378), .B(new_n371), .C1(new_n373), .C2(new_n374), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT5), .A4(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT80), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n368), .B1(new_n359), .B2(new_n366), .ZN(new_n382));
  AOI211_X1 g181(.A(KEYINPUT3), .B(new_n355), .C1(new_n358), .C2(new_n350), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n354), .B(new_n360), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n381), .B1(new_n384), .B2(new_n371), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n361), .A2(KEYINPUT80), .A3(new_n363), .A4(new_n369), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n380), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n362), .B1(new_n375), .B2(KEYINPUT81), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n377), .B1(new_n388), .B2(new_n379), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n301), .B(new_n370), .C1(new_n387), .C2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT6), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n364), .A2(new_n368), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n363), .B1(new_n393), .B2(new_n352), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT5), .B1(new_n394), .B2(new_n378), .ZN(new_n395));
  INV_X1    g194(.A(new_n379), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT82), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n397), .A2(new_n380), .A3(new_n385), .A4(new_n386), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n301), .B1(new_n398), .B2(new_n370), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n392), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n370), .B1(new_n387), .B2(new_n389), .ZN(new_n401));
  INV_X1    g200(.A(new_n301), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(KEYINPUT6), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n297), .B1(new_n400), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n368), .B1(new_n229), .B2(new_n255), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT72), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n282), .A2(KEYINPUT72), .A3(new_n368), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n269), .A2(new_n274), .A3(new_n321), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT71), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n269), .A2(new_n274), .A3(KEYINPUT71), .A4(new_n321), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(G227gat), .A2(G233gat), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT34), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n408), .A2(new_n409), .B1(new_n413), .B2(new_n414), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT34), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(new_n421), .A3(new_n417), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT33), .B1(new_n416), .B2(new_n418), .ZN(new_n423));
  XOR2_X1   g222(.A(G15gat), .B(G43gat), .Z(new_n424));
  XNOR2_X1  g223(.A(G71gat), .B(G99gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n419), .B(new_n422), .C1(new_n423), .C2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT33), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n429), .B1(new_n420), .B2(new_n417), .ZN(new_n430));
  AND4_X1   g229(.A1(new_n421), .A2(new_n410), .A3(new_n417), .A4(new_n415), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n421), .B1(new_n420), .B2(new_n417), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n430), .B(new_n426), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n416), .A2(new_n418), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT32), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT31), .B(G50gat), .ZN(new_n438));
  INV_X1    g237(.A(G106gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G228gat), .A2(G233gat), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n264), .B1(new_n367), .B2(new_n283), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n264), .A2(new_n283), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n359), .B1(new_n444), .B2(new_n366), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n442), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n366), .B1(new_n281), .B2(KEYINPUT29), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n442), .B1(new_n447), .B2(new_n364), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n448), .B1(new_n443), .B2(KEYINPUT83), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT83), .ZN(new_n450));
  AOI211_X1 g249(.A(new_n450), .B(new_n264), .C1(new_n367), .C2(new_n283), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n446), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(G22gat), .ZN(new_n453));
  INV_X1    g252(.A(G78gat), .ZN(new_n454));
  INV_X1    g253(.A(G22gat), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n446), .B(new_n455), .C1(new_n449), .C2(new_n451), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n453), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n454), .B1(new_n453), .B2(new_n456), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n441), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n453), .A2(new_n456), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(G78gat), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n453), .A2(new_n454), .A3(new_n456), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n462), .A3(new_n440), .ZN(new_n463));
  INV_X1    g262(.A(new_n436), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n428), .A2(new_n433), .A3(new_n464), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n437), .A2(new_n459), .A3(new_n463), .A4(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n202), .B1(new_n405), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n466), .ZN(new_n468));
  NOR3_X1   g267(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n469), .A2(new_n295), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n401), .A2(new_n402), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n471), .A2(new_n391), .A3(new_n390), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n470), .B1(new_n472), .B2(new_n403), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n468), .A2(KEYINPUT35), .A3(new_n473), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n459), .A2(new_n463), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT39), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT84), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n384), .A2(new_n477), .A3(new_n371), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n477), .B1(new_n384), .B2(new_n371), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n384), .A2(new_n371), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT84), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n384), .A2(new_n477), .A3(new_n371), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n373), .A2(new_n374), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n476), .B1(new_n484), .B2(new_n363), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n480), .A2(new_n486), .A3(new_n301), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT40), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n480), .A2(new_n486), .A3(KEYINPUT40), .A4(new_n301), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n471), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT85), .B1(new_n491), .B2(new_n297), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n293), .A2(KEYINPUT37), .ZN(new_n493));
  XNOR2_X1  g292(.A(KEYINPUT87), .B(KEYINPUT37), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n278), .A2(new_n285), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n294), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT38), .B1(new_n493), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n257), .B1(new_n265), .B2(new_n277), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT86), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(new_n499), .A3(new_n281), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n498), .A2(new_n281), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n284), .A2(new_n275), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT86), .B1(new_n502), .B2(new_n281), .ZN(new_n503));
  OAI211_X1 g302(.A(KEYINPUT37), .B(new_n500), .C1(new_n501), .C2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT38), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n495), .A2(new_n505), .A3(new_n294), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n289), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n472), .A2(new_n403), .A3(new_n497), .A4(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n490), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n509), .A2(new_n399), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT85), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n510), .A2(new_n511), .A3(new_n470), .A4(new_n489), .ZN(new_n512));
  AND4_X1   g311(.A1(new_n475), .A2(new_n492), .A3(new_n508), .A4(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n437), .A2(KEYINPUT36), .A3(new_n465), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(KEYINPUT36), .B1(new_n437), .B2(new_n465), .ZN(new_n516));
  OAI22_X1  g315(.A1(new_n515), .A2(new_n516), .B1(new_n473), .B2(new_n475), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n467), .B(new_n474), .C1(new_n513), .C2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G15gat), .B(G22gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(KEYINPUT93), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT16), .ZN(new_n521));
  OR2_X1    g320(.A1(new_n521), .A2(G1gat), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n520), .A2(G1gat), .ZN(new_n524));
  OAI21_X1  g323(.A(G8gat), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n520), .B1(new_n521), .B2(G1gat), .ZN(new_n526));
  INV_X1    g325(.A(G8gat), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n526), .B(new_n527), .C1(G1gat), .C2(new_n520), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(G50gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(G43gat), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT15), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n530), .A2(G43gat), .ZN(new_n534));
  NOR3_X1   g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(G29gat), .ZN(new_n536));
  INV_X1    g335(.A(G36gat), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n536), .A2(new_n537), .A3(KEYINPUT14), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT14), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n539), .B1(G29gat), .B2(G36gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n536), .A2(new_n537), .ZN(new_n542));
  NOR3_X1   g341(.A1(new_n535), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT91), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n534), .B1(new_n544), .B2(new_n531), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n532), .A2(KEYINPUT91), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(new_n533), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT89), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n541), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n538), .A2(new_n540), .A3(KEYINPUT89), .ZN(new_n552));
  INV_X1    g351(.A(new_n542), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(KEYINPUT90), .A3(new_n535), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT90), .B1(new_n554), .B2(new_n535), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n549), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n529), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n529), .A2(new_n558), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G229gat), .A2(G233gat), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n563), .B(KEYINPUT13), .Z(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT17), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT94), .B1(new_n558), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n554), .A2(new_n535), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT90), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(new_n555), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT94), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n572), .A2(new_n573), .A3(KEYINPUT17), .A4(new_n549), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n568), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n529), .ZN(new_n576));
  XOR2_X1   g375(.A(KEYINPUT92), .B(KEYINPUT17), .Z(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n558), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n575), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n580), .A2(new_n563), .A3(new_n559), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT18), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n566), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n580), .A2(KEYINPUT18), .A3(new_n563), .A4(new_n559), .ZN(new_n584));
  XNOR2_X1  g383(.A(G113gat), .B(G141gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G169gat), .B(G197gat), .Z(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT12), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n583), .A2(new_n584), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n590), .B1(new_n583), .B2(new_n584), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n518), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G85gat), .A2(G92gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT7), .ZN(new_n597));
  NAND2_X1  g396(.A1(G99gat), .A2(G106gat), .ZN(new_n598));
  INV_X1    g397(.A(G85gat), .ZN(new_n599));
  INV_X1    g398(.A(G92gat), .ZN(new_n600));
  AOI22_X1  g399(.A1(KEYINPUT8), .A2(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G99gat), .B(G106gat), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT97), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n604), .B(KEYINPUT97), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(new_n602), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT98), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n607), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n603), .A2(new_n606), .A3(KEYINPUT98), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n558), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g413(.A1(G232gat), .A2(G233gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT41), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G190gat), .B(G218gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n568), .A2(new_n574), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n613), .A2(KEYINPUT99), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT99), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n611), .A2(new_n623), .A3(new_n612), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n579), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n618), .B(new_n620), .C1(new_n621), .C2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT100), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n579), .A2(new_n624), .A3(new_n622), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n617), .B1(new_n629), .B2(new_n575), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n630), .A2(KEYINPUT100), .A3(new_n620), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(G134gat), .B(G162gat), .Z(new_n633));
  NOR2_X1   g432(.A1(new_n615), .A2(KEYINPUT41), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n630), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n635), .B1(new_n636), .B2(new_n619), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n632), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT102), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n632), .A2(KEYINPUT102), .A3(new_n637), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT101), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n626), .A2(new_n627), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT100), .B1(new_n630), .B2(new_n620), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n628), .A2(KEYINPUT101), .A3(new_n631), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n636), .A2(new_n619), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n635), .ZN(new_n650));
  XOR2_X1   g449(.A(G57gat), .B(G64gat), .Z(new_n651));
  INV_X1    g450(.A(KEYINPUT9), .ZN(new_n652));
  INV_X1    g451(.A(G71gat), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n652), .B1(new_n653), .B2(new_n454), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G71gat), .B(G78gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n657), .A2(KEYINPUT21), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT95), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n529), .B1(KEYINPUT21), .B2(new_n657), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT96), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n662), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(G127gat), .B(G155gat), .ZN(new_n668));
  NAND2_X1  g467(.A1(G231gat), .A2(G233gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(G183gat), .B(G211gat), .Z(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n665), .A2(new_n666), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n661), .ZN(new_n674));
  AND3_X1   g473(.A1(new_n667), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n672), .B1(new_n667), .B2(new_n674), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n657), .A2(KEYINPUT10), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n613), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(KEYINPUT103), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT10), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n657), .A2(new_n607), .A3(new_n609), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n681), .B(new_n682), .C1(new_n613), .C2(new_n657), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n613), .A2(new_n678), .A3(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n680), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(G230gat), .A2(G233gat), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n682), .B1(new_n613), .B2(new_n657), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n689), .A2(G230gat), .A3(G233gat), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(G120gat), .B(G148gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(G176gat), .B(G204gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT104), .B(KEYINPUT105), .Z(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n691), .A2(new_n696), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n642), .A2(new_n650), .A3(new_n677), .A4(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT106), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI22_X1  g502(.A1(new_n640), .A2(new_n641), .B1(new_n649), .B2(new_n635), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n704), .A2(KEYINPUT106), .A3(new_n677), .A4(new_n700), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n595), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n472), .A2(new_n403), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g509(.A1(new_n707), .A2(new_n297), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT16), .B(G8gat), .Z(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n713), .B1(new_n527), .B2(new_n711), .ZN(new_n714));
  MUX2_X1   g513(.A(new_n713), .B(new_n714), .S(KEYINPUT42), .Z(G1325gat));
  NOR2_X1   g514(.A1(new_n515), .A2(new_n516), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(G15gat), .B1(new_n707), .B2(new_n717), .ZN(new_n718));
  AND3_X1   g517(.A1(new_n428), .A2(new_n433), .A3(new_n464), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n464), .B1(new_n428), .B2(new_n433), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  OR2_X1    g521(.A1(new_n722), .A2(G15gat), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n718), .B1(new_n707), .B2(new_n723), .ZN(G1326gat));
  NAND2_X1  g523(.A1(new_n459), .A2(new_n463), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n595), .A2(new_n725), .A3(new_n706), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT107), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT43), .B(G22gat), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1327gat));
  NOR3_X1   g528(.A1(new_n704), .A2(new_n677), .A3(new_n699), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n595), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n708), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n732), .A2(new_n536), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT45), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n474), .A2(new_n467), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT36), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n719), .B2(new_n720), .ZN(new_n739));
  AOI22_X1  g538(.A1(new_n405), .A2(new_n725), .B1(new_n739), .B2(new_n514), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n492), .A2(new_n508), .A3(new_n512), .A4(new_n475), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n740), .A2(KEYINPUT108), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT108), .B1(new_n740), .B2(new_n741), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n737), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n642), .A2(new_n650), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT44), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n518), .A2(KEYINPUT44), .A3(new_n745), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n593), .A2(new_n677), .A3(new_n699), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G29gat), .B1(new_n750), .B2(new_n708), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n751), .ZN(G1328gat));
  NOR3_X1   g551(.A1(new_n731), .A2(G36gat), .A3(new_n297), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT46), .ZN(new_n754));
  OAI21_X1  g553(.A(G36gat), .B1(new_n750), .B2(new_n297), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(G1329gat));
  AOI21_X1  g555(.A(G43gat), .B1(new_n732), .B2(new_n721), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n757), .B1(KEYINPUT109), .B2(KEYINPUT47), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n716), .A2(G43gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n758), .B1(new_n750), .B2(new_n759), .ZN(new_n760));
  OR2_X1    g559(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n760), .B(new_n761), .ZN(G1330gat));
  OAI21_X1  g561(.A(G50gat), .B1(new_n750), .B2(new_n475), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT110), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT48), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n732), .A2(new_n530), .A3(new_n725), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n765), .B(new_n767), .ZN(G1331gat));
  INV_X1    g567(.A(new_n677), .ZN(new_n769));
  NOR4_X1   g568(.A1(new_n745), .A2(new_n594), .A3(new_n769), .A4(new_n700), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n744), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n733), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g573(.A1(new_n771), .A2(new_n297), .ZN(new_n775));
  NOR2_X1   g574(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n776));
  AND2_X1   g575(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n775), .B2(new_n776), .ZN(G1333gat));
  OAI21_X1  g578(.A(G71gat), .B1(new_n771), .B2(new_n717), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n721), .A2(new_n653), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n780), .B1(new_n771), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g581(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n782), .B(new_n783), .ZN(G1334gat));
  NOR2_X1   g583(.A1(new_n771), .A2(new_n475), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(new_n454), .ZN(G1335gat));
  NOR2_X1   g585(.A1(new_n594), .A2(new_n677), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n700), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n746), .A2(new_n747), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(G85gat), .B1(new_n792), .B2(new_n708), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n744), .A2(new_n794), .A3(new_n745), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n787), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n794), .B1(new_n744), .B2(new_n745), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n798), .B(new_n799), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n800), .A2(new_n700), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n733), .A2(new_n599), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n793), .B1(new_n801), .B2(new_n802), .ZN(G1336gat));
  AOI21_X1  g602(.A(new_n600), .B1(new_n791), .B2(new_n470), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n804), .A2(KEYINPUT52), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n470), .A2(new_n699), .A3(new_n600), .ZN(new_n806));
  XOR2_X1   g605(.A(new_n806), .B(KEYINPUT113), .Z(new_n807));
  OAI21_X1  g606(.A(new_n805), .B1(new_n800), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n799), .A2(KEYINPUT114), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n810), .B1(new_n796), .B2(new_n797), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT108), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n812), .B1(new_n513), .B2(new_n517), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n740), .A2(KEYINPUT108), .A3(new_n741), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n736), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT112), .B1(new_n815), .B2(new_n704), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n816), .A2(new_n795), .A3(new_n787), .A4(new_n809), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n807), .B1(new_n811), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT52), .B1(new_n818), .B2(new_n804), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n808), .A2(new_n819), .ZN(G1337gat));
  OR2_X1    g619(.A1(new_n722), .A2(G99gat), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n792), .A2(KEYINPUT115), .A3(new_n717), .ZN(new_n822));
  OAI21_X1  g621(.A(KEYINPUT115), .B1(new_n792), .B2(new_n717), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G99gat), .ZN(new_n824));
  OAI22_X1  g623(.A1(new_n801), .A2(new_n821), .B1(new_n822), .B2(new_n824), .ZN(G1338gat));
  AOI21_X1  g624(.A(new_n439), .B1(new_n791), .B2(new_n725), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n826), .A2(KEYINPUT53), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n475), .A2(G106gat), .A3(new_n700), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n827), .B1(new_n800), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n813), .A2(new_n814), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n704), .B1(new_n831), .B2(new_n737), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n788), .B1(new_n832), .B2(new_n794), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n809), .B1(new_n833), .B2(new_n816), .ZN(new_n834));
  INV_X1    g633(.A(new_n817), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n828), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n826), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT116), .B1(new_n838), .B2(KEYINPUT53), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n829), .B1(new_n811), .B2(new_n817), .ZN(new_n840));
  OAI211_X1 g639(.A(KEYINPUT116), .B(KEYINPUT53), .C1(new_n840), .C2(new_n826), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n830), .B1(new_n839), .B2(new_n842), .ZN(G1339gat));
  NOR2_X1   g642(.A1(new_n708), .A2(new_n470), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n721), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT55), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n686), .A2(new_n687), .ZN(new_n847));
  AND3_X1   g646(.A1(new_n847), .A2(new_n688), .A3(KEYINPUT54), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n696), .B1(new_n688), .B2(KEYINPUT54), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n846), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n847), .A2(new_n688), .A3(KEYINPUT54), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n688), .A2(KEYINPUT54), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n851), .A2(new_n852), .A3(KEYINPUT55), .A4(new_n696), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n850), .A2(new_n697), .A3(new_n853), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n560), .A2(new_n561), .A3(new_n564), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT117), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n563), .B1(new_n580), .B2(new_n559), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n589), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n583), .A2(new_n584), .A3(new_n590), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI22_X1  g659(.A1(new_n593), .A2(new_n854), .B1(new_n860), .B2(new_n700), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n704), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n854), .A2(new_n860), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n745), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n677), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  NOR4_X1   g664(.A1(new_n745), .A2(new_n594), .A3(new_n769), .A4(new_n699), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(KEYINPUT118), .A3(new_n475), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n865), .A2(new_n866), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n869), .B1(new_n870), .B2(new_n725), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n845), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n302), .B1(new_n872), .B2(new_n594), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n870), .A2(new_n708), .A3(new_n470), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n468), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n875), .A2(new_n319), .A3(new_n593), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n873), .A2(new_n876), .ZN(G1340gat));
  AOI21_X1  g676(.A(new_n303), .B1(new_n872), .B2(new_n699), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n875), .A2(G120gat), .A3(new_n700), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g679(.A(new_n880), .B(KEYINPUT119), .Z(G1341gat));
  INV_X1    g680(.A(new_n872), .ZN(new_n882));
  OAI21_X1  g681(.A(G127gat), .B1(new_n882), .B2(new_n769), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n677), .A2(new_n308), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n883), .B1(new_n875), .B2(new_n884), .ZN(G1342gat));
  NAND4_X1  g684(.A1(new_n874), .A2(new_n306), .A3(new_n468), .A4(new_n745), .ZN(new_n886));
  XOR2_X1   g685(.A(new_n886), .B(KEYINPUT56), .Z(new_n887));
  OAI21_X1  g686(.A(G134gat), .B1(new_n882), .B2(new_n704), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1343gat));
  NAND2_X1  g688(.A1(new_n867), .A2(new_n725), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n717), .A2(new_n844), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n322), .A3(new_n594), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n890), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n867), .A2(KEYINPUT57), .A3(new_n725), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XOR2_X1   g699(.A(new_n892), .B(KEYINPUT120), .Z(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n902), .A2(new_n593), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n328), .A2(new_n330), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n896), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT58), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT58), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n907), .B(new_n896), .C1(new_n903), .C2(new_n904), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(G1344gat));
  NAND3_X1  g708(.A1(new_n895), .A2(new_n325), .A3(new_n699), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n911));
  INV_X1    g710(.A(new_n899), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n594), .B1(new_n703), .B2(new_n705), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n914), .B2(new_n865), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n725), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n914), .A2(new_n865), .A3(new_n913), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n897), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n912), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI211_X1 g719(.A(KEYINPUT122), .B(new_n897), .C1(new_n916), .C2(new_n917), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n901), .A2(new_n699), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n911), .B1(new_n924), .B2(G148gat), .ZN(new_n925));
  INV_X1    g724(.A(new_n902), .ZN(new_n926));
  AOI211_X1 g725(.A(KEYINPUT59), .B(new_n325), .C1(new_n926), .C2(new_n699), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n910), .B1(new_n925), .B2(new_n927), .ZN(G1345gat));
  NOR3_X1   g727(.A1(new_n902), .A2(new_n336), .A3(new_n769), .ZN(new_n929));
  OAI21_X1  g728(.A(KEYINPUT123), .B1(new_n894), .B2(new_n769), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n894), .A2(KEYINPUT123), .A3(new_n769), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n931), .A2(G155gat), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n929), .B1(new_n930), .B2(new_n932), .ZN(G1346gat));
  XOR2_X1   g732(.A(KEYINPUT79), .B(G162gat), .Z(new_n934));
  AND4_X1   g733(.A1(new_n745), .A2(new_n900), .A3(new_n901), .A4(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n895), .B2(new_n745), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT124), .ZN(G1347gat));
  NOR2_X1   g737(.A1(new_n870), .A2(new_n733), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n939), .A2(new_n470), .A3(new_n468), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(G169gat), .B1(new_n941), .B2(new_n594), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n733), .A2(new_n297), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(new_n721), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n944), .B1(new_n868), .B2(new_n871), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n594), .A2(G169gat), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n942), .B1(new_n945), .B2(new_n946), .ZN(G1348gat));
  INV_X1    g746(.A(G176gat), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n941), .A2(new_n948), .A3(new_n699), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n945), .A2(new_n699), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n950), .B2(new_n948), .ZN(G1349gat));
  AOI21_X1  g750(.A(new_n214), .B1(new_n945), .B2(new_n677), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n677), .A2(new_n246), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n952), .B1(new_n941), .B2(new_n953), .ZN(new_n954));
  XOR2_X1   g753(.A(new_n954), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g754(.A1(new_n941), .A2(new_n213), .A3(new_n745), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n945), .A2(new_n745), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n958), .B2(G190gat), .ZN(new_n959));
  AOI211_X1 g758(.A(KEYINPUT61), .B(new_n216), .C1(new_n945), .C2(new_n745), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT125), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI211_X1 g762(.A(KEYINPUT125), .B(new_n956), .C1(new_n959), .C2(new_n960), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1351gat));
  NOR3_X1   g764(.A1(new_n716), .A2(new_n297), .A3(new_n475), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n939), .A2(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(G197gat), .B1(new_n968), .B2(new_n594), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n717), .A2(new_n943), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n970), .B1(new_n920), .B2(new_n921), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n594), .A2(G197gat), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(G1352gat));
  NOR3_X1   g772(.A1(new_n967), .A2(G204gat), .A3(new_n700), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT62), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n971), .A2(new_n699), .ZN(new_n976));
  INV_X1    g775(.A(G204gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(G1353gat));
  AOI211_X1 g777(.A(new_n769), .B(new_n970), .C1(new_n920), .C2(new_n921), .ZN(new_n979));
  OAI21_X1  g778(.A(KEYINPUT63), .B1(new_n979), .B2(new_n259), .ZN(new_n980));
  INV_X1    g779(.A(new_n970), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n922), .A2(new_n677), .A3(new_n981), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT63), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n982), .A2(new_n983), .A3(G211gat), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n968), .A2(new_n259), .A3(new_n677), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT126), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n980), .A2(new_n984), .A3(new_n986), .ZN(G1354gat));
  AOI21_X1  g786(.A(G218gat), .B1(new_n968), .B2(new_n745), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n704), .A2(new_n260), .ZN(new_n989));
  XNOR2_X1  g788(.A(new_n989), .B(KEYINPUT127), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n988), .B1(new_n971), .B2(new_n990), .ZN(G1355gat));
endmodule


