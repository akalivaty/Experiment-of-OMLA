//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 0 0 0 1 1 0 1 1 1 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n796, new_n797, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n998, new_n999;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G228gat), .A2(G233gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n207));
  INV_X1    g006(.A(G211gat), .ZN(new_n208));
  INV_X1    g007(.A(G218gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT76), .ZN(new_n211));
  NOR2_X1   g010(.A1(G211gat), .A2(G218gat), .ZN(new_n212));
  OR3_X1    g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n211), .B1(new_n210), .B2(new_n212), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT88), .ZN(new_n216));
  OR2_X1    g015(.A1(G197gat), .A2(G204gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(G197gat), .A2(G204gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(KEYINPUT22), .B2(new_n210), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT88), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n213), .A2(new_n222), .A3(new_n214), .ZN(new_n223));
  AND3_X1   g022(.A1(new_n216), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT29), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(new_n216), .B2(new_n221), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n207), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G155gat), .A2(G162gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT2), .ZN(new_n229));
  INV_X1    g028(.A(G148gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n230), .A2(G141gat), .ZN(new_n231));
  INV_X1    g030(.A(G141gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n232), .A2(G148gat), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n229), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  OR2_X1    g033(.A1(G155gat), .A2(G162gat), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n235), .A2(KEYINPUT78), .A3(new_n228), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT78), .B1(new_n235), .B2(new_n228), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n234), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT79), .B1(new_n232), .B2(G148gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT79), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(new_n230), .A3(G141gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n232), .A2(G148gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n239), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT80), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n235), .A2(new_n244), .A3(new_n228), .ZN(new_n245));
  AND2_X1   g044(.A1(G155gat), .A2(G162gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(G155gat), .A2(G162gat), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT80), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n243), .A2(new_n229), .A3(new_n245), .A4(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n238), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n206), .B1(new_n227), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n213), .A2(KEYINPUT75), .A3(new_n214), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(new_n220), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n238), .A2(new_n249), .A3(new_n207), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(new_n225), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  OR2_X1    g055(.A1(new_n256), .A2(KEYINPUT89), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(KEYINPUT89), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n251), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n238), .A2(new_n249), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n252), .B(new_n221), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(new_n225), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n260), .B1(new_n262), .B2(new_n207), .ZN(new_n263));
  INV_X1    g062(.A(new_n256), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n206), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT31), .B(G50gat), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n259), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n267), .B1(new_n259), .B2(new_n265), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n204), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n259), .A2(new_n265), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(new_n266), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n259), .A2(new_n265), .A3(new_n267), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n272), .A2(new_n203), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  OR2_X1    g074(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n276));
  INV_X1    g075(.A(G183gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G183gat), .A2(G190gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT65), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT24), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT24), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n280), .A2(KEYINPUT65), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n279), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT64), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(KEYINPUT23), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT25), .ZN(new_n291));
  INV_X1    g090(.A(new_n286), .ZN(new_n292));
  NAND2_X1  g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT23), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n291), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n285), .A2(new_n290), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n283), .A2(new_n277), .ZN(new_n297));
  NAND2_X1  g096(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(G190gat), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G190gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n300), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n286), .A2(KEYINPUT23), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT23), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n304), .B1(G169gat), .B2(G176gat), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n303), .B1(new_n305), .B2(new_n286), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n291), .B1(new_n302), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n296), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT69), .ZN(new_n309));
  INV_X1    g108(.A(G120gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G113gat), .ZN(new_n311));
  INV_X1    g110(.A(G113gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G120gat), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT1), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G127gat), .B(G134gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n309), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G134gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G127gat), .ZN(new_n318));
  INV_X1    g117(.A(G127gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G134gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(G113gat), .B(G120gat), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n321), .B(KEYINPUT69), .C1(new_n322), .C2(KEYINPUT1), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT70), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n313), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n312), .A2(KEYINPUT70), .A3(G120gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(new_n311), .A3(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n321), .A2(KEYINPUT1), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n316), .A2(new_n323), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT68), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n331), .A2(new_n332), .A3(new_n292), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT26), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n288), .A2(new_n334), .A3(new_n289), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT68), .B1(new_n330), .B2(new_n286), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  XOR2_X1   g136(.A(KEYINPUT27), .B(G183gat), .Z(new_n338));
  NAND2_X1  g137(.A1(new_n276), .A2(new_n278), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT28), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n278), .ZN(new_n341));
  NOR2_X1   g140(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT28), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT27), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n345), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT67), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT27), .B1(new_n347), .B2(new_n277), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n343), .A2(new_n344), .A3(new_n346), .A4(new_n348), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n337), .A2(new_n340), .A3(new_n280), .A4(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n308), .A2(new_n329), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT71), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n308), .A2(new_n350), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n328), .A2(new_n327), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT1), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n312), .A2(G120gat), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n310), .A2(G113gat), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT69), .B1(new_n359), .B2(new_n321), .ZN(new_n360));
  NOR3_X1   g159(.A1(new_n314), .A2(new_n309), .A3(new_n315), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n355), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n354), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G227gat), .A2(G233gat), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n308), .A2(new_n350), .A3(new_n329), .A4(KEYINPUT71), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n353), .A2(new_n363), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n366), .B(KEYINPUT34), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT32), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n353), .A2(new_n365), .A3(new_n363), .ZN(new_n369));
  INV_X1    g168(.A(new_n364), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT33), .B1(new_n369), .B2(new_n370), .ZN(new_n372));
  XNOR2_X1  g171(.A(G15gat), .B(G43gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n373), .B(KEYINPUT72), .ZN(new_n374));
  XNOR2_X1  g173(.A(G71gat), .B(G99gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NOR3_X1   g176(.A1(new_n371), .A2(new_n372), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n369), .A2(new_n370), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT33), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT73), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n380), .B1(new_n376), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n382), .B1(new_n381), .B2(new_n376), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n379), .A2(KEYINPUT32), .A3(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n367), .B1(new_n378), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n371), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n379), .A2(new_n380), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n386), .A2(new_n387), .A3(new_n376), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT34), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n366), .B(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n371), .A2(new_n383), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n388), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n385), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n275), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G226gat), .A2(G233gat), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n396), .B1(new_n354), .B2(new_n225), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n395), .B1(new_n308), .B2(new_n350), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n253), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n398), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT29), .B1(new_n308), .B2(new_n350), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n400), .B(new_n261), .C1(new_n396), .C2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G8gat), .B(G36gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(KEYINPUT77), .ZN(new_n406));
  XNOR2_X1  g205(.A(G64gat), .B(G92gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n404), .A2(KEYINPUT30), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n408), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n403), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT30), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n412), .B1(new_n403), .B2(new_n410), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n409), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n207), .B1(new_n238), .B2(new_n249), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT81), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n362), .B(new_n254), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n417), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n316), .A2(new_n323), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n422), .A2(new_n238), .A3(new_n249), .A4(new_n355), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT4), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT4), .B1(new_n260), .B2(new_n329), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT85), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n424), .B1(new_n362), .B2(new_n250), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT85), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n260), .A2(new_n329), .A3(KEYINPUT4), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n421), .B1(new_n427), .B2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(G225gat), .A2(G233gat), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(G1gat), .B(G29gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n439), .B(KEYINPUT0), .ZN(new_n440));
  XNOR2_X1  g239(.A(G57gat), .B(G85gat), .ZN(new_n441));
  XOR2_X1   g240(.A(new_n440), .B(new_n441), .Z(new_n442));
  NAND2_X1  g241(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n428), .A2(new_n435), .A3(new_n430), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT81), .B1(new_n260), .B2(new_n207), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n445), .A2(new_n419), .A3(new_n362), .A4(new_n254), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n423), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n422), .A2(new_n355), .B1(new_n238), .B2(new_n249), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n436), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT83), .B1(new_n450), .B2(new_n434), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n362), .A2(new_n250), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n435), .B1(new_n452), .B2(new_n423), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT83), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n453), .A2(new_n454), .A3(new_n433), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n447), .B1(new_n451), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT84), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n450), .A2(KEYINPUT83), .A3(new_n434), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n454), .B1(new_n453), .B2(new_n433), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT84), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n461), .A3(new_n447), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n443), .B1(new_n457), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT86), .B1(new_n463), .B2(KEYINPUT6), .ZN(new_n464));
  AOI221_X4 g263(.A(KEYINPUT84), .B1(new_n444), .B2(new_n446), .C1(new_n458), .C2(new_n459), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n461), .B1(new_n460), .B2(new_n447), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n438), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n442), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n468), .B1(new_n432), .B2(new_n437), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n470), .B1(new_n465), .B2(new_n466), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT86), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n464), .A2(new_n469), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n467), .A2(KEYINPUT6), .A3(new_n468), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT87), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n467), .A2(KEYINPUT87), .A3(KEYINPUT6), .A4(new_n468), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n394), .B(new_n415), .C1(new_n475), .C2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n438), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n482), .B1(new_n457), .B2(new_n462), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n473), .B(new_n471), .C1(new_n483), .C2(new_n442), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n478), .A2(new_n479), .A3(new_n484), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n275), .A2(KEYINPUT35), .A3(new_n414), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT74), .B1(new_n385), .B2(new_n392), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT74), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n371), .A2(new_n377), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n384), .B1(new_n387), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n489), .B1(new_n491), .B2(new_n390), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT94), .B1(new_n488), .B2(new_n492), .ZN(new_n493));
  NOR3_X1   g292(.A1(new_n378), .A2(new_n367), .A3(new_n384), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n390), .B1(new_n388), .B2(new_n391), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n489), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n491), .A2(new_n390), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT74), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT94), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n493), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g300(.A1(KEYINPUT35), .A2(new_n481), .B1(new_n487), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT92), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT37), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n340), .A2(new_n280), .A3(new_n349), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n505), .A2(new_n337), .B1(new_n307), .B2(new_n296), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n395), .B1(new_n506), .B2(KEYINPUT29), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n261), .B1(new_n507), .B2(new_n400), .ZN(new_n508));
  NOR3_X1   g307(.A1(new_n397), .A2(new_n398), .A3(new_n253), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n504), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n399), .A2(new_n402), .A3(KEYINPUT37), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n408), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT38), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n503), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n399), .A2(new_n402), .A3(KEYINPUT37), .ZN(new_n515));
  AOI21_X1  g314(.A(KEYINPUT37), .B1(new_n399), .B2(new_n402), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n410), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(KEYINPUT92), .A3(KEYINPUT38), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  OAI22_X1  g318(.A1(new_n517), .A2(KEYINPUT38), .B1(new_n403), .B2(new_n410), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n484), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n480), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT93), .ZN(new_n524));
  INV_X1    g323(.A(new_n275), .ZN(new_n525));
  XOR2_X1   g324(.A(KEYINPUT91), .B(KEYINPUT39), .Z(new_n526));
  INV_X1    g325(.A(KEYINPUT90), .ZN(new_n527));
  NOR3_X1   g326(.A1(new_n432), .A2(new_n527), .A3(new_n435), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n429), .B1(new_n428), .B2(new_n430), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n446), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT90), .B1(new_n531), .B2(new_n436), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n526), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n527), .B1(new_n432), .B2(new_n435), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n531), .A2(KEYINPUT90), .A3(new_n436), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT39), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n448), .A2(new_n449), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n536), .B1(new_n537), .B2(new_n435), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n534), .A2(new_n535), .A3(new_n538), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n533), .A2(KEYINPUT40), .A3(new_n442), .A4(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n540), .A2(new_n469), .A3(new_n414), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n534), .A2(new_n535), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n468), .B1(new_n542), .B2(new_n526), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT40), .B1(new_n543), .B2(new_n539), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n525), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  NOR3_X1   g344(.A1(new_n523), .A2(new_n524), .A3(new_n545), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n540), .A2(new_n469), .A3(new_n414), .ZN(new_n547));
  INV_X1    g346(.A(new_n544), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n275), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n457), .A2(new_n462), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT6), .B1(new_n550), .B2(new_n470), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n520), .B1(new_n551), .B2(new_n469), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n552), .A2(new_n479), .A3(new_n478), .A4(new_n519), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT93), .B1(new_n549), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n546), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT36), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n393), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n496), .A2(new_n498), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n557), .B1(new_n558), .B2(new_n556), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n415), .B1(new_n475), .B2(new_n480), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n559), .B1(new_n560), .B2(new_n275), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n502), .B1(new_n555), .B2(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(G43gat), .B(G50gat), .Z(new_n563));
  INV_X1    g362(.A(KEYINPUT15), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NOR3_X1   g365(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(G29gat), .A2(G36gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n563), .A2(new_n564), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n566), .A2(new_n570), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT96), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n567), .B1(new_n574), .B2(new_n569), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n575), .B1(new_n574), .B2(new_n569), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n571), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT97), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n577), .A2(new_n578), .A3(new_n565), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n578), .B1(new_n577), .B2(new_n565), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n573), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT17), .ZN(new_n582));
  INV_X1    g381(.A(G8gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(G15gat), .B(G22gat), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT16), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n584), .B1(new_n585), .B2(G1gat), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n583), .B1(new_n586), .B2(KEYINPUT98), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n586), .B1(G1gat), .B2(new_n584), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n582), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G229gat), .A2(G233gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n581), .A2(new_n589), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT18), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n581), .B(new_n589), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n592), .B(KEYINPUT13), .Z(new_n597));
  AOI22_X1  g396(.A1(new_n594), .A2(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n591), .A2(KEYINPUT18), .A3(new_n592), .A4(new_n593), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n599), .A2(KEYINPUT99), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(KEYINPUT99), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n598), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n594), .A2(new_n595), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT100), .ZN(new_n604));
  XNOR2_X1  g403(.A(G113gat), .B(G141gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(G169gat), .B(G197gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT95), .B(KEYINPUT11), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n609), .B(KEYINPUT12), .Z(new_n610));
  NAND3_X1  g409(.A1(new_n602), .A2(new_n604), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n604), .A2(new_n610), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n599), .B(KEYINPUT99), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n612), .A2(new_n613), .A3(new_n598), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT101), .B1(new_n562), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n560), .A2(new_n275), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n524), .B1(new_n523), .B2(new_n545), .ZN(new_n619));
  INV_X1    g418(.A(new_n559), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n549), .A2(KEYINPUT93), .A3(new_n553), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n618), .A2(new_n619), .A3(new_n620), .A4(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n481), .A2(KEYINPUT35), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n487), .A2(new_n501), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT101), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n626), .A2(new_n627), .A3(new_n615), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n617), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G232gat), .A2(G233gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT103), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT41), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G134gat), .B(G162gat), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n633), .B(new_n634), .Z(new_n635));
  XOR2_X1   g434(.A(KEYINPUT104), .B(KEYINPUT105), .Z(new_n636));
  XOR2_X1   g435(.A(new_n635), .B(new_n636), .Z(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G85gat), .A2(G92gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT7), .ZN(new_n640));
  NAND2_X1  g439(.A1(G99gat), .A2(G106gat), .ZN(new_n641));
  INV_X1    g440(.A(G85gat), .ZN(new_n642));
  INV_X1    g441(.A(G92gat), .ZN(new_n643));
  AOI22_X1  g442(.A1(KEYINPUT8), .A2(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G99gat), .B(G106gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n581), .A2(KEYINPUT17), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n581), .A2(KEYINPUT17), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(KEYINPUT106), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT106), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n582), .A2(new_n653), .A3(new_n648), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G190gat), .B(G218gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n656), .B(KEYINPUT107), .Z(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n631), .A2(new_n632), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n659), .B1(new_n581), .B2(new_n647), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n655), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n658), .B1(new_n655), .B2(new_n660), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n638), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n663), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n665), .A2(new_n637), .A3(new_n661), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  XOR2_X1   g467(.A(G57gat), .B(G64gat), .Z(new_n669));
  INV_X1    g468(.A(KEYINPUT9), .ZN(new_n670));
  INV_X1    g469(.A(G71gat), .ZN(new_n671));
  INV_X1    g470(.A(G78gat), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g473(.A(G71gat), .B(G78gat), .Z(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT21), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(G231gat), .A2(G233gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(G127gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n676), .B(KEYINPUT102), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n589), .B1(new_n682), .B2(KEYINPUT21), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n681), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(G155gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(G183gat), .B(G211gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n684), .A2(new_n688), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n668), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(G230gat), .ZN(new_n693));
  INV_X1    g492(.A(G233gat), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n647), .B(new_n676), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT10), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n682), .A2(KEYINPUT10), .A3(new_n647), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n696), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(new_n696), .B2(new_n697), .ZN(new_n702));
  XNOR2_X1  g501(.A(G120gat), .B(G148gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(G176gat), .B(G204gat), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n703), .B(new_n704), .Z(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n702), .A2(new_n706), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n692), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n629), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n475), .A2(new_n480), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g513(.A(new_n714), .B(G1gat), .Z(G1324gat));
  AOI21_X1  g514(.A(new_n627), .B1(new_n626), .B2(new_n615), .ZN(new_n716));
  AOI211_X1 g515(.A(KEYINPUT101), .B(new_n616), .C1(new_n622), .C2(new_n625), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n414), .B(new_n710), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n629), .A2(KEYINPUT108), .A3(new_n414), .A4(new_n710), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT16), .B(G8gat), .Z(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT42), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n720), .A2(new_n721), .A3(G8gat), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n723), .A2(KEYINPUT42), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n718), .A2(new_n728), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n726), .A2(new_n730), .A3(KEYINPUT109), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT109), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT42), .B1(new_n722), .B2(new_n723), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n727), .A2(new_n729), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n731), .A2(new_n735), .ZN(G1325gat));
  OAI21_X1  g535(.A(G15gat), .B1(new_n711), .B2(new_n620), .ZN(new_n737));
  INV_X1    g536(.A(new_n501), .ZN(new_n738));
  OR2_X1    g537(.A1(new_n738), .A2(G15gat), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n737), .B1(new_n711), .B2(new_n739), .ZN(G1326gat));
  NOR2_X1   g539(.A1(new_n711), .A2(new_n525), .ZN(new_n741));
  XOR2_X1   g540(.A(KEYINPUT43), .B(G22gat), .Z(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1327gat));
  NOR2_X1   g542(.A1(new_n691), .A2(new_n709), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  AOI211_X1 g544(.A(new_n668), .B(new_n745), .C1(new_n617), .C2(new_n628), .ZN(new_n746));
  INV_X1    g545(.A(G29gat), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n746), .A2(new_n747), .A3(new_n712), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT45), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n562), .A2(new_n668), .ZN(new_n751));
  XOR2_X1   g550(.A(KEYINPUT110), .B(KEYINPUT44), .Z(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n626), .A2(new_n667), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n754), .B1(new_n755), .B2(KEYINPUT44), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n616), .A2(new_n745), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(G29gat), .B1(new_n759), .B2(new_n713), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n748), .A2(new_n749), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n750), .A2(new_n760), .A3(new_n761), .ZN(G1328gat));
  INV_X1    g561(.A(G36gat), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n746), .A2(new_n763), .A3(new_n414), .ZN(new_n764));
  XNOR2_X1  g563(.A(KEYINPUT111), .B(KEYINPUT46), .ZN(new_n765));
  OR2_X1    g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(G36gat), .B1(new_n759), .B2(new_n415), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n764), .A2(new_n765), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(G1329gat));
  AND4_X1   g568(.A1(G43gat), .A2(new_n757), .A3(new_n559), .A4(new_n758), .ZN(new_n770));
  AOI21_X1  g569(.A(G43gat), .B1(new_n746), .B2(new_n501), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT47), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(G1330gat));
  OAI21_X1  g573(.A(G50gat), .B1(new_n759), .B2(new_n525), .ZN(new_n775));
  INV_X1    g574(.A(G50gat), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n746), .A2(new_n776), .A3(new_n275), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT48), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(G1331gat));
  INV_X1    g579(.A(new_n709), .ZN(new_n781));
  NOR4_X1   g580(.A1(new_n562), .A2(new_n615), .A3(new_n692), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n712), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(G57gat), .ZN(G1332gat));
  INV_X1    g583(.A(KEYINPUT49), .ZN(new_n785));
  INV_X1    g584(.A(G64gat), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n414), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  XOR2_X1   g586(.A(new_n787), .B(KEYINPUT112), .Z(new_n788));
  NAND2_X1  g587(.A1(new_n782), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n785), .A2(new_n786), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n789), .B(new_n790), .ZN(G1333gat));
  AOI21_X1  g590(.A(new_n671), .B1(new_n782), .B2(new_n559), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n738), .A2(G71gat), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n792), .B1(new_n782), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g594(.A1(new_n782), .A2(new_n275), .ZN(new_n796));
  XNOR2_X1  g595(.A(KEYINPUT113), .B(G78gat), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n796), .B(new_n797), .ZN(G1335gat));
  NOR2_X1   g597(.A1(new_n615), .A2(new_n691), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n751), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n781), .B1(new_n800), .B2(KEYINPUT51), .ZN(new_n801));
  INV_X1    g600(.A(new_n799), .ZN(new_n802));
  OR3_X1    g601(.A1(new_n754), .A2(KEYINPUT51), .A3(new_n802), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n804), .A2(new_n642), .A3(new_n712), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n802), .A2(new_n781), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n757), .A2(new_n806), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n807), .A2(new_n712), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n805), .B1(new_n808), .B2(new_n642), .ZN(G1336gat));
  NAND2_X1  g608(.A1(new_n800), .A2(KEYINPUT51), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n415), .A2(G92gat), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n810), .A2(new_n803), .A3(new_n709), .A4(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n757), .A2(new_n414), .A3(new_n806), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(G92gat), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n812), .A2(new_n813), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT52), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n812), .A2(KEYINPUT115), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n812), .A2(KEYINPUT115), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n820), .A2(new_n821), .A3(new_n816), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n819), .A2(new_n823), .ZN(G1337gat));
  AOI21_X1  g623(.A(G99gat), .B1(new_n804), .B2(new_n501), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n559), .A2(G99gat), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n825), .B1(new_n807), .B2(new_n826), .ZN(G1338gat));
  INV_X1    g626(.A(G106gat), .ZN(new_n828));
  AND4_X1   g627(.A1(new_n828), .A2(new_n801), .A3(new_n275), .A4(new_n803), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n807), .A2(new_n275), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n830), .B(new_n831), .C1(new_n832), .C2(new_n828), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n828), .B1(new_n807), .B2(new_n275), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT53), .B1(new_n834), .B2(new_n829), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(G1339gat));
  NOR3_X1   g635(.A1(new_n692), .A2(new_n615), .A3(new_n709), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT55), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n699), .A2(new_n700), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n695), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n840), .A2(KEYINPUT54), .A3(new_n701), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n706), .B1(new_n701), .B2(KEYINPUT54), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n838), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n842), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n840), .A2(KEYINPUT54), .A3(new_n701), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(KEYINPUT55), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n843), .A2(new_n707), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n847), .B1(new_n611), .B2(new_n614), .ZN(new_n848));
  INV_X1    g647(.A(new_n610), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n849), .B(new_n598), .C1(new_n600), .C2(new_n601), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n592), .B1(new_n591), .B2(new_n593), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n596), .A2(new_n597), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n609), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(new_n781), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n668), .B1(new_n848), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n847), .B1(new_n664), .B2(new_n666), .ZN(new_n857));
  INV_X1    g656(.A(new_n854), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n691), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n837), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n713), .A2(new_n414), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n738), .A2(new_n275), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n866), .A2(new_n312), .A3(new_n616), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n863), .A2(new_n712), .A3(new_n394), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n868), .A2(new_n414), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n615), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n867), .B1(new_n870), .B2(new_n312), .ZN(G1340gat));
  NOR3_X1   g670(.A1(new_n866), .A2(new_n310), .A3(new_n781), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n869), .A2(new_n709), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n872), .B1(new_n873), .B2(new_n310), .ZN(G1341gat));
  NAND3_X1  g673(.A1(new_n869), .A2(new_n319), .A3(new_n691), .ZN(new_n875));
  OAI21_X1  g674(.A(G127gat), .B1(new_n866), .B2(new_n861), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(G1342gat));
  NAND3_X1  g676(.A1(new_n667), .A2(new_n317), .A3(new_n415), .ZN(new_n878));
  OR3_X1    g677(.A1(new_n868), .A2(KEYINPUT56), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(G134gat), .B1(new_n866), .B2(new_n668), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT56), .B1(new_n868), .B2(new_n878), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT116), .ZN(G1343gat));
  OR3_X1    g682(.A1(new_n862), .A2(KEYINPUT118), .A3(new_n713), .ZN(new_n884));
  OAI21_X1  g683(.A(KEYINPUT118), .B1(new_n862), .B2(new_n713), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n559), .A2(new_n525), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n887), .A2(new_n414), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n232), .A3(new_n615), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT58), .ZN(new_n890));
  OR2_X1    g689(.A1(new_n890), .A2(KEYINPUT119), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n892), .B1(new_n862), .B2(new_n525), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n691), .B1(new_n856), .B2(new_n859), .ZN(new_n894));
  OAI211_X1 g693(.A(KEYINPUT57), .B(new_n275), .C1(new_n894), .C2(new_n837), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n864), .A2(new_n620), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(new_n616), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n890), .A2(G141gat), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n889), .B(new_n891), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n615), .A2(new_n232), .ZN(new_n903));
  NOR4_X1   g702(.A1(new_n887), .A2(KEYINPUT119), .A3(new_n414), .A4(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT117), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n899), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n896), .A2(KEYINPUT117), .A3(new_n898), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(new_n615), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n904), .B1(new_n908), .B2(G141gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n902), .B1(new_n909), .B2(new_n890), .ZN(G1344gat));
  NAND3_X1  g709(.A1(new_n888), .A2(new_n230), .A3(new_n709), .ZN(new_n911));
  XOR2_X1   g710(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n912));
  AOI21_X1  g711(.A(new_n781), .B1(new_n897), .B2(KEYINPUT121), .ZN(new_n913));
  INV_X1    g712(.A(new_n837), .ZN(new_n914));
  INV_X1    g713(.A(new_n847), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n615), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n858), .A2(new_n709), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n854), .B1(new_n857), .B2(KEYINPUT122), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n667), .A2(new_n915), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT122), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI22_X1  g721(.A1(new_n918), .A2(new_n668), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n914), .B1(new_n923), .B2(new_n691), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT57), .B1(new_n924), .B2(new_n275), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT123), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n895), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n919), .A2(new_n922), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n856), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n837), .B1(new_n929), .B2(new_n861), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n892), .B1(new_n930), .B2(new_n525), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n931), .A2(KEYINPUT123), .ZN(new_n932));
  OAI221_X1 g731(.A(new_n913), .B1(KEYINPUT121), .B2(new_n897), .C1(new_n927), .C2(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n912), .B1(new_n933), .B2(G148gat), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n230), .A2(KEYINPUT59), .ZN(new_n935));
  AOI21_X1  g734(.A(KEYINPUT117), .B1(new_n896), .B2(new_n898), .ZN(new_n936));
  AOI211_X1 g735(.A(new_n905), .B(new_n897), .C1(new_n893), .C2(new_n895), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n935), .B1(new_n938), .B2(new_n709), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n911), .B1(new_n934), .B2(new_n939), .ZN(G1345gat));
  INV_X1    g739(.A(G155gat), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n888), .A2(new_n941), .A3(new_n691), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n936), .A2(new_n937), .A3(new_n861), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n942), .B1(new_n943), .B2(new_n941), .ZN(G1346gat));
  OR4_X1    g743(.A1(G162gat), .A2(new_n887), .A3(new_n414), .A4(new_n668), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n936), .A2(new_n937), .A3(new_n668), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n947));
  OAI21_X1  g746(.A(G162gat), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NOR4_X1   g747(.A1(new_n936), .A2(new_n937), .A3(KEYINPUT124), .A4(new_n668), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(G1347gat));
  NAND4_X1  g749(.A1(new_n863), .A2(new_n713), .A3(new_n414), .A4(new_n865), .ZN(new_n951));
  INV_X1    g750(.A(G169gat), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n951), .A2(new_n952), .A3(new_n616), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n862), .A2(new_n712), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n275), .A2(new_n393), .A3(new_n415), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(new_n615), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n953), .B1(new_n958), .B2(new_n952), .ZN(G1348gat));
  INV_X1    g758(.A(new_n951), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n960), .A2(G176gat), .A3(new_n709), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT125), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n961), .A2(new_n962), .ZN(new_n964));
  AOI21_X1  g763(.A(G176gat), .B1(new_n957), .B2(new_n709), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(G1349gat));
  OR3_X1    g765(.A1(new_n956), .A2(new_n338), .A3(new_n861), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n968), .B1(new_n951), .B2(new_n861), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(G183gat), .ZN(new_n970));
  NOR3_X1   g769(.A1(new_n951), .A2(new_n968), .A3(new_n861), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n967), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g772(.A(G190gat), .B1(new_n951), .B2(new_n668), .ZN(new_n974));
  OR2_X1    g773(.A1(new_n974), .A2(KEYINPUT127), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(KEYINPUT127), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n975), .A2(KEYINPUT61), .A3(new_n976), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n957), .A2(new_n343), .A3(new_n667), .ZN(new_n978));
  OAI211_X1 g777(.A(new_n977), .B(new_n978), .C1(KEYINPUT61), .C2(new_n976), .ZN(G1351gat));
  NOR3_X1   g778(.A1(new_n712), .A2(new_n559), .A3(new_n415), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n980), .B1(new_n927), .B2(new_n932), .ZN(new_n981));
  INV_X1    g780(.A(G197gat), .ZN(new_n982));
  NOR3_X1   g781(.A1(new_n981), .A2(new_n982), .A3(new_n616), .ZN(new_n983));
  NOR3_X1   g782(.A1(new_n559), .A2(new_n415), .A3(new_n525), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n954), .A2(new_n984), .ZN(new_n985));
  INV_X1    g784(.A(new_n985), .ZN(new_n986));
  AOI21_X1  g785(.A(G197gat), .B1(new_n986), .B2(new_n615), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n983), .A2(new_n987), .ZN(G1352gat));
  OAI21_X1  g787(.A(G204gat), .B1(new_n981), .B2(new_n781), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n985), .A2(G204gat), .A3(new_n781), .ZN(new_n990));
  XNOR2_X1  g789(.A(new_n990), .B(KEYINPUT62), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n989), .A2(new_n991), .ZN(G1353gat));
  NAND3_X1  g791(.A1(new_n986), .A2(new_n208), .A3(new_n691), .ZN(new_n993));
  OAI211_X1 g792(.A(new_n691), .B(new_n980), .C1(new_n927), .C2(new_n932), .ZN(new_n994));
  AND3_X1   g793(.A1(new_n994), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n995));
  AOI21_X1  g794(.A(KEYINPUT63), .B1(new_n994), .B2(G211gat), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n993), .B1(new_n995), .B2(new_n996), .ZN(G1354gat));
  OAI21_X1  g796(.A(G218gat), .B1(new_n981), .B2(new_n668), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n986), .A2(new_n209), .A3(new_n667), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(new_n999), .ZN(G1355gat));
endmodule


