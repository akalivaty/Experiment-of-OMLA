//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 0 1 0 1 0 0 0 0 0 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n626, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XNOR2_X1  g016(.A(KEYINPUT65), .B(G108), .ZN(G238));
  AND2_X1   g017(.A1(G2072), .A2(G2078), .ZN(new_n443));
  NAND3_X1  g018(.A1(new_n443), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n448));
  AND2_X1   g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  NAND2_X1  g025(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n449), .A2(G2106), .ZN(G217));
  OR4_X1    g027(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n453), .B(new_n454), .Z(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT68), .Z(G325));
  XOR2_X1   g034(.A(G325), .B(KEYINPUT69), .Z(G261));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT70), .Z(new_n463));
  AOI21_X1  g038(.A(new_n463), .B1(new_n455), .B2(G2106), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G125), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n465), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  OAI211_X1 g046(.A(G137), .B(new_n465), .C1(new_n466), .C2(new_n467), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n465), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G112), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n466), .A2(new_n467), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT71), .Z(new_n485));
  NOR2_X1   g060(.A1(new_n482), .A2(new_n465), .ZN(new_n486));
  AOI211_X1 g061(.A(new_n481), .B(new_n485), .C1(G124), .C2(new_n486), .ZN(G162));
  OAI211_X1 g062(.A(G126), .B(G2105), .C1(new_n466), .C2(new_n467), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n493), .A2(new_n465), .A3(G138), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT72), .B1(new_n482), .B2(new_n494), .ZN(new_n495));
  OR2_X1    g070(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n496));
  NAND2_X1  g071(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT72), .ZN(new_n499));
  AND3_X1   g074(.A1(new_n493), .A2(new_n465), .A3(G138), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g077(.A(G138), .B(new_n465), .C1(new_n466), .C2(new_n467), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n492), .B1(new_n502), .B2(new_n504), .ZN(G164));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT6), .B(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  AND2_X1   g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  AND2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n515), .A2(new_n516), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n513), .A2(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  INV_X1    g100(.A(new_n521), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT76), .B(G89), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n526), .A2(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g106(.A(KEYINPUT73), .B1(new_n518), .B2(new_n517), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT73), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n508), .A2(new_n533), .A3(new_n509), .ZN(new_n534));
  AND2_X1   g109(.A1(G63), .A2(G651), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT75), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT74), .B(G51), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n514), .A2(new_n538), .A3(G543), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n537), .B1(new_n536), .B2(new_n539), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n531), .B1(new_n540), .B2(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  AND2_X1   g118(.A1(new_n532), .A2(new_n534), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n544), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n512), .ZN(new_n546));
  INV_X1    g121(.A(G52), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n515), .A2(new_n547), .B1(new_n521), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(G171));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n532), .A2(new_n534), .ZN(new_n552));
  INV_X1    g127(.A(G56), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G651), .ZN(new_n555));
  INV_X1    g130(.A(new_n515), .ZN(new_n556));
  AOI22_X1  g131(.A1(G43), .A2(new_n556), .B1(new_n526), .B2(G81), .ZN(new_n557));
  AND2_X1   g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT77), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  NAND3_X1  g140(.A1(new_n526), .A2(KEYINPUT78), .A3(G91), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT78), .ZN(new_n567));
  INV_X1    g142(.A(G91), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n521), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(new_n510), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n566), .A2(new_n569), .B1(new_n573), .B2(G651), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n514), .A2(G53), .A3(G543), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT9), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(G299));
  INV_X1    g152(.A(G171), .ZN(G301));
  OAI21_X1  g153(.A(G651), .B1(new_n544), .B2(G74), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n514), .A2(G49), .A3(G543), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n514), .A2(KEYINPUT79), .A3(G49), .A4(G543), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n526), .A2(G87), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n579), .A2(new_n584), .A3(new_n585), .ZN(G288));
  NAND3_X1  g161(.A1(new_n510), .A2(new_n514), .A3(G86), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n514), .A2(G48), .A3(G543), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(G61), .B1(new_n518), .B2(new_n517), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n512), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G305));
  NAND2_X1  g169(.A1(new_n544), .A2(G60), .ZN(new_n595));
  NAND2_X1  g170(.A1(G72), .A2(G543), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n512), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(G47), .ZN(new_n598));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  OAI22_X1  g174(.A1(new_n515), .A2(new_n598), .B1(new_n521), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n526), .A2(G92), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT81), .ZN(new_n605));
  XOR2_X1   g180(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n604), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(new_n606), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n510), .A2(G66), .ZN(new_n612));
  INV_X1    g187(.A(G79), .ZN(new_n613));
  OAI21_X1  g188(.A(KEYINPUT82), .B1(new_n613), .B2(new_n507), .ZN(new_n614));
  OR3_X1    g189(.A1(new_n613), .A2(new_n507), .A3(KEYINPUT82), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n612), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n616), .A2(G651), .B1(new_n556), .B2(G54), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n608), .A2(new_n611), .A3(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n603), .B1(new_n619), .B2(G868), .ZN(G284));
  OAI21_X1  g195(.A(new_n603), .B1(new_n619), .B2(G868), .ZN(G321));
  NAND2_X1  g196(.A1(G286), .A2(G868), .ZN(new_n622));
  INV_X1    g197(.A(G299), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G868), .ZN(G297));
  OAI21_X1  g199(.A(new_n622), .B1(new_n623), .B2(G868), .ZN(G280));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n619), .B1(new_n626), .B2(G860), .ZN(G148));
  NAND2_X1  g202(.A1(new_n619), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G868), .B2(new_n560), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n498), .A2(new_n473), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n635), .A2(G2100), .ZN(new_n636));
  OAI21_X1  g211(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n637));
  INV_X1    g212(.A(G111), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(G2105), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n486), .A2(G123), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT83), .Z(new_n641));
  AOI211_X1 g216(.A(new_n639), .B(new_n641), .C1(G135), .C2(new_n483), .ZN(new_n642));
  INV_X1    g217(.A(G2096), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n636), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n635), .A2(G2100), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n644), .B(new_n645), .C1(new_n643), .C2(new_n642), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT84), .ZN(G156));
  XNOR2_X1  g222(.A(G2427), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2430), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(KEYINPUT14), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2451), .B(G2454), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT85), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n655), .A2(new_n658), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT86), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT87), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n660), .B1(new_n659), .B2(new_n661), .ZN(new_n665));
  INV_X1    g240(.A(G14), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AND3_X1   g242(.A1(new_n663), .A2(new_n664), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n664), .B1(new_n663), .B2(new_n667), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(G401));
  XOR2_X1   g245(.A(G2067), .B(G2678), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT88), .ZN(new_n672));
  NOR2_X1   g247(.A1(G2072), .A2(G2078), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n443), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2084), .B(G2090), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n672), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n672), .A2(new_n674), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n674), .B(KEYINPUT17), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n679), .B(new_n675), .C1(new_n672), .C2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n675), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n672), .A2(new_n682), .A3(new_n680), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n678), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2096), .B(G2100), .Z(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n684), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT90), .B(KEYINPUT91), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(G227));
  XOR2_X1   g266(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n692));
  XNOR2_X1  g267(.A(G1971), .B(G1976), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1956), .B(G2474), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1961), .B(G1966), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT20), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n695), .B(new_n696), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n699), .B(new_n700), .C1(new_n694), .C2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(G1991), .B(G1996), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1981), .B(G1986), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n705), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n704), .B(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n707), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n708), .A2(new_n712), .ZN(G229));
  NOR2_X1   g288(.A1(G16), .A2(G23), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT95), .Z(new_n715));
  INV_X1    g290(.A(G288), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(G16), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT33), .B(G1976), .Z(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G16), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G22), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G166), .B2(new_n720), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT96), .Z(new_n723));
  AOI21_X1  g298(.A(new_n719), .B1(new_n723), .B2(G1971), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n720), .A2(G6), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(new_n593), .B2(new_n720), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT32), .B(G1981), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT94), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n726), .B(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n717), .B2(new_n718), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n724), .B(new_n730), .C1(G1971), .C2(new_n723), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(KEYINPUT34), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(KEYINPUT34), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n601), .A2(new_n720), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n720), .B2(G24), .ZN(new_n735));
  INV_X1    g310(.A(G1986), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G29), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G25), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT93), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n483), .A2(G131), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n486), .A2(G119), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n465), .A2(G107), .ZN(new_n743));
  OAI21_X1  g318(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n741), .B(new_n742), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n740), .B1(new_n745), .B2(G29), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT35), .B(G1991), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n735), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(G1986), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n732), .A2(new_n733), .A3(new_n737), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(KEYINPUT97), .A2(KEYINPUT36), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT98), .B(KEYINPUT28), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n738), .A2(G26), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n483), .A2(G140), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n486), .A2(G128), .ZN(new_n758));
  OR2_X1    g333(.A1(G104), .A2(G2105), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n759), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n756), .B1(new_n762), .B2(new_n738), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G2067), .ZN(new_n764));
  INV_X1    g339(.A(G11), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(KEYINPUT31), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(KEYINPUT31), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT30), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n768), .A2(G28), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n738), .B1(new_n768), .B2(G28), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n766), .B(new_n767), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n642), .B2(G29), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT24), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n773), .A2(G34), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(G34), .ZN(new_n776));
  AOI21_X1  g351(.A(G29), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n477), .B2(G29), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(G2084), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(G2084), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n772), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n738), .A2(G35), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G162), .B2(new_n738), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT29), .Z(new_n785));
  INV_X1    g360(.A(G2090), .ZN(new_n786));
  AOI211_X1 g361(.A(new_n764), .B(new_n782), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n738), .A2(G27), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G164), .B2(new_n738), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(G2078), .Z(new_n790));
  INV_X1    g365(.A(KEYINPUT103), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n720), .A2(G21), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G168), .B2(new_n720), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT101), .B(G1966), .Z(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n790), .A2(new_n791), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n787), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(G4), .A2(G16), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n619), .B2(G16), .ZN(new_n799));
  INV_X1    g374(.A(G1348), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n560), .A2(new_n720), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n720), .B2(G19), .ZN(new_n803));
  INV_X1    g378(.A(G1341), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT25), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n498), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n809));
  AND3_X1   g384(.A1(new_n483), .A2(KEYINPUT99), .A3(G139), .ZN(new_n810));
  AOI21_X1  g385(.A(KEYINPUT99), .B1(new_n483), .B2(G139), .ZN(new_n811));
  OAI221_X1 g386(.A(new_n808), .B1(new_n465), .B2(new_n809), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  MUX2_X1   g387(.A(G33), .B(new_n812), .S(G29), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G2072), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT104), .B(KEYINPUT23), .Z(new_n815));
  NAND2_X1  g390(.A1(new_n720), .A2(G20), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n623), .B2(new_n720), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(G1956), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n818), .A2(G1956), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n814), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n720), .A2(G5), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G171), .B2(new_n720), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT102), .ZN(new_n824));
  INV_X1    g399(.A(G1961), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n801), .A2(new_n805), .A3(new_n821), .A4(new_n826), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n793), .A2(new_n795), .ZN(new_n828));
  OAI221_X1 g403(.A(new_n828), .B1(new_n791), .B2(new_n790), .C1(new_n785), .C2(new_n786), .ZN(new_n829));
  NOR3_X1   g404(.A1(new_n797), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  OR2_X1    g405(.A1(KEYINPUT97), .A2(KEYINPUT36), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n751), .A2(new_n752), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n738), .A2(G32), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n486), .A2(G129), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT100), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n473), .A2(G105), .ZN(new_n836));
  NAND3_X1  g411(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT26), .ZN(new_n838));
  AOI211_X1 g413(.A(new_n836), .B(new_n838), .C1(G141), .C2(new_n483), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n833), .B1(new_n841), .B2(new_n738), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT27), .ZN(new_n843));
  INV_X1    g418(.A(G1996), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n803), .A2(new_n804), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n824), .A2(new_n825), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n753), .A2(new_n830), .A3(new_n832), .A4(new_n848), .ZN(G150));
  INV_X1    g424(.A(G150), .ZN(G311));
  INV_X1    g425(.A(G55), .ZN(new_n851));
  INV_X1    g426(.A(G93), .ZN(new_n852));
  OAI22_X1  g427(.A1(new_n515), .A2(new_n851), .B1(new_n521), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(G80), .A2(G543), .ZN(new_n854));
  INV_X1    g429(.A(G67), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n552), .B2(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n856), .A2(KEYINPUT105), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n512), .B1(new_n856), .B2(KEYINPUT105), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n853), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(new_n558), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(new_n560), .B2(new_n859), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT38), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n618), .A2(new_n626), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n864), .A2(KEYINPUT39), .ZN(new_n865));
  INV_X1    g440(.A(G860), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(KEYINPUT39), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n859), .A2(new_n866), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT37), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT106), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n868), .A2(KEYINPUT106), .A3(new_n870), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(G145));
  XNOR2_X1  g450(.A(new_n840), .B(new_n812), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n486), .A2(G130), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n465), .A2(G118), .ZN(new_n878));
  OAI21_X1  g453(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n880), .B1(G142), .B2(new_n483), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n633), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n876), .B(new_n882), .ZN(new_n883));
  AOI22_X1  g458(.A1(new_n495), .A2(new_n501), .B1(KEYINPUT4), .B2(new_n503), .ZN(new_n884));
  NAND2_X1  g459(.A1(G126), .A2(G2105), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(new_n496), .B2(new_n497), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n465), .A2(G114), .ZN(new_n887));
  OAI21_X1  g462(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT107), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT107), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n488), .A2(new_n491), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n884), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n761), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n745), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n883), .B(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n642), .B(new_n477), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(G162), .ZN(new_n899));
  AOI21_X1  g474(.A(G37), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(new_n899), .B2(new_n897), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g477(.A1(new_n619), .A2(new_n623), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n618), .A2(G299), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n903), .A2(KEYINPUT41), .A3(new_n904), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI211_X1 g484(.A(new_n628), .B(new_n860), .C1(new_n560), .C2(new_n859), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n861), .A2(new_n626), .A3(new_n619), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n910), .A2(new_n911), .A3(new_n905), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT42), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT42), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n913), .A2(new_n917), .A3(new_n914), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n601), .B(G303), .ZN(new_n920));
  XNOR2_X1  g495(.A(G288), .B(new_n593), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n920), .B(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n919), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n916), .A2(new_n922), .A3(new_n918), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(G868), .A3(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n859), .A2(G868), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n927), .A2(KEYINPUT108), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n924), .A2(KEYINPUT108), .A3(new_n925), .A4(G868), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(G295));
  AND2_X1   g506(.A1(new_n929), .A2(new_n930), .ZN(G331));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n933));
  INV_X1    g508(.A(G37), .ZN(new_n934));
  XNOR2_X1  g509(.A(G171), .B(G168), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n861), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n936), .A2(new_n905), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n861), .A2(new_n935), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(KEYINPUT109), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n861), .A2(new_n941), .A3(new_n935), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n936), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n939), .B1(new_n943), .B2(new_n909), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n934), .B1(new_n944), .B2(new_n923), .ZN(new_n945));
  INV_X1    g520(.A(new_n936), .ZN(new_n946));
  INV_X1    g521(.A(new_n942), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n941), .B1(new_n861), .B2(new_n935), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n909), .ZN(new_n950));
  AOI22_X1  g525(.A1(new_n949), .A2(new_n950), .B1(new_n938), .B2(new_n937), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n951), .A2(new_n922), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n933), .B1(new_n945), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(G37), .B1(new_n951), .B2(new_n922), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n946), .A2(new_n938), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n940), .A2(new_n942), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n950), .A2(new_n955), .B1(new_n956), .B2(new_n937), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT110), .B1(new_n957), .B2(new_n922), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n956), .A2(new_n937), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n909), .B1(new_n946), .B2(new_n938), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n959), .B(new_n923), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n954), .A2(new_n958), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n953), .B1(new_n963), .B2(new_n933), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT44), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n954), .A2(new_n958), .A3(new_n962), .A4(new_n933), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT43), .B1(new_n945), .B2(new_n952), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n965), .A2(new_n970), .ZN(G397));
  XNOR2_X1  g546(.A(new_n840), .B(new_n844), .ZN(new_n972));
  INV_X1    g547(.A(G2067), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n761), .B(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n747), .ZN(new_n976));
  OR2_X1    g551(.A1(new_n745), .A2(new_n976), .ZN(new_n977));
  OAI22_X1  g552(.A1(new_n975), .A2(new_n977), .B1(G2067), .B2(new_n761), .ZN(new_n978));
  INV_X1    g553(.A(G1384), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(new_n884), .B2(new_n893), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(KEYINPUT111), .B(G40), .Z(new_n983));
  NOR3_X1   g558(.A1(new_n470), .A2(new_n475), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n978), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n974), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n986), .B1(new_n988), .B2(new_n840), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n986), .A2(new_n844), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n990), .A2(KEYINPUT46), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n990), .A2(KEYINPUT46), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  XOR2_X1   g568(.A(new_n993), .B(KEYINPUT47), .Z(new_n994));
  NAND3_X1  g569(.A1(new_n986), .A2(new_n736), .A3(new_n601), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT48), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n995), .A2(new_n996), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n745), .A2(new_n976), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n972), .A2(new_n974), .A3(new_n977), .A4(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n998), .B1(new_n1000), .B2(new_n986), .ZN(new_n1001));
  AOI211_X1 g576(.A(new_n987), .B(new_n994), .C1(new_n997), .C2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n1003));
  OAI211_X1 g578(.A(G303), .B(G8), .C1(new_n1003), .C2(KEYINPUT55), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(KEYINPUT55), .ZN(new_n1005));
  XOR2_X1   g580(.A(new_n1005), .B(KEYINPUT115), .Z(new_n1006));
  XNOR2_X1  g581(.A(new_n1004), .B(new_n1006), .ZN(new_n1007));
  XOR2_X1   g582(.A(KEYINPUT113), .B(G2090), .Z(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT50), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1011), .B(new_n979), .C1(new_n884), .C2(new_n893), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1010), .A2(KEYINPUT112), .A3(new_n1012), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n890), .A2(new_n892), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n502), .A2(new_n504), .ZN(new_n1015));
  AOI21_X1  g590(.A(G1384), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(new_n1017), .A3(new_n1011), .ZN(new_n1018));
  AOI211_X1 g593(.A(new_n985), .B(new_n1009), .C1(new_n1013), .C2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n981), .B1(G164), .B2(G1384), .ZN(new_n1020));
  OAI211_X1 g595(.A(KEYINPUT45), .B(new_n979), .C1(new_n884), .C2(new_n893), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1020), .A2(new_n984), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G1971), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  OAI211_X1 g600(.A(G8), .B(new_n1007), .C1(new_n1019), .C2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g601(.A(new_n1004), .B(new_n1006), .Z(new_n1027));
  NOR2_X1   g602(.A1(new_n1016), .A2(new_n1011), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1011), .B(new_n979), .C1(new_n884), .C2(new_n492), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n984), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  AOI22_X1  g606(.A1(new_n1031), .A2(new_n1008), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1032));
  INV_X1    g607(.A(G8), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1027), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n984), .B(new_n979), .C1(new_n884), .C2(new_n893), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n579), .A2(new_n584), .A3(G1976), .A4(new_n585), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n1035), .A2(G8), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G1976), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT52), .B1(G288), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(G1981), .B1(new_n589), .B2(new_n592), .ZN(new_n1040));
  INV_X1    g615(.A(G61), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1041), .B1(new_n508), .B2(new_n509), .ZN(new_n1042));
  INV_X1    g617(.A(new_n591), .ZN(new_n1043));
  OAI21_X1  g618(.A(G651), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1981), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1044), .A2(new_n1045), .A3(new_n587), .A4(new_n588), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1040), .A2(KEYINPUT49), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT49), .B1(new_n1040), .B2(new_n1046), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1033), .B1(new_n1016), .B2(new_n984), .ZN(new_n1050));
  AOI22_X1  g625(.A1(new_n1037), .A2(new_n1039), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1035), .A2(G8), .A3(new_n1036), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT116), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1035), .A2(new_n1054), .A3(new_n1036), .A4(G8), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1053), .A2(KEYINPUT52), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1051), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1057), .B1(new_n1051), .B2(new_n1056), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1026), .B(new_n1034), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1013), .A2(new_n1018), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n985), .A2(G2084), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n985), .B1(new_n980), .B2(new_n981), .ZN(new_n1064));
  INV_X1    g639(.A(G164), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1065), .A2(KEYINPUT118), .A3(KEYINPUT45), .A4(new_n979), .ZN(new_n1066));
  OAI211_X1 g641(.A(KEYINPUT45), .B(new_n979), .C1(new_n884), .C2(new_n492), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT118), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1064), .A2(new_n1066), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n794), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1063), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1072), .A2(G8), .A3(G168), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT119), .B1(new_n1060), .B2(new_n1073), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1029), .A2(new_n984), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n980), .A2(KEYINPUT50), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1075), .A2(new_n1008), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1024), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1007), .B1(G8), .B2(new_n1078), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1053), .A2(KEYINPUT52), .A3(new_n1055), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT117), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1051), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1079), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1073), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1086), .A2(new_n1087), .A3(new_n1026), .A4(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT63), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1074), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(G8), .B1(new_n1019), .B2(new_n1025), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n1027), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1080), .A2(new_n1083), .A3(new_n1090), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1088), .A2(new_n1093), .A3(new_n1026), .A4(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1091), .A2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(G299), .B(KEYINPUT57), .ZN(new_n1097));
  AOI21_X1  g672(.A(G1956), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1098));
  XNOR2_X1  g673(.A(KEYINPUT56), .B(G2072), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1020), .A2(new_n984), .A3(new_n1021), .A4(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1097), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n1104));
  XNOR2_X1  g679(.A(G299), .B(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(G1956), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1105), .A2(new_n1107), .A3(new_n1100), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1108), .A2(new_n619), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1061), .A2(new_n984), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n800), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1035), .A2(G2067), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1112), .B(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1103), .B1(new_n1109), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1035), .ZN(new_n1117));
  XNOR2_X1  g692(.A(KEYINPUT58), .B(G1341), .ZN(new_n1118));
  OAI22_X1  g693(.A1(new_n1022), .A2(G1996), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n560), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(KEYINPUT59), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1119), .A2(new_n560), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1111), .A2(KEYINPUT60), .A3(new_n618), .A4(new_n1114), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT61), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1102), .A2(new_n1108), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1126), .B1(new_n1102), .B2(new_n1108), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1124), .B(new_n1125), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT60), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n985), .B1(new_n1013), .B2(new_n1018), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1131), .A2(G1348), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1112), .B(KEYINPUT120), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1130), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1114), .B(KEYINPUT60), .C1(G1348), .C2(new_n1131), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1134), .A2(new_n619), .A3(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1116), .B1(new_n1129), .B2(new_n1136), .ZN(new_n1137));
  AND3_X1   g712(.A1(G286), .A2(KEYINPUT121), .A3(G8), .ZN(new_n1138));
  AOI21_X1  g713(.A(KEYINPUT121), .B1(G286), .B2(G8), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1138), .A2(new_n1139), .A3(KEYINPUT51), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1061), .A2(new_n1062), .B1(new_n1070), .B2(new_n794), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1140), .B1(new_n1141), .B2(new_n1033), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1143), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1144));
  NAND2_X1  g719(.A1(G286), .A2(G8), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(G286), .A2(KEYINPUT121), .A3(G8), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1147), .A2(KEYINPUT123), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1144), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1150), .B1(new_n1072), .B2(G8), .ZN(new_n1151));
  XNOR2_X1  g726(.A(KEYINPUT122), .B(KEYINPUT51), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1142), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1141), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT54), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT53), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1158), .B1(new_n1022), .B2(G2078), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1158), .A2(G2078), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1064), .A2(new_n1066), .A3(new_n1069), .A4(new_n1160), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1159), .B(new_n1161), .C1(new_n1131), .C2(G1961), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1157), .B1(new_n1163), .B2(G301), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n1160), .A2(G40), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n982), .A2(G160), .A3(new_n1021), .A4(new_n1165), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1159), .B(new_n1166), .C1(new_n1131), .C2(G1961), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(G171), .ZN(new_n1168));
  AOI22_X1  g743(.A1(new_n1153), .A2(new_n1156), .B1(new_n1164), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1060), .ZN(new_n1170));
  OR3_X1    g745(.A1(new_n1167), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1163), .A2(G301), .ZN(new_n1172));
  OAI21_X1  g747(.A(KEYINPUT124), .B1(new_n1167), .B2(G171), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n1171), .B(new_n1157), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1137), .A2(new_n1169), .A3(new_n1170), .A4(new_n1174), .ZN(new_n1175));
  AND2_X1   g750(.A1(new_n1144), .A2(new_n1149), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1176), .B1(new_n1141), .B2(new_n1033), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1152), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1072), .A2(G8), .ZN(new_n1179));
  AOI22_X1  g754(.A1(new_n1177), .A2(new_n1178), .B1(new_n1179), .B2(new_n1140), .ZN(new_n1180));
  OAI21_X1  g755(.A(KEYINPUT62), .B1(new_n1180), .B2(new_n1155), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT62), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1153), .A2(new_n1182), .A3(new_n1156), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1181), .A2(new_n1170), .A3(new_n1183), .A4(new_n1172), .ZN(new_n1184));
  NOR3_X1   g759(.A1(new_n1026), .A2(new_n1080), .A3(new_n1083), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1082), .A2(new_n1038), .A3(new_n716), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(new_n1046), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1185), .B1(new_n1050), .B2(new_n1187), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1096), .A2(new_n1175), .A3(new_n1184), .A4(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n601), .B(new_n736), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n986), .B1(new_n1000), .B2(new_n1190), .ZN(new_n1191));
  AND3_X1   g766(.A1(new_n1189), .A2(KEYINPUT125), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(KEYINPUT125), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1002), .B1(new_n1192), .B2(new_n1193), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g769(.A(G319), .B1(new_n689), .B2(new_n690), .ZN(new_n1196));
  AOI21_X1  g770(.A(new_n1196), .B1(new_n708), .B2(new_n712), .ZN(new_n1197));
  OAI21_X1  g771(.A(new_n1197), .B1(new_n668), .B2(new_n669), .ZN(new_n1198));
  INV_X1    g772(.A(KEYINPUT126), .ZN(new_n1199));
  NAND2_X1  g773(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  OAI211_X1 g774(.A(new_n1197), .B(KEYINPUT126), .C1(new_n669), .C2(new_n668), .ZN(new_n1201));
  AND4_X1   g775(.A1(new_n901), .A2(new_n968), .A3(new_n1200), .A4(new_n1201), .ZN(G308));
  NAND4_X1  g776(.A1(new_n968), .A2(new_n901), .A3(new_n1200), .A4(new_n1201), .ZN(G225));
endmodule


