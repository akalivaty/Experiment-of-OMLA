//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1204, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  INV_X1    g0009(.A(G77), .ZN(new_n210));
  INV_X1    g0010(.A(G244), .ZN(new_n211));
  INV_X1    g0011(.A(G97), .ZN(new_n212));
  INV_X1    g0012(.A(G257), .ZN(new_n213));
  OAI22_X1  g0013(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT65), .Z(new_n216));
  AOI211_X1 g0016(.A(new_n214), .B(new_n216), .C1(G50), .C2(G226), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G116), .A2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n217), .B(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AND2_X1   g0021(.A1(G68), .A2(G238), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n206), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT64), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n209), .B(new_n224), .C1(new_n227), .C2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  AND2_X1   g0047(.A1(KEYINPUT67), .A2(G1), .ZN(new_n248));
  NOR2_X1   g0048(.A1(KEYINPUT67), .A2(G1), .ZN(new_n249));
  OAI211_X1 g0049(.A(G13), .B(G20), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  OAI21_X1  g0050(.A(G33), .B1(new_n248), .B2(new_n249), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n225), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  AND3_X1   g0054(.A1(new_n250), .A2(new_n251), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G107), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT86), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n257), .B(KEYINPUT25), .C1(new_n250), .C2(G107), .ZN(new_n258));
  INV_X1    g0058(.A(new_n250), .ZN(new_n259));
  INV_X1    g0059(.A(G107), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(KEYINPUT25), .ZN(new_n261));
  OR2_X1    g0061(.A1(new_n257), .A2(KEYINPUT25), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n259), .A2(new_n260), .A3(new_n261), .A4(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n256), .A2(new_n258), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT87), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n256), .A2(KEYINPUT87), .A3(new_n258), .A4(new_n263), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT3), .B(G33), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(new_n226), .A3(G87), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT22), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT23), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n272), .B1(new_n226), .B2(G107), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n260), .A2(KEYINPUT23), .A3(G20), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n270), .A2(new_n271), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  NOR3_X1   g0076(.A1(new_n276), .A2(KEYINPUT72), .A3(G33), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT3), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT72), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n280), .B1(new_n278), .B2(KEYINPUT3), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n277), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n282), .A2(KEYINPUT22), .A3(new_n226), .A4(G87), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n226), .A2(G33), .A3(G116), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n275), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT24), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n275), .A2(new_n283), .A3(KEYINPUT24), .A4(new_n284), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(new_n253), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n268), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n280), .A2(new_n278), .A3(KEYINPUT3), .ZN(new_n291));
  INV_X1    g0091(.A(G1698), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n220), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(KEYINPUT72), .B1(new_n276), .B2(G33), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n276), .A2(G33), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n291), .B(new_n293), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n292), .A2(G257), .ZN(new_n297));
  INV_X1    g0097(.A(G294), .ZN(new_n298));
  OAI22_X1  g0098(.A1(new_n296), .A2(new_n297), .B1(new_n278), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT88), .ZN(new_n300));
  INV_X1    g0100(.A(G41), .ZN(new_n301));
  OAI211_X1 g0101(.A(G1), .B(G13), .C1(new_n278), .C2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT88), .ZN(new_n304));
  OAI221_X1 g0104(.A(new_n304), .B1(new_n278), .B2(new_n298), .C1(new_n296), .C2(new_n297), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n300), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G45), .ZN(new_n307));
  OR2_X1    g0107(.A1(KEYINPUT67), .A2(G1), .ZN(new_n308));
  NAND2_X1  g0108(.A1(KEYINPUT67), .A2(G1), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT5), .B(G41), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n310), .A2(G274), .A3(new_n311), .A4(new_n302), .ZN(new_n312));
  INV_X1    g0112(.A(new_n311), .ZN(new_n313));
  OAI21_X1  g0113(.A(G45), .B1(new_n248), .B2(new_n249), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n302), .B(G264), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n306), .A2(new_n312), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G169), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G179), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n306), .A2(new_n319), .A3(new_n312), .A4(new_n315), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n290), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT89), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT89), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n290), .A2(new_n318), .A3(new_n323), .A4(new_n320), .ZN(new_n324));
  NOR3_X1   g0124(.A1(new_n316), .A2(KEYINPUT90), .A3(G190), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n325), .A2(new_n290), .ZN(new_n326));
  INV_X1    g0126(.A(G200), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n316), .A2(new_n327), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n328), .B(KEYINPUT90), .C1(G190), .C2(new_n316), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n322), .A2(new_n324), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n248), .A2(new_n249), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n253), .B1(new_n332), .B2(G20), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G50), .ZN(new_n334));
  XNOR2_X1  g0134(.A(KEYINPUT8), .B(G58), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n226), .A2(G33), .ZN(new_n336));
  INV_X1    g0136(.A(G150), .ZN(new_n337));
  NOR2_X1   g0137(.A1(G20), .A2(G33), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  OAI22_X1  g0139(.A1(new_n335), .A2(new_n336), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n340), .B1(G20), .B2(new_n203), .ZN(new_n341));
  OAI221_X1 g0141(.A(new_n334), .B1(G50), .B2(new_n250), .C1(new_n341), .C2(new_n254), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT9), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  XOR2_X1   g0144(.A(new_n344), .B(KEYINPUT70), .Z(new_n345));
  INV_X1    g0145(.A(KEYINPUT10), .ZN(new_n346));
  OAI22_X1  g0146(.A1(new_n248), .A2(new_n249), .B1(G41), .B2(G45), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT68), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT68), .ZN(new_n349));
  OAI221_X1 g0149(.A(new_n349), .B1(G41), .B2(G45), .C1(new_n248), .C2(new_n249), .ZN(new_n350));
  AND3_X1   g0150(.A1(new_n348), .A2(new_n302), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G226), .ZN(new_n352));
  INV_X1    g0152(.A(G1), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT66), .B(G45), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n353), .B(G274), .C1(new_n354), .C2(G41), .ZN(new_n355));
  NOR2_X1   g0155(.A1(G222), .A2(G1698), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n292), .A2(G223), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n269), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n358), .B(new_n303), .C1(G77), .C2(new_n269), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n352), .A2(new_n355), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G200), .ZN(new_n361));
  XOR2_X1   g0161(.A(new_n361), .B(KEYINPUT71), .Z(new_n362));
  INV_X1    g0162(.A(new_n360), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n363), .A2(G190), .B1(new_n343), .B2(new_n342), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n345), .A2(new_n346), .A3(new_n362), .A4(new_n364), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n345), .A2(new_n364), .A3(new_n361), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n365), .B1(new_n366), .B2(new_n346), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n363), .A2(new_n319), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n360), .A2(new_n317), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n368), .A2(new_n342), .A3(new_n369), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n348), .A2(new_n350), .A3(G232), .A4(new_n302), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n355), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n281), .A2(new_n279), .ZN(new_n374));
  OR2_X1    g0174(.A1(G223), .A2(G1698), .ZN(new_n375));
  OR2_X1    g0175(.A1(new_n292), .A2(G226), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n374), .A2(new_n291), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(G33), .A2(G87), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n302), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n327), .B1(new_n373), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n377), .A2(new_n378), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n303), .ZN(new_n382));
  INV_X1    g0182(.A(G190), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n382), .A2(new_n383), .A3(new_n372), .A4(new_n355), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(G58), .ZN(new_n386));
  INV_X1    g0186(.A(G68), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(G20), .B1(new_n388), .B2(new_n201), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n338), .A2(G159), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(G20), .B1(new_n374), .B2(new_n291), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT7), .ZN(new_n394));
  OAI21_X1  g0194(.A(G68), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n291), .B1(new_n294), .B2(new_n295), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n226), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n397), .A2(KEYINPUT7), .ZN(new_n398));
  OAI211_X1 g0198(.A(KEYINPUT16), .B(new_n392), .C1(new_n395), .C2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT16), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n394), .B1(new_n269), .B2(G20), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n276), .A2(G33), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n279), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n403), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n387), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n400), .B1(new_n405), .B2(new_n391), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n399), .A2(new_n253), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n250), .A2(new_n335), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n333), .B2(new_n335), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n385), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n410), .B(KEYINPUT17), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT18), .ZN(new_n412));
  INV_X1    g0212(.A(new_n409), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n387), .B1(new_n397), .B2(KEYINPUT7), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n393), .A2(new_n394), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n391), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n254), .B1(new_n416), .B2(KEYINPUT16), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n413), .B1(new_n417), .B2(new_n406), .ZN(new_n418));
  OAI21_X1  g0218(.A(G169), .B1(new_n373), .B2(new_n379), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n382), .A2(G179), .A3(new_n372), .A4(new_n355), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n412), .B1(new_n418), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n407), .A2(new_n409), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n419), .A2(new_n420), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(KEYINPUT18), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G20), .A2(G77), .ZN(new_n427));
  OR2_X1    g0227(.A1(KEYINPUT15), .A2(G87), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT69), .ZN(new_n429));
  NAND2_X1  g0229(.A1(KEYINPUT15), .A2(G87), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  AND2_X1   g0231(.A1(KEYINPUT15), .A2(G87), .ZN(new_n432));
  NOR2_X1   g0232(.A1(KEYINPUT15), .A2(G87), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT69), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  OAI221_X1 g0235(.A(new_n427), .B1(new_n339), .B2(new_n335), .C1(new_n435), .C2(new_n336), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n436), .A2(new_n253), .B1(new_n210), .B2(new_n259), .ZN(new_n437));
  INV_X1    g0237(.A(new_n333), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n437), .B1(new_n210), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(G232), .A2(G1698), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n292), .A2(G238), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n269), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n442), .B(new_n303), .C1(G107), .C2(new_n269), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n348), .A2(new_n302), .A3(new_n350), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n443), .B(new_n355), .C1(new_n444), .C2(new_n211), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n445), .A2(G200), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n439), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(new_n383), .B2(new_n445), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n371), .A2(new_n411), .A3(new_n426), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n351), .A2(G238), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n233), .A2(G1698), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(G226), .B2(G1698), .ZN(new_n452));
  OAI22_X1  g0252(.A1(new_n452), .A2(new_n403), .B1(new_n278), .B2(new_n212), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n303), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n450), .A2(new_n355), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT13), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT13), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n450), .A2(new_n454), .A3(new_n457), .A4(new_n355), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G169), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT14), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT14), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n459), .A2(new_n462), .A3(G169), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n461), .B(new_n463), .C1(new_n319), .C2(new_n459), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n387), .A2(G20), .ZN(new_n465));
  OAI221_X1 g0265(.A(new_n465), .B1(new_n336), .B2(new_n210), .C1(new_n339), .C2(new_n202), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n253), .ZN(new_n467));
  XNOR2_X1  g0267(.A(new_n467), .B(KEYINPUT11), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(new_n387), .B2(new_n438), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n250), .A2(G68), .ZN(new_n470));
  XNOR2_X1  g0270(.A(new_n470), .B(KEYINPUT12), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n464), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n445), .A2(new_n317), .ZN(new_n475));
  OR2_X1    g0275(.A1(new_n445), .A2(G179), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n439), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n459), .A2(G200), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n478), .B(new_n472), .C1(new_n383), .C2(new_n459), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n474), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n449), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n310), .A2(G274), .A3(new_n302), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n314), .A2(G250), .A3(new_n302), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT77), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n211), .A2(G1698), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(G238), .B2(G1698), .ZN(new_n487));
  INV_X1    g0287(.A(G116), .ZN(new_n488));
  OAI22_X1  g0288(.A1(new_n396), .A2(new_n487), .B1(new_n278), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n303), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT77), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n482), .A2(new_n483), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n485), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n317), .ZN(new_n494));
  OR2_X1    g0294(.A1(new_n493), .A2(G179), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n431), .A2(new_n434), .A3(KEYINPUT79), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT79), .B1(new_n431), .B2(new_n434), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n255), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT80), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT79), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n435), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n431), .A2(new_n434), .A3(KEYINPUT79), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT80), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n503), .A2(new_n504), .A3(new_n255), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT81), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n282), .A2(new_n226), .A3(G68), .ZN(new_n508));
  NOR3_X1   g0308(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n509), .A2(KEYINPUT78), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n509), .A2(KEYINPUT78), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT19), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n512), .A2(new_n278), .A3(new_n212), .ZN(new_n513));
  OAI22_X1  g0313(.A1(new_n510), .A2(new_n511), .B1(G20), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n512), .B1(new_n336), .B2(new_n212), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n508), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n516), .A2(new_n253), .B1(new_n259), .B2(new_n435), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n506), .A2(new_n507), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n507), .B1(new_n506), .B2(new_n517), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n494), .B(new_n495), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n255), .A2(G87), .ZN(new_n522));
  XNOR2_X1  g0322(.A(new_n522), .B(KEYINPUT82), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n523), .A2(new_n517), .ZN(new_n524));
  OR3_X1    g0324(.A1(new_n493), .A2(KEYINPUT83), .A3(new_n383), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n493), .A2(G200), .ZN(new_n526));
  OAI21_X1  g0326(.A(KEYINPUT83), .B1(new_n493), .B2(new_n383), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n524), .A2(new_n525), .A3(new_n526), .A4(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n521), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n403), .A2(G303), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n374), .B(new_n291), .C1(G257), .C2(G1698), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n292), .A2(G264), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n303), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n302), .B(G270), .C1(new_n313), .C2(new_n314), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT84), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n535), .A2(new_n312), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n536), .B1(new_n535), .B2(new_n312), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n534), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G200), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n250), .A2(G116), .ZN(new_n541));
  AND4_X1   g0341(.A1(G116), .A2(new_n250), .A3(new_n251), .A4(new_n254), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G283), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n543), .B(new_n226), .C1(G33), .C2(new_n212), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n544), .B(new_n253), .C1(new_n226), .C2(G116), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT20), .ZN(new_n546));
  OAI21_X1  g0346(.A(KEYINPUT85), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n546), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n545), .A2(KEYINPUT85), .A3(new_n546), .ZN(new_n550));
  AOI211_X1 g0350(.A(new_n541), .B(new_n542), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n540), .B(new_n551), .C1(new_n383), .C2(new_n539), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT21), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n539), .A2(G169), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n553), .B1(new_n554), .B2(new_n551), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n541), .B1(new_n549), .B2(new_n550), .ZN(new_n556));
  INV_X1    g0356(.A(new_n542), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n558), .A2(KEYINPUT21), .A3(G169), .A4(new_n539), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n534), .B(G179), .C1(new_n537), .C2(new_n538), .ZN(new_n560));
  OR2_X1    g0360(.A1(new_n551), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n552), .A2(new_n555), .A3(new_n559), .A4(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n529), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n250), .A2(G97), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n564), .B1(new_n255), .B2(G97), .ZN(new_n565));
  NOR3_X1   g0365(.A1(new_n269), .A2(new_n394), .A3(G20), .ZN(new_n566));
  AOI21_X1  g0366(.A(KEYINPUT7), .B1(new_n403), .B2(new_n226), .ZN(new_n567));
  OAI21_X1  g0367(.A(G107), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n260), .A2(KEYINPUT6), .A3(G97), .ZN(new_n569));
  AND2_X1   g0369(.A1(G97), .A2(G107), .ZN(new_n570));
  NOR2_X1   g0370(.A1(G97), .A2(G107), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n569), .B1(new_n572), .B2(KEYINPUT6), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n573), .A2(G20), .B1(G77), .B2(new_n338), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n568), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(KEYINPUT73), .B1(new_n575), .B2(new_n253), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT73), .ZN(new_n577));
  AOI211_X1 g0377(.A(new_n577), .B(new_n254), .C1(new_n568), .C2(new_n574), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n565), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n211), .A2(G1698), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n291), .B(new_n580), .C1(new_n294), .C2(new_n295), .ZN(new_n581));
  XNOR2_X1  g0381(.A(KEYINPUT74), .B(KEYINPUT4), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n292), .A2(G244), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT4), .ZN(new_n584));
  OAI22_X1  g0384(.A1(new_n583), .A2(new_n584), .B1(new_n220), .B2(new_n292), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n581), .A2(new_n582), .B1(new_n269), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n302), .B1(new_n586), .B2(new_n543), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n302), .B(G257), .C1(new_n313), .C2(new_n314), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n312), .ZN(new_n589));
  OAI21_X1  g0389(.A(KEYINPUT75), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n588), .A2(new_n312), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT75), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n581), .A2(new_n582), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n585), .A2(new_n269), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n593), .A2(new_n543), .A3(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n591), .B(new_n592), .C1(new_n595), .C2(new_n302), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n383), .B1(new_n590), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n587), .A2(new_n589), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n598), .A2(new_n327), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n579), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n590), .A2(new_n596), .A3(new_n317), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n598), .A2(new_n319), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n579), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT76), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n579), .A2(KEYINPUT76), .A3(new_n601), .A4(new_n602), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n600), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AND4_X1   g0407(.A1(new_n330), .A2(new_n481), .A3(new_n563), .A4(new_n607), .ZN(G372));
  OR2_X1    g0408(.A1(new_n493), .A2(new_n383), .ZN(new_n609));
  AND4_X1   g0409(.A1(new_n517), .A2(new_n609), .A3(new_n526), .A4(new_n523), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n506), .A2(new_n517), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT81), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n612), .A2(new_n518), .B1(new_n317), .B2(new_n493), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n610), .B1(new_n613), .B2(new_n495), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n326), .A2(new_n329), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n321), .A2(new_n555), .A3(new_n559), .A4(new_n561), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n607), .A2(new_n614), .A3(new_n615), .A4(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n613), .A2(KEYINPUT91), .A3(new_n495), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT91), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n521), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n605), .A2(new_n521), .A3(new_n528), .A4(new_n606), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT26), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT26), .ZN(new_n624));
  INV_X1    g0424(.A(new_n603), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n614), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n617), .A2(new_n621), .A3(new_n623), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n481), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n370), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n474), .A2(new_n477), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n630), .A2(new_n411), .A3(new_n479), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n426), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n629), .B1(new_n632), .B2(new_n367), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n628), .A2(new_n633), .ZN(G369));
  NAND3_X1  g0434(.A1(new_n555), .A2(new_n561), .A3(new_n559), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(G13), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n637), .A2(G20), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n332), .A2(new_n638), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n639), .A2(KEYINPUT27), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(KEYINPUT27), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(G213), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(G343), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n636), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n330), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n321), .ZN(new_n648));
  INV_X1    g0448(.A(new_n644), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n330), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n649), .B1(new_n268), .B2(new_n289), .ZN(new_n652));
  OAI22_X1  g0452(.A1(new_n651), .A2(new_n652), .B1(new_n321), .B2(new_n649), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n649), .A2(new_n551), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n635), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n562), .B2(new_n654), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n656), .A2(G330), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n650), .A2(new_n658), .ZN(G399));
  OR3_X1    g0459(.A1(new_n510), .A2(new_n511), .A3(G116), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n207), .A2(new_n301), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(G1), .ZN(new_n662));
  OAI22_X1  g0462(.A1(new_n660), .A2(new_n662), .B1(new_n228), .B2(new_n661), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT28), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n563), .A2(new_n330), .A3(new_n607), .A4(new_n649), .ZN(new_n665));
  INV_X1    g0465(.A(new_n598), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n316), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT92), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n539), .A2(new_n319), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n316), .A2(new_n666), .A3(KEYINPUT92), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n669), .A2(new_n493), .A3(new_n670), .A4(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n560), .A2(new_n493), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n306), .A2(new_n315), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n590), .A2(new_n596), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT30), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n673), .A2(KEYINPUT30), .A3(new_n675), .A4(new_n674), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n672), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n644), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT31), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n680), .A2(KEYINPUT31), .A3(new_n644), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n665), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n685), .A2(G330), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n524), .A2(new_n609), .A3(new_n526), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n521), .A2(new_n625), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT26), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n621), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n622), .A2(KEYINPUT26), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n322), .A2(new_n324), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n636), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n695), .A2(new_n615), .A3(new_n607), .A4(new_n614), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n644), .B1(new_n693), .B2(new_n696), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n697), .A2(KEYINPUT29), .ZN(new_n698));
  AOI21_X1  g0498(.A(KEYINPUT29), .B1(new_n627), .B2(new_n649), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n687), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n664), .B1(new_n701), .B2(G1), .ZN(G364));
  AOI21_X1  g0502(.A(new_n662), .B1(G45), .B2(new_n638), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n657), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(G330), .B2(new_n656), .ZN(new_n705));
  INV_X1    g0505(.A(new_n703), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n396), .A2(new_n207), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT93), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n243), .A2(G45), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n708), .B(new_n709), .C1(new_n229), .C2(new_n354), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n269), .A2(G355), .A3(new_n207), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n710), .B(new_n711), .C1(G116), .C2(new_n207), .ZN(new_n712));
  NOR2_X1   g0512(.A1(G13), .A2(G33), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G20), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n225), .B1(G20), .B2(new_n317), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n712), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n226), .A2(new_n383), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n319), .A2(G200), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n226), .A2(G190), .ZN(new_n723));
  NOR2_X1   g0523(.A1(G179), .A2(G200), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI22_X1  g0526(.A1(G322), .A2(new_n722), .B1(new_n726), .B2(G329), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n403), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n319), .A2(new_n327), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n719), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n728), .B1(G326), .B2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n226), .B1(new_n724), .B2(G190), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G294), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n327), .A2(G179), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n723), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G283), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n729), .A2(new_n723), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  XNOR2_X1  g0541(.A(KEYINPUT33), .B(G317), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n723), .A2(new_n720), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI22_X1  g0544(.A1(new_n741), .A2(new_n742), .B1(new_n744), .B2(G311), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n732), .A2(new_n735), .A3(new_n739), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n719), .A2(new_n736), .ZN(new_n747));
  INV_X1    g0547(.A(G303), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n734), .A2(KEYINPUT95), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n734), .A2(KEYINPUT95), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G97), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n747), .A2(new_n219), .B1(new_n743), .B2(new_n210), .ZN(new_n755));
  AOI211_X1 g0555(.A(new_n403), .B(new_n755), .C1(G58), .C2(new_n722), .ZN(new_n756));
  AOI22_X1  g0556(.A1(G68), .A2(new_n741), .B1(new_n738), .B2(G107), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n731), .A2(G50), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n754), .A2(new_n756), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G159), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n725), .A2(new_n760), .ZN(new_n761));
  XOR2_X1   g0561(.A(KEYINPUT94), .B(KEYINPUT32), .Z(new_n762));
  XNOR2_X1  g0562(.A(new_n761), .B(new_n762), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n746), .A2(new_n749), .B1(new_n759), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(new_n716), .ZN(new_n765));
  INV_X1    g0565(.A(new_n715), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n718), .B(new_n765), .C1(new_n656), .C2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n705), .B1(new_n706), .B2(new_n767), .ZN(G396));
  NAND2_X1  g0568(.A1(new_n627), .A2(new_n649), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n477), .A2(new_n644), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n439), .A2(new_n644), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n448), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n771), .B1(new_n477), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n769), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n627), .A2(new_n649), .A3(new_n774), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(new_n686), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n706), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n775), .A2(new_n713), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n754), .B1(new_n298), .B2(new_n721), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT96), .ZN(new_n783));
  INV_X1    g0583(.A(new_n747), .ZN(new_n784));
  AOI22_X1  g0584(.A1(G107), .A2(new_n784), .B1(new_n741), .B2(G283), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n738), .A2(G87), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(new_n488), .B2(new_n743), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n269), .B(new_n787), .C1(G303), .C2(new_n731), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n783), .A2(new_n785), .A3(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G311), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n725), .A2(new_n790), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n747), .A2(new_n202), .B1(new_n737), .B2(new_n387), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT97), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G143), .A2(new_n722), .B1(new_n744), .B2(G159), .ZN(new_n795));
  INV_X1    g0595(.A(G137), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n795), .B1(new_n796), .B2(new_n730), .C1(new_n337), .C2(new_n740), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT34), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n396), .B1(new_n797), .B2(new_n798), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n726), .A2(G132), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n792), .A2(new_n793), .B1(G58), .B2(new_n734), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n799), .A2(new_n800), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n789), .A2(new_n791), .B1(new_n794), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n716), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n716), .A2(new_n713), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(new_n210), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n781), .A2(new_n703), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n780), .A2(new_n808), .ZN(G384));
  INV_X1    g0609(.A(KEYINPUT38), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n417), .B1(KEYINPUT16), .B2(new_n416), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n642), .B1(new_n811), .B2(new_n409), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(new_n411), .B2(new_n426), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT37), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n399), .A2(new_n253), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n414), .A2(new_n415), .ZN(new_n817));
  AOI21_X1  g0617(.A(KEYINPUT16), .B1(new_n817), .B2(new_n392), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n642), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n819), .A2(new_n413), .B1(new_n424), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n815), .B1(new_n821), .B2(new_n410), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n421), .A2(new_n642), .B1(new_n407), .B2(new_n409), .ZN(new_n823));
  AND3_X1   g0623(.A1(new_n385), .A2(new_n407), .A3(new_n409), .ZN(new_n824));
  NOR3_X1   g0624(.A1(new_n823), .A2(new_n824), .A3(KEYINPUT37), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n810), .B1(new_n814), .B2(new_n826), .ZN(new_n827));
  AND3_X1   g0627(.A1(new_n423), .A2(KEYINPUT18), .A3(new_n424), .ZN(new_n828));
  AOI21_X1  g0628(.A(KEYINPUT18), .B1(new_n423), .B2(new_n424), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n418), .A2(KEYINPUT17), .A3(new_n385), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT17), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n410), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n812), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n811), .A2(new_n409), .B1(new_n421), .B2(new_n642), .ZN(new_n836));
  OAI21_X1  g0636(.A(KEYINPUT37), .B1(new_n836), .B2(new_n824), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n423), .A2(new_n424), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n423), .A2(new_n820), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n838), .A2(new_n839), .A3(new_n815), .A4(new_n410), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n835), .A2(new_n841), .A3(KEYINPUT38), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n827), .A2(KEYINPUT99), .A3(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT99), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n844), .B(new_n810), .C1(new_n814), .C2(new_n826), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n473), .A2(new_n644), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n479), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n462), .B1(new_n459), .B2(G169), .ZN(new_n848));
  AOI211_X1 g0648(.A(KEYINPUT14), .B(new_n317), .C1(new_n456), .C2(new_n458), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n459), .A2(new_n319), .ZN(new_n850));
  NOR3_X1   g0650(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n847), .B1(new_n851), .B2(new_n472), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n464), .A2(new_n473), .A3(new_n649), .ZN(new_n853));
  AND3_X1   g0653(.A1(new_n852), .A2(new_n853), .A3(new_n774), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n843), .A2(new_n685), .A3(new_n845), .A4(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT40), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XOR2_X1   g0657(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n858));
  AOI21_X1  g0658(.A(new_n839), .B1(new_n411), .B2(new_n426), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT37), .B1(new_n823), .B2(new_n824), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n860), .A2(new_n840), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n858), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n856), .B1(new_n862), .B2(new_n842), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n863), .A2(new_n685), .A3(new_n854), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n857), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT102), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n865), .B(new_n866), .ZN(new_n867));
  XOR2_X1   g0667(.A(new_n867), .B(KEYINPUT103), .Z(new_n868));
  NAND2_X1  g0668(.A1(new_n481), .A2(new_n685), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n868), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(G330), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n698), .A2(new_n699), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n481), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n633), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n871), .B(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n852), .A2(new_n853), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(new_n777), .B2(new_n770), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(new_n845), .A3(new_n843), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n843), .A2(KEYINPUT39), .A3(new_n845), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT39), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n862), .A2(new_n880), .A3(new_n842), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n853), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n830), .A2(new_n642), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n878), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT101), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n878), .A2(new_n884), .A3(KEYINPUT101), .A4(new_n885), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n875), .B(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n332), .B2(new_n638), .ZN(new_n892));
  OAI211_X1 g0692(.A(G116), .B(new_n227), .C1(new_n573), .C2(KEYINPUT35), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n893), .B(KEYINPUT98), .Z(new_n894));
  NAND2_X1  g0694(.A1(new_n573), .A2(KEYINPUT35), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n896), .B(KEYINPUT36), .ZN(new_n897));
  OAI21_X1  g0697(.A(G77), .B1(new_n386), .B2(new_n387), .ZN(new_n898));
  OAI22_X1  g0698(.A1(new_n898), .A2(new_n228), .B1(G50), .B2(new_n387), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n899), .A2(new_n637), .A3(new_n331), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n892), .A2(new_n897), .A3(new_n900), .ZN(G367));
  OR2_X1    g0701(.A1(new_n524), .A2(new_n649), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n614), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n621), .B2(new_n902), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT43), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n905), .B(KEYINPUT105), .Z(new_n906));
  NAND2_X1  g0706(.A1(new_n579), .A2(new_n644), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n607), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n603), .B2(new_n649), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n647), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(KEYINPUT42), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n909), .A2(new_n322), .A3(new_n324), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n605), .A2(new_n606), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n644), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n906), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n909), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n658), .A2(new_n916), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n915), .B(new_n917), .Z(new_n918));
  XOR2_X1   g0718(.A(new_n904), .B(KEYINPUT104), .Z(new_n919));
  NOR2_X1   g0719(.A1(new_n919), .A2(KEYINPUT43), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n918), .B(new_n920), .Z(new_n921));
  XOR2_X1   g0721(.A(new_n661), .B(KEYINPUT41), .Z(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n646), .B1(new_n653), .B2(new_n645), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n657), .A2(KEYINPUT106), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n924), .B(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n700), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT107), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n650), .A2(new_n909), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT45), .Z(new_n930));
  NOR2_X1   g0730(.A1(new_n650), .A2(new_n909), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT44), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n930), .A2(new_n658), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n658), .B1(new_n930), .B2(new_n932), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n928), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n923), .B1(new_n936), .B2(new_n701), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n353), .B1(new_n638), .B2(G45), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n921), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n708), .ZN(new_n941));
  OAI221_X1 g0741(.A(new_n717), .B1(new_n207), .B2(new_n435), .C1(new_n941), .C2(new_n239), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n703), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT108), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n722), .A2(G303), .B1(new_n734), .B2(G107), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n738), .A2(G97), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n945), .B(new_n946), .C1(new_n298), .C2(new_n740), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(G317), .B2(new_n726), .ZN(new_n948));
  AOI22_X1  g0748(.A1(G311), .A2(new_n731), .B1(new_n744), .B2(G283), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n784), .A2(G116), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT46), .ZN(new_n951));
  AND4_X1   g0751(.A1(new_n396), .A2(new_n948), .A3(new_n949), .A4(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(G143), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n269), .B1(new_n721), .B2(new_n337), .C1(new_n953), .C2(new_n730), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n753), .A2(G68), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n738), .A2(G77), .ZN(new_n956));
  AOI22_X1  g0756(.A1(G58), .A2(new_n784), .B1(new_n744), .B2(G50), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n954), .B(new_n958), .C1(G159), .C2(new_n741), .ZN(new_n959));
  XNOR2_X1  g0759(.A(KEYINPUT109), .B(G137), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n726), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n952), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n963));
  XNOR2_X1  g0763(.A(new_n962), .B(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n716), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n944), .B1(new_n904), .B2(new_n766), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n940), .A2(new_n966), .ZN(G387));
  INV_X1    g0767(.A(new_n927), .ZN(new_n968));
  INV_X1    g0768(.A(new_n661), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n700), .A2(new_n926), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n784), .A2(G294), .B1(new_n734), .B2(G283), .ZN(new_n972));
  AOI22_X1  g0772(.A1(G322), .A2(new_n731), .B1(new_n741), .B2(G311), .ZN(new_n973));
  INV_X1    g0773(.A(G317), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n973), .B1(new_n748), .B2(new_n743), .C1(new_n974), .C2(new_n721), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT48), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n972), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT112), .Z(new_n978));
  NAND2_X1  g0778(.A1(new_n975), .A2(new_n976), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT49), .ZN(new_n981));
  AOI22_X1  g0781(.A1(G116), .A2(new_n738), .B1(new_n726), .B2(G326), .ZN(new_n982));
  AND3_X1   g0782(.A1(new_n981), .A2(new_n396), .A3(new_n982), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n721), .A2(new_n202), .B1(new_n743), .B2(new_n387), .ZN(new_n984));
  INV_X1    g0784(.A(new_n503), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n985), .A2(new_n752), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n984), .B(new_n986), .C1(G159), .C2(new_n731), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n210), .B2(new_n747), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n725), .A2(new_n337), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n946), .B1(new_n335), .B2(new_n740), .ZN(new_n990));
  NOR4_X1   g0790(.A1(new_n988), .A2(new_n396), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n716), .B1(new_n983), .B2(new_n991), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n653), .A2(new_n766), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n660), .A2(new_n207), .A3(new_n269), .ZN(new_n994));
  AOI211_X1 g0794(.A(G45), .B(new_n660), .C1(G68), .C2(G77), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT111), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n335), .A2(G50), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT50), .Z(new_n998));
  NOR2_X1   g0798(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n354), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n708), .B1(new_n236), .B2(new_n1000), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n994), .B1(G107), .B2(new_n207), .C1(new_n999), .C2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n717), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n992), .A2(new_n703), .A3(new_n993), .A4(new_n1003), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n971), .B(new_n1004), .C1(new_n938), .C2(new_n926), .ZN(G393));
  OAI211_X1 g0805(.A(new_n936), .B(new_n969), .C1(new_n935), .C2(new_n927), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n730), .A2(new_n337), .B1(new_n721), .B2(new_n760), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT51), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1008), .B(new_n282), .C1(new_n953), .C2(new_n725), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n753), .A2(G77), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n740), .A2(new_n202), .B1(new_n743), .B2(new_n335), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1011), .A2(KEYINPUT114), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(KEYINPUT114), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1010), .A2(new_n786), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1009), .B(new_n1014), .C1(G68), .C2(new_n784), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n730), .A2(new_n974), .B1(new_n721), .B2(new_n790), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT52), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n726), .A2(G322), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n784), .A2(G283), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n740), .A2(new_n748), .B1(new_n743), .B2(new_n298), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(G116), .B2(new_n734), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .A4(new_n1021), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n269), .B(new_n1022), .C1(G107), .C2(new_n738), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n716), .B1(new_n1015), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n717), .B1(new_n212), .B2(new_n207), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n708), .B2(new_n246), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT113), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1024), .A2(new_n703), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n916), .B2(new_n715), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n935), .B2(new_n939), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1006), .A2(new_n1030), .ZN(G390));
  NAND3_X1  g0831(.A1(new_n879), .A2(new_n713), .A3(new_n881), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n747), .A2(new_n337), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT53), .ZN(new_n1034));
  XOR2_X1   g0834(.A(KEYINPUT54), .B(G143), .Z(new_n1035));
  AOI22_X1  g0835(.A1(new_n1033), .A2(new_n1034), .B1(new_n744), .B2(new_n1035), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n741), .A2(new_n960), .B1(new_n726), .B2(G125), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n403), .B1(new_n731), .B2(G128), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n753), .A2(G159), .B1(G50), .B2(new_n738), .ZN(new_n1040));
  INV_X1    g0840(.A(G132), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1040), .B1(new_n1041), .B2(new_n721), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1033), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1039), .B(new_n1042), .C1(KEYINPUT53), .C2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n731), .A2(G283), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1010), .B(new_n1045), .C1(new_n212), .C2(new_n743), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n219), .A2(new_n747), .B1(new_n740), .B2(new_n260), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n403), .B1(new_n721), .B2(new_n488), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n737), .A2(new_n387), .B1(new_n725), .B2(new_n298), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT116), .ZN(new_n1050));
  NOR4_X1   g0850(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .A4(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n716), .B1(new_n1044), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n806), .A2(new_n335), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1032), .A2(new_n703), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n686), .A2(new_n854), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n777), .A2(new_n770), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n876), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n882), .B1(new_n1059), .B2(new_n853), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n862), .A2(new_n842), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n853), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n696), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n690), .B(new_n621), .C1(KEYINPUT26), .C2(new_n622), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n649), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n773), .A2(new_n477), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n770), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1062), .B1(new_n1068), .B2(new_n1058), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1056), .B1(new_n1060), .B2(new_n1069), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n879), .B(new_n881), .C1(new_n877), .C2(new_n883), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n771), .B1(new_n697), .B2(new_n1066), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1072), .A2(new_n876), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1071), .B(new_n1055), .C1(new_n1073), .C2(new_n1062), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1070), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1054), .B1(new_n1075), .B2(new_n938), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n481), .A2(G330), .A3(new_n685), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n873), .A2(new_n633), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n685), .A2(G330), .A3(new_n774), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n686), .A2(new_n854), .B1(new_n1081), .B2(new_n876), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1057), .ZN(new_n1083));
  OAI21_X1  g0883(.A(KEYINPUT115), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1082), .A2(new_n1072), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1081), .A2(new_n876), .ZN(new_n1087));
  AND4_X1   g0887(.A1(KEYINPUT115), .A2(new_n1055), .A3(new_n1072), .A4(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1080), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n969), .B1(new_n1091), .B2(new_n1075), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1090), .A2(new_n1080), .B1(new_n1070), .B2(new_n1074), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1077), .B1(new_n1092), .B2(new_n1093), .ZN(G378));
  AOI21_X1  g0894(.A(new_n1088), .B1(new_n1085), .B2(new_n1084), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1080), .B1(new_n1075), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT120), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n857), .A2(G330), .A3(new_n864), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT119), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n857), .A2(new_n864), .A3(KEYINPUT119), .A4(G330), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n342), .A2(new_n820), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n371), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1102), .B1(new_n367), .B2(new_n370), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1103), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1106), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n367), .A2(new_n370), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1102), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1108), .B1(new_n1111), .B2(new_n1104), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1100), .A2(new_n1101), .A3(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1098), .A2(new_n1099), .A3(new_n1113), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n890), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1115), .A2(new_n888), .A3(new_n889), .A4(new_n1116), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1097), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(KEYINPUT120), .B1(new_n1117), .B2(new_n890), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1096), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT57), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  AND4_X1   g0924(.A1(new_n888), .A2(new_n1115), .A3(new_n889), .A4(new_n1116), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1115), .A2(new_n1116), .B1(new_n888), .B2(new_n889), .ZN(new_n1126));
  OAI211_X1 g0926(.A(KEYINPUT57), .B(new_n1096), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n969), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1124), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1114), .A2(new_n713), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n301), .B1(new_n396), .B2(new_n278), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n202), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n722), .A2(G107), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n503), .A2(new_n744), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(G116), .A2(new_n731), .B1(new_n738), .B2(G58), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n955), .A2(new_n1134), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(G97), .A2(new_n741), .B1(new_n726), .B2(G283), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1138), .B(new_n301), .C1(new_n210), .C2(new_n747), .ZN(new_n1139));
  NOR3_X1   g0939(.A1(new_n1137), .A2(new_n282), .A3(new_n1139), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1035), .A2(new_n784), .B1(new_n722), .B2(G128), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT118), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n753), .A2(G150), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n740), .A2(new_n1041), .B1(new_n743), .B2(new_n796), .ZN(new_n1144));
  XOR2_X1   g0944(.A(new_n1144), .B(KEYINPUT117), .Z(new_n1145));
  NAND2_X1  g0945(.A1(new_n731), .A2(G125), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1142), .A2(new_n1143), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1147), .A2(KEYINPUT59), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n738), .A2(G159), .ZN(new_n1149));
  AOI21_X1  g0949(.A(G41), .B1(new_n726), .B2(G124), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1148), .A2(new_n278), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1147), .A2(KEYINPUT59), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1133), .B1(KEYINPUT58), .B2(new_n1140), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n1140), .A2(KEYINPUT58), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n716), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n806), .A2(new_n202), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1131), .A2(new_n703), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1121), .B1(new_n1158), .B2(KEYINPUT120), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1157), .B1(new_n1159), .B2(new_n938), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(KEYINPUT121), .B1(new_n1130), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1128), .B1(new_n1123), .B2(new_n1122), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT121), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n1163), .A2(new_n1164), .A3(new_n1160), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(G375));
  NAND2_X1  g0967(.A1(new_n1095), .A2(new_n1079), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1091), .A2(new_n922), .A3(new_n1168), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1058), .A2(new_n714), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n986), .B1(G294), .B2(new_n731), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n744), .A2(G107), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n956), .B1(new_n488), .B2(new_n740), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n269), .B(new_n1173), .C1(G283), .C2(new_n722), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n747), .A2(new_n212), .B1(new_n725), .B2(new_n748), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT123), .Z(new_n1176));
  NAND4_X1  g0976(.A1(new_n1171), .A2(new_n1172), .A3(new_n1174), .A4(new_n1176), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(G132), .A2(new_n731), .B1(new_n741), .B2(new_n1035), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n726), .A2(G128), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n722), .A2(new_n960), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(G159), .B2(new_n784), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n738), .A2(G58), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n396), .B1(new_n744), .B2(G150), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n753), .A2(G50), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .A4(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n965), .B1(new_n1177), .B2(new_n1186), .ZN(new_n1187));
  NOR3_X1   g0987(.A1(new_n716), .A2(G68), .A3(new_n713), .ZN(new_n1188));
  NOR4_X1   g0988(.A1(new_n1170), .A2(new_n706), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n938), .B(KEYINPUT122), .Z(new_n1190));
  AOI21_X1  g0990(.A(new_n1189), .B1(new_n1090), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1169), .A2(new_n1191), .ZN(G381));
  INV_X1    g0992(.A(G384), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n1169), .A2(new_n1191), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(G378), .A2(KEYINPUT124), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT124), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1196), .B(new_n1077), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1166), .A2(new_n1193), .A3(new_n1194), .A4(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(G390), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1200), .A2(new_n940), .A3(new_n966), .ZN(new_n1201));
  OR3_X1    g1001(.A1(new_n1201), .A2(G396), .A3(G393), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1199), .A2(new_n1202), .ZN(G407));
  NAND3_X1  g1003(.A1(new_n1166), .A2(new_n643), .A3(new_n1198), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(G407), .A2(G213), .A3(new_n1204), .ZN(G409));
  NAND2_X1  g1005(.A1(new_n643), .A2(G213), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT60), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1168), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1095), .A2(KEYINPUT60), .A3(new_n1079), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1208), .A2(new_n969), .A3(new_n1091), .A4(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n1191), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n1193), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1210), .A2(G384), .A3(new_n1191), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(G378), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1163), .A2(new_n1216), .A3(new_n1160), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n922), .B(new_n1096), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1157), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n1158), .B2(new_n1190), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1195), .A2(new_n1197), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1206), .B(new_n1215), .C1(new_n1217), .C2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(KEYINPUT62), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT61), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1206), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(G2897), .ZN(new_n1226));
  XOR2_X1   g1026(.A(new_n1226), .B(KEYINPUT126), .Z(new_n1227));
  XNOR2_X1  g1027(.A(new_n1214), .B(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1160), .B1(new_n1124), .B2(new_n1129), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1221), .B1(new_n1229), .B2(G378), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1228), .B1(new_n1230), .B2(new_n1225), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1130), .A2(G378), .A3(new_n1161), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1221), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT62), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1234), .A2(new_n1235), .A3(new_n1206), .A4(new_n1215), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1223), .A2(new_n1224), .A3(new_n1231), .A4(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(G387), .A2(G390), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n1201), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(G393), .B(G396), .ZN(new_n1240));
  OR2_X1    g1040(.A1(new_n1240), .A2(KEYINPUT127), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1240), .B(KEYINPUT127), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1243), .A2(new_n1201), .A3(new_n1238), .ZN(new_n1244));
  AND2_X1   g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1237), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT125), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n1230), .B2(new_n1225), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1234), .A2(KEYINPUT125), .A3(new_n1206), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1248), .A2(new_n1228), .A3(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT61), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT63), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1222), .A2(new_n1252), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1234), .A2(KEYINPUT63), .A3(new_n1206), .A4(new_n1215), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1250), .A2(new_n1251), .A3(new_n1253), .A4(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1246), .A2(new_n1255), .ZN(G405));
  INV_X1    g1056(.A(new_n1198), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1232), .B(new_n1214), .C1(new_n1166), .C2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1130), .A2(KEYINPUT121), .A3(new_n1161), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1164), .B1(new_n1163), .B2(new_n1160), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1257), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1215), .B1(new_n1261), .B2(new_n1217), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1258), .A2(new_n1262), .A3(new_n1245), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1245), .B1(new_n1258), .B2(new_n1262), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1263), .A2(new_n1264), .ZN(G402));
endmodule


