//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 0 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1204, new_n1205, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT64), .Z(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  XOR2_X1   g0010(.A(KEYINPUT65), .B(G238), .Z(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(new_n203), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G107), .A2(G264), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n210), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT66), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT1), .ZN(new_n220));
  OR2_X1    g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n220), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n210), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT0), .Z(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n202), .A2(new_n203), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n225), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  AND3_X1   g0032(.A1(new_n221), .A2(new_n222), .A3(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  INV_X1    g0038(.A(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(KEYINPUT2), .B(G226), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n237), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT68), .ZN(new_n247));
  XOR2_X1   g0047(.A(G50), .B(G68), .Z(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(KEYINPUT86), .ZN(new_n252));
  AND2_X1   g0052(.A1(KEYINPUT69), .A2(G41), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT69), .A2(G41), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G45), .ZN(new_n256));
  AOI21_X1  g0056(.A(G1), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G274), .ZN(new_n258));
  AND2_X1   g0058(.A1(G1), .A2(G13), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n257), .A2(KEYINPUT70), .A3(new_n261), .ZN(new_n262));
  OR2_X1    g0062(.A1(KEYINPUT69), .A2(G41), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT69), .A2(G41), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(new_n256), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(new_n261), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT70), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n259), .A2(new_n260), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n262), .A2(new_n269), .B1(G232), .B2(new_n273), .ZN(new_n274));
  AND2_X1   g0074(.A1(KEYINPUT85), .A2(G190), .ZN(new_n275));
  NOR2_X1   g0075(.A1(KEYINPUT85), .A2(G190), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT72), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n270), .B(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G1698), .ZN(new_n280));
  AND2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  OAI211_X1 g0082(.A(G223), .B(new_n280), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G33), .A2(G87), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AND2_X1   g0085(.A1(G226), .A2(G1698), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n286), .B1(new_n281), .B2(new_n282), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT83), .ZN(new_n288));
  OR2_X1    g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT83), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(new_n292), .A3(new_n286), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n285), .B1(new_n288), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT84), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n279), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n293), .A2(new_n288), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n283), .A2(new_n284), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n297), .A2(new_n295), .A3(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n274), .B(new_n277), .C1(new_n296), .C2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(KEYINPUT70), .B1(new_n257), .B2(new_n261), .ZN(new_n301));
  AND4_X1   g0101(.A1(KEYINPUT70), .A2(new_n265), .A3(new_n261), .A4(new_n266), .ZN(new_n302));
  OAI22_X1  g0102(.A1(new_n301), .A2(new_n302), .B1(new_n239), .B2(new_n272), .ZN(new_n303));
  INV_X1    g0103(.A(new_n279), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n297), .A2(new_n298), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n304), .B1(new_n305), .B2(KEYINPUT84), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n294), .A2(new_n295), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n303), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n300), .B1(new_n308), .B2(G200), .ZN(new_n309));
  INV_X1    g0109(.A(G33), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n226), .B1(new_n210), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n311), .B(KEYINPUT73), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n266), .A2(G13), .A3(G20), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT8), .B(G58), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n227), .A2(G1), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n315), .ZN(new_n319));
  OAI22_X1  g0119(.A1(new_n314), .A2(new_n318), .B1(new_n313), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(G58), .A2(G68), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT80), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT80), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n323), .A2(G58), .A3(G68), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n322), .A2(new_n324), .A3(new_n229), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G20), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT81), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n227), .A2(new_n310), .ZN(new_n328));
  INV_X1    g0128(.A(G159), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(G20), .A2(G33), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(KEYINPUT81), .A3(G159), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT82), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n326), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n334), .B1(new_n326), .B2(new_n333), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT16), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n289), .A2(new_n227), .A3(new_n290), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT7), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n289), .A2(KEYINPUT7), .A3(new_n227), .A4(new_n290), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n338), .B1(new_n343), .B2(G68), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n312), .B1(new_n337), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n326), .A2(new_n333), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT82), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n326), .A2(new_n333), .A3(new_n334), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n343), .A2(G68), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n338), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n320), .B1(new_n345), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n309), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT17), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G179), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n356), .B(new_n274), .C1(new_n296), .C2(new_n299), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n308), .B2(G169), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT18), .B1(new_n358), .B2(new_n352), .ZN(new_n359));
  INV_X1    g0159(.A(new_n320), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT16), .B1(new_n337), .B2(new_n349), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n344), .A2(new_n347), .A3(new_n348), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT73), .ZN(new_n363));
  XNOR2_X1  g0163(.A(new_n311), .B(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n360), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n274), .B1(new_n296), .B2(new_n299), .ZN(new_n367));
  INV_X1    g0167(.A(G169), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT18), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n366), .A2(new_n369), .A3(new_n370), .A4(new_n357), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n309), .A2(KEYINPUT17), .A3(new_n352), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n355), .A2(new_n359), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT77), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n319), .A2(new_n331), .B1(G20), .B2(G77), .ZN(new_n375));
  XNOR2_X1  g0175(.A(KEYINPUT15), .B(G87), .ZN(new_n376));
  XNOR2_X1  g0176(.A(new_n376), .B(KEYINPUT74), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n227), .A2(G33), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n375), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G77), .ZN(new_n380));
  INV_X1    g0180(.A(new_n313), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n379), .A2(new_n364), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n316), .A2(new_n380), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n312), .A2(new_n313), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT75), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT75), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n312), .A2(new_n386), .A3(new_n313), .A4(new_n383), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT76), .B1(new_n382), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n281), .A2(new_n282), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT71), .B1(new_n391), .B2(new_n280), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT71), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n291), .A2(new_n393), .A3(G1698), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n211), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n291), .A2(G232), .A3(new_n280), .ZN(new_n396));
  INV_X1    g0196(.A(G107), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n396), .B1(new_n397), .B2(new_n291), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n279), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n262), .A2(new_n269), .ZN(new_n401));
  INV_X1    g0201(.A(G244), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n401), .B1(new_n402), .B2(new_n272), .ZN(new_n403));
  OAI21_X1  g0203(.A(G200), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n382), .A2(new_n388), .A3(KEYINPUT76), .ZN(new_n405));
  INV_X1    g0205(.A(new_n403), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n406), .A2(G190), .A3(new_n399), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n390), .A2(new_n404), .A3(new_n405), .A4(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n368), .B1(new_n400), .B2(new_n403), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n406), .A2(new_n356), .A3(new_n399), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n382), .A2(new_n388), .A3(KEYINPUT76), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n409), .B(new_n410), .C1(new_n411), .C2(new_n389), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n374), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n408), .A2(new_n412), .A3(new_n374), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n373), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT78), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT10), .ZN(new_n418));
  OR2_X1    g0218(.A1(new_n417), .A2(KEYINPUT10), .ZN(new_n419));
  INV_X1    g0219(.A(new_n316), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n312), .A2(G50), .A3(new_n313), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n204), .A2(G20), .ZN(new_n422));
  INV_X1    g0222(.A(G150), .ZN(new_n423));
  OAI221_X1 g0223(.A(new_n422), .B1(new_n423), .B2(new_n328), .C1(new_n315), .C2(new_n378), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n364), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n381), .A2(new_n201), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n421), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n427), .A2(KEYINPUT9), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(KEYINPUT9), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(G190), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n301), .A2(new_n302), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(G226), .B2(new_n273), .ZN(new_n433));
  INV_X1    g0233(.A(G223), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(new_n392), .B2(new_n394), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n291), .A2(new_n280), .ZN(new_n436));
  INV_X1    g0236(.A(G222), .ZN(new_n437));
  OAI22_X1  g0237(.A1(new_n436), .A2(new_n437), .B1(new_n380), .B2(new_n291), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n279), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n433), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n430), .B1(new_n431), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(G200), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n418), .B(new_n419), .C1(new_n441), .C2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n440), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n445), .A2(G190), .B1(new_n429), .B2(new_n428), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n446), .A2(new_n417), .A3(KEYINPUT10), .A4(new_n442), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n440), .A2(new_n368), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n448), .B(new_n427), .C1(G179), .C2(new_n440), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n444), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n416), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n381), .A2(KEYINPUT79), .A3(new_n203), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT12), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT79), .B1(new_n381), .B2(new_n203), .ZN(new_n455));
  XOR2_X1   g0255(.A(new_n454), .B(new_n455), .Z(new_n456));
  INV_X1    g0256(.A(KEYINPUT11), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n331), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(new_n380), .B2(new_n378), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n364), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n456), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n457), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n420), .A2(G68), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(new_n314), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(G1698), .B1(new_n289), .B2(new_n290), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G226), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n291), .A2(G232), .A3(G1698), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G97), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n471), .A2(new_n279), .B1(G238), .B2(new_n273), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT13), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(new_n401), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n473), .B1(new_n472), .B2(new_n401), .ZN(new_n476));
  OAI21_X1  g0276(.A(G169), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n472), .A2(new_n401), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT13), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n474), .ZN(new_n480));
  OAI22_X1  g0280(.A1(new_n477), .A2(KEYINPUT14), .B1(new_n480), .B2(new_n356), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT14), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n482), .B1(new_n480), .B2(G169), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n466), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(G200), .B1(new_n475), .B2(new_n476), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n479), .A2(G190), .A3(new_n474), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n485), .A2(new_n465), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n252), .B1(new_n452), .B2(new_n489), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n408), .A2(new_n412), .A3(new_n374), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(new_n413), .ZN(new_n492));
  NOR3_X1   g0292(.A1(new_n492), .A2(new_n450), .A3(new_n373), .ZN(new_n493));
  INV_X1    g0293(.A(new_n489), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n493), .A2(KEYINPUT86), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G283), .ZN(new_n497));
  INV_X1    g0297(.A(G97), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n497), .B(new_n227), .C1(G33), .C2(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n499), .B(new_n311), .C1(new_n227), .C2(G116), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT20), .ZN(new_n501));
  XNOR2_X1  g0301(.A(new_n500), .B(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n266), .A2(G33), .ZN(new_n503));
  XNOR2_X1  g0303(.A(new_n503), .B(KEYINPUT88), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n312), .A2(G116), .A3(new_n313), .A4(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n313), .A2(G116), .ZN(new_n506));
  XNOR2_X1  g0306(.A(new_n506), .B(KEYINPUT91), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n502), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n291), .A2(G264), .A3(G1698), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n291), .A2(G257), .A3(new_n280), .ZN(new_n510));
  INV_X1    g0310(.A(G303), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n509), .B(new_n510), .C1(new_n511), .C2(new_n291), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n279), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n266), .A2(G45), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n263), .A2(new_n264), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT5), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(G41), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT5), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n520), .A2(G270), .A3(new_n270), .ZN(new_n521));
  XOR2_X1   g0321(.A(new_n519), .B(KEYINPUT89), .Z(new_n522));
  NAND3_X1  g0322(.A1(new_n522), .A2(new_n261), .A3(new_n517), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n513), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n508), .A2(new_n524), .A3(G169), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT21), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n524), .A2(new_n356), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n508), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n508), .A2(new_n524), .A3(KEYINPUT21), .A4(G169), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n508), .B1(G200), .B2(new_n524), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT92), .ZN(new_n533));
  OR2_X1    g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n277), .ZN(new_n535));
  INV_X1    g0335(.A(new_n524), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n532), .A2(new_n533), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n531), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n291), .A2(new_n227), .A3(G87), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT22), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT22), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n291), .A2(new_n541), .A3(new_n227), .A4(G87), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT23), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n227), .B2(G107), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n397), .A2(KEYINPUT23), .A3(G20), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT93), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G116), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n548), .B1(new_n549), .B2(G20), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n227), .A2(KEYINPUT93), .A3(G33), .A4(G116), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n547), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n543), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT24), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT24), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n543), .A2(new_n555), .A3(new_n552), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n312), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n312), .A2(new_n313), .A3(new_n504), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(new_n397), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n381), .A2(new_n397), .ZN(new_n560));
  XNOR2_X1  g0360(.A(new_n560), .B(KEYINPUT25), .ZN(new_n561));
  OR2_X1    g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(KEYINPUT94), .B1(new_n557), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n556), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n555), .B1(new_n543), .B2(new_n552), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n364), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT94), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n559), .A2(new_n561), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(G250), .ZN(new_n570));
  INV_X1    g0370(.A(G294), .ZN(new_n571));
  OAI22_X1  g0371(.A1(new_n436), .A2(new_n570), .B1(new_n310), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n291), .A2(G257), .A3(G1698), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n279), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n520), .A2(G264), .A3(new_n270), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n575), .A2(new_n576), .A3(new_n523), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G169), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n356), .B2(new_n577), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n563), .A2(new_n569), .A3(new_n579), .ZN(new_n580));
  OR2_X1    g0380(.A1(new_n577), .A2(new_n431), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n577), .A2(G200), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n581), .A2(new_n566), .A3(new_n568), .A4(new_n582), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n291), .A2(new_n227), .A3(G68), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT19), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n227), .B1(new_n470), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(G87), .B2(new_n207), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n586), .B1(new_n378), .B2(new_n498), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n585), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n364), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n377), .A2(new_n381), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n591), .B(new_n592), .C1(new_n558), .C2(new_n377), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n514), .A2(new_n570), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n266), .A2(new_n258), .A3(G45), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n270), .A3(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n291), .A2(G244), .A3(G1698), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n291), .A2(G238), .A3(new_n280), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(new_n599), .A3(new_n549), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n597), .B1(new_n600), .B2(new_n279), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n356), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n593), .B(new_n602), .C1(G169), .C2(new_n601), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n467), .A2(KEYINPUT4), .A3(G244), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n291), .A2(G250), .A3(G1698), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n604), .A2(new_n497), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT4), .B1(new_n467), .B2(G244), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n279), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n520), .A2(G257), .A3(new_n270), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n608), .A2(new_n356), .A3(new_n523), .A4(new_n609), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n604), .A2(new_n497), .A3(new_n605), .ZN(new_n611));
  INV_X1    g0411(.A(new_n607), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n304), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n609), .A2(new_n523), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n368), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n343), .A2(G107), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT87), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n343), .A2(KEYINPUT87), .A3(G107), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n397), .A2(KEYINPUT6), .A3(G97), .ZN(new_n620));
  XOR2_X1   g0420(.A(G97), .B(G107), .Z(new_n621));
  OAI21_X1  g0421(.A(new_n620), .B1(new_n621), .B2(KEYINPUT6), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n622), .A2(G20), .B1(G77), .B2(new_n331), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n618), .A2(new_n619), .A3(new_n623), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n624), .A2(new_n364), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n381), .A2(new_n498), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(new_n558), .B2(new_n498), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n610), .B(new_n615), .C1(new_n625), .C2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n601), .A2(G190), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT90), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT90), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n601), .A2(new_n631), .A3(G190), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n600), .A2(new_n279), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n596), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G200), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n312), .A2(G87), .A3(new_n313), .A4(new_n504), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n636), .A2(new_n591), .A3(new_n592), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n630), .A2(new_n632), .A3(new_n635), .A4(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n627), .B1(new_n624), .B2(new_n364), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n608), .A2(new_n523), .A3(new_n609), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(G200), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n639), .B(new_n641), .C1(new_n431), .C2(new_n640), .ZN(new_n642));
  AND4_X1   g0442(.A1(new_n603), .A2(new_n628), .A3(new_n638), .A4(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n496), .A2(new_n538), .A3(new_n584), .A4(new_n643), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n644), .B(KEYINPUT95), .ZN(G372));
  INV_X1    g0445(.A(new_n449), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n359), .A2(new_n371), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n484), .B1(new_n487), .B2(new_n412), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT96), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n651), .A2(new_n355), .A3(new_n372), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n649), .A2(new_n650), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n648), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n444), .A2(new_n447), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n646), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n496), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n635), .A2(new_n637), .A3(new_n629), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(new_n603), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n628), .A2(new_n642), .A3(new_n660), .A4(new_n583), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n579), .B1(new_n557), .B2(new_n562), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n659), .A2(new_n603), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n615), .A2(new_n610), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n665), .A2(new_n639), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT26), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n638), .A2(new_n603), .ZN(new_n670));
  OAI21_X1  g0470(.A(KEYINPUT26), .B1(new_n628), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n669), .A2(new_n671), .A3(new_n603), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n664), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n657), .B1(new_n658), .B2(new_n674), .ZN(G369));
  INV_X1    g0475(.A(new_n508), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n266), .A2(new_n227), .A3(G13), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n676), .A2(new_n683), .ZN(new_n684));
  MUX2_X1   g0484(.A(new_n538), .B(new_n531), .S(new_n684), .Z(new_n685));
  XOR2_X1   g0485(.A(new_n685), .B(KEYINPUT97), .Z(new_n686));
  NAND3_X1  g0486(.A1(new_n563), .A2(new_n569), .A3(new_n682), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n584), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n580), .B2(new_n683), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n686), .A2(G330), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT98), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n662), .A2(new_n682), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n584), .A2(new_n692), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n691), .B(new_n693), .C1(new_n663), .C2(new_n682), .ZN(G399));
  INV_X1    g0494(.A(new_n223), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(new_n515), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G1), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n230), .B2(new_n697), .ZN(new_n700));
  XOR2_X1   g0500(.A(KEYINPUT99), .B(KEYINPUT28), .Z(new_n701));
  XNOR2_X1  g0501(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT31), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n601), .A2(new_n575), .A3(new_n576), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT100), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n613), .A2(new_n614), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT100), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n601), .A2(new_n575), .A3(new_n576), .A4(new_n707), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n705), .A2(new_n528), .A3(new_n706), .A4(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n709), .A2(KEYINPUT101), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n710), .B1(new_n709), .B2(KEYINPUT101), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n524), .A2(new_n356), .A3(new_n634), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n640), .A2(new_n577), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(KEYINPUT102), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT102), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n640), .A2(new_n716), .A3(new_n577), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n713), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n711), .A2(new_n712), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n703), .B1(new_n719), .B2(new_n683), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n712), .A2(new_n718), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n709), .A2(KEYINPUT101), .A3(new_n710), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(KEYINPUT31), .A3(new_n682), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n584), .A2(new_n643), .A3(new_n538), .A4(new_n683), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n720), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G330), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n580), .A2(new_n662), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT106), .ZN(new_n730));
  INV_X1    g0530(.A(new_n661), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT106), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n580), .A2(new_n662), .A3(new_n732), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n730), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n668), .B1(new_n628), .B2(new_n670), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n666), .A2(new_n639), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n736), .A2(new_n660), .A3(KEYINPUT26), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n735), .A2(KEYINPUT105), .A3(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT105), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n736), .A2(new_n660), .A3(new_n739), .A4(KEYINPUT26), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n738), .A2(new_n603), .A3(new_n740), .ZN(new_n741));
  OAI211_X1 g0541(.A(KEYINPUT29), .B(new_n683), .C1(new_n734), .C2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n683), .B1(new_n664), .B2(new_n672), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT103), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI211_X1 g0545(.A(KEYINPUT103), .B(new_n683), .C1(new_n664), .C2(new_n672), .ZN(new_n746));
  XNOR2_X1  g0546(.A(KEYINPUT104), .B(KEYINPUT29), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n728), .B1(new_n742), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n702), .B1(new_n749), .B2(G1), .ZN(G364));
  INV_X1    g0550(.A(G13), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n266), .B1(new_n752), .B2(G45), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n696), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n695), .A2(new_n391), .ZN(new_n757));
  INV_X1    g0557(.A(G116), .ZN(new_n758));
  AOI22_X1  g0558(.A1(G355), .A2(new_n757), .B1(new_n758), .B2(new_n695), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n250), .A2(new_n256), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n695), .A2(new_n291), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n761), .B1(G45), .B2(new_n230), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n759), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G13), .A2(G33), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT107), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n226), .B1(G20), .B2(new_n368), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n756), .B1(new_n763), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n767), .ZN(new_n770));
  INV_X1    g0570(.A(G200), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n227), .A2(new_n356), .A3(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G190), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n227), .A2(new_n356), .A3(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n431), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n775), .A2(new_n203), .B1(new_n777), .B2(new_n380), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n773), .A2(new_n277), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n535), .A2(new_n776), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n780), .A2(new_n201), .B1(new_n202), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n771), .A2(G179), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n783), .A2(G20), .A3(G190), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G87), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n227), .A2(G190), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n783), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n786), .B(new_n291), .C1(new_n397), .C2(new_n788), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n778), .A2(new_n782), .A3(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n787), .ZN(new_n791));
  OR3_X1    g0591(.A1(KEYINPUT108), .A2(G179), .A3(G200), .ZN(new_n792));
  OAI21_X1  g0592(.A(KEYINPUT108), .B1(G179), .B2(G200), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G159), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT32), .Z(new_n796));
  AOI21_X1  g0596(.A(new_n431), .B1(new_n792), .B2(new_n793), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n227), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n798), .A2(KEYINPUT109), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(KEYINPUT109), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n790), .B(new_n796), .C1(new_n498), .C2(new_n801), .ZN(new_n802));
  XOR2_X1   g0602(.A(KEYINPUT110), .B(G326), .Z(new_n803));
  INV_X1    g0603(.A(G311), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n780), .A2(new_n803), .B1(new_n804), .B2(new_n777), .ZN(new_n805));
  XOR2_X1   g0605(.A(KEYINPUT33), .B(G317), .Z(new_n806));
  INV_X1    g0606(.A(G322), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n775), .A2(new_n806), .B1(new_n807), .B2(new_n781), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(G283), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n391), .B1(new_n788), .B2(new_n810), .C1(new_n511), .C2(new_n784), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(G329), .B2(new_n794), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n809), .B(new_n812), .C1(new_n571), .C2(new_n798), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n802), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n766), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n769), .B1(new_n770), .B2(new_n814), .C1(new_n686), .C2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n686), .A2(G330), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n756), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n686), .A2(G330), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n816), .B1(new_n818), .B2(new_n819), .ZN(G396));
  OAI21_X1  g0620(.A(new_n682), .B1(new_n411), .B2(new_n389), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n408), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n412), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n412), .A2(new_n682), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n745), .A2(new_n746), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n824), .B1(new_n412), .B2(new_n822), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n828), .B(new_n683), .C1(new_n664), .C2(new_n672), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n755), .B1(new_n830), .B2(new_n727), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n727), .B2(new_n830), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n767), .A2(new_n764), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n755), .B1(G77), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n788), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n779), .A2(G303), .B1(G87), .B2(new_n836), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n837), .B1(new_n758), .B2(new_n777), .C1(new_n571), .C2(new_n781), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n774), .B(KEYINPUT111), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n838), .B1(G283), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n794), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n391), .B1(new_n784), .B2(new_n397), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n842), .A2(new_n804), .B1(new_n843), .B2(KEYINPUT112), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(KEYINPUT112), .B2(new_n843), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n841), .B(new_n845), .C1(new_n498), .C2(new_n801), .ZN(new_n846));
  INV_X1    g0646(.A(new_n777), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n779), .A2(G137), .B1(new_n847), .B2(G159), .ZN(new_n848));
  INV_X1    g0648(.A(G143), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n848), .B1(new_n849), .B2(new_n781), .C1(new_n423), .C2(new_n775), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT34), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n836), .A2(G68), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n854), .B(new_n291), .C1(new_n201), .C2(new_n784), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(G132), .B2(new_n794), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n853), .B(new_n856), .C1(new_n202), .C2(new_n798), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n846), .B1(new_n852), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n835), .B1(new_n858), .B2(new_n767), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n828), .B2(new_n765), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n832), .A2(new_n860), .ZN(G384));
  NAND2_X1  g0661(.A1(new_n231), .A2(G77), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n322), .A2(new_n324), .ZN(new_n863));
  OAI22_X1  g0663(.A1(new_n862), .A2(new_n863), .B1(G50), .B2(new_n203), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n864), .A2(G1), .A3(new_n751), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n865), .B(KEYINPUT113), .Z(new_n866));
  INV_X1    g0666(.A(KEYINPUT36), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n228), .A2(G116), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(new_n622), .B2(KEYINPUT35), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(KEYINPUT35), .B2(new_n622), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n866), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n867), .B2(new_n870), .ZN(new_n872));
  INV_X1    g0672(.A(G330), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n466), .A2(new_n682), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n484), .A2(new_n488), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n477), .A2(KEYINPUT14), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n480), .A2(new_n482), .A3(G169), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n876), .B(new_n877), .C1(new_n356), .C2(new_n480), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n466), .B(new_n682), .C1(new_n878), .C2(new_n487), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n826), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n726), .A2(KEYINPUT40), .A3(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT38), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n366), .A2(new_n357), .A3(new_n369), .ZN(new_n883));
  INV_X1    g0683(.A(new_n680), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n366), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n883), .A2(new_n353), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT37), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n883), .A2(new_n353), .A3(new_n885), .A4(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n887), .A2(KEYINPUT115), .A3(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n885), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n373), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT115), .B1(new_n887), .B2(new_n889), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n882), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT116), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT116), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n897), .B(new_n882), .C1(new_n893), .C2(new_n894), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT114), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n892), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n373), .A2(KEYINPUT114), .A3(new_n891), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n887), .A2(new_n889), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n901), .A2(KEYINPUT38), .A3(new_n902), .A4(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n881), .B1(new_n899), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT40), .ZN(new_n906));
  INV_X1    g0706(.A(new_n904), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n892), .A2(new_n900), .B1(new_n887), .B2(new_n889), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT38), .B1(new_n908), .B2(new_n902), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n726), .B(new_n880), .C1(new_n907), .C2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n905), .B1(new_n906), .B2(new_n910), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n496), .A2(new_n726), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n873), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n911), .B2(new_n912), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n879), .A2(new_n875), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n829), .B2(new_n825), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n907), .B2(new_n909), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n647), .A2(new_n680), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT39), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n904), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n898), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT115), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n903), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(new_n892), .A3(new_n890), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n897), .B1(new_n925), .B2(new_n882), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n921), .B1(new_n922), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(KEYINPUT39), .B1(new_n907), .B2(new_n909), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n878), .A2(new_n466), .A3(new_n683), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n919), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n452), .A2(new_n252), .A3(new_n489), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT86), .B1(new_n493), .B2(new_n494), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n748), .B(new_n742), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n935), .A2(new_n657), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n932), .B(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n914), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n266), .B2(new_n752), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n914), .A2(new_n937), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n872), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT117), .ZN(G367));
  INV_X1    g0742(.A(KEYINPUT120), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n628), .B(new_n642), .C1(new_n639), .C2(new_n683), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n736), .A2(new_n682), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n693), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT42), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n628), .B1(new_n944), .B2(new_n580), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n683), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n637), .A2(new_n683), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n660), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n603), .B2(new_n954), .ZN(new_n956));
  XOR2_X1   g0756(.A(KEYINPUT118), .B(KEYINPUT43), .Z(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n952), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT119), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n952), .A2(KEYINPUT119), .A3(new_n958), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n958), .B1(KEYINPUT43), .B2(new_n956), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n951), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n943), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  AOI211_X1 g0767(.A(KEYINPUT120), .B(new_n965), .C1(new_n961), .C2(new_n962), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n691), .A2(new_n946), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  OR3_X1    g0770(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n970), .B1(new_n967), .B2(new_n968), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n696), .B(KEYINPUT41), .Z(new_n973));
  OAI21_X1  g0773(.A(new_n693), .B1(new_n663), .B2(new_n682), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n946), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT44), .Z(new_n976));
  NOR2_X1   g0776(.A1(new_n974), .A2(new_n946), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT45), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n691), .B(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n693), .B1(new_n689), .B2(new_n692), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n817), .B(new_n981), .Z(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n749), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n973), .B1(new_n985), .B2(new_n749), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n971), .B(new_n972), .C1(new_n986), .C2(new_n754), .ZN(new_n987));
  INV_X1    g0787(.A(new_n768), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(new_n236), .B2(new_n761), .ZN(new_n989));
  INV_X1    g0789(.A(new_n377), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n695), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n756), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n781), .A2(new_n511), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n784), .A2(new_n758), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n780), .A2(new_n804), .B1(new_n994), .B2(KEYINPUT46), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n993), .B(new_n995), .C1(KEYINPUT46), .C2(new_n994), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n391), .B1(new_n788), .B2(new_n498), .C1(new_n777), .C2(new_n810), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G317), .B2(new_n794), .ZN(new_n998));
  INV_X1    g0798(.A(new_n798), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n840), .A2(G294), .B1(G107), .B2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n996), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n801), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(G68), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n840), .A2(G159), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n780), .A2(new_n849), .B1(new_n423), .B2(new_n781), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(G50), .B2(new_n847), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n291), .B1(new_n788), .B2(new_n380), .C1(new_n202), .C2(new_n784), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(G137), .B2(new_n794), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1003), .A2(new_n1004), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1001), .A2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT47), .Z(new_n1011));
  OAI221_X1 g0811(.A(new_n992), .B1(new_n956), .B2(new_n815), .C1(new_n1011), .C2(new_n770), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n987), .A2(new_n1012), .ZN(G387));
  OR2_X1    g0813(.A1(new_n689), .A2(new_n815), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n757), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n1015), .A2(new_n698), .B1(G107), .B2(new_n223), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n242), .A2(new_n256), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n761), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n698), .ZN(new_n1019));
  AOI211_X1 g0819(.A(G45), .B(new_n1019), .C1(G68), .C2(G77), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n315), .A2(G50), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT50), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1018), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1016), .B1(new_n1017), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n755), .B1(new_n1024), .B2(new_n988), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1002), .A2(new_n990), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n774), .A2(new_n319), .B1(new_n847), .B2(G68), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n781), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n1028), .A2(G50), .B1(new_n779), .B2(G159), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n291), .B1(new_n788), .B2(new_n498), .C1(new_n380), .C2(new_n784), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G150), .B2(new_n794), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1026), .A2(new_n1027), .A3(new_n1029), .A4(new_n1031), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n798), .A2(new_n810), .B1(new_n571), .B2(new_n784), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n1028), .A2(G317), .B1(G303), .B2(new_n847), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n807), .B2(new_n780), .C1(new_n839), .C2(new_n804), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT48), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1033), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n1036), .B2(new_n1035), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT49), .Z(new_n1039));
  OAI221_X1 g0839(.A(new_n391), .B1(new_n758), .B2(new_n788), .C1(new_n842), .C2(new_n803), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1032), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1025), .B1(new_n1041), .B2(new_n767), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n982), .A2(new_n754), .B1(new_n1014), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n983), .A2(new_n696), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n982), .A2(new_n749), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(G393));
  AOI21_X1  g0846(.A(new_n697), .B1(new_n980), .B2(new_n984), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n984), .B2(new_n980), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n946), .A2(new_n766), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n842), .A2(new_n849), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n391), .B1(new_n836), .B2(G87), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n203), .B2(new_n784), .C1(new_n315), .C2(new_n777), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1050), .B(new_n1052), .C1(new_n840), .C2(G50), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1002), .A2(G77), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n780), .A2(new_n423), .B1(new_n329), .B2(new_n781), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT51), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1053), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n1028), .A2(G311), .B1(new_n779), .B2(G317), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT52), .Z(new_n1059));
  AOI21_X1  g0859(.A(new_n291), .B1(new_n836), .B2(G107), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(new_n810), .B2(new_n784), .C1(new_n571), .C2(new_n777), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(G322), .B2(new_n794), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n840), .A2(G303), .B1(G116), .B2(new_n999), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1059), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n770), .B1(new_n1057), .B2(new_n1064), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n246), .A2(new_n1018), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n988), .B1(G97), .B2(new_n695), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n756), .B(new_n1065), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n980), .A2(new_n754), .B1(new_n1049), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1048), .A2(new_n1069), .ZN(G390));
  NAND2_X1  g0870(.A1(new_n496), .A2(new_n728), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n935), .A2(new_n1071), .A3(new_n657), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n915), .B1(new_n727), .B2(new_n826), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n915), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1074), .A2(new_n726), .A3(G330), .A4(new_n828), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n829), .A2(new_n825), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n683), .B(new_n823), .C1(new_n734), .C2(new_n741), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1073), .A2(new_n825), .A3(new_n1075), .A4(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1072), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n916), .A2(new_n931), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n927), .A2(new_n928), .A3(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n904), .B1(new_n922), .B2(new_n926), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1079), .A2(new_n825), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n931), .B1(new_n1086), .B2(new_n1074), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  AND3_X1   g0888(.A1(new_n1084), .A2(new_n1075), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1075), .B1(new_n1084), .B2(new_n1088), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1082), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1084), .A2(new_n1088), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1075), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1084), .A2(new_n1088), .A3(new_n1075), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1094), .A2(new_n1081), .A3(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1091), .A2(new_n696), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n794), .A2(G125), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n391), .B1(new_n836), .B2(G50), .ZN(new_n1099));
  INV_X1    g0899(.A(G132), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1098), .B(new_n1099), .C1(new_n1100), .C2(new_n781), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n784), .A2(new_n423), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT53), .ZN(new_n1103));
  INV_X1    g0903(.A(G128), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(KEYINPUT54), .B(G143), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1103), .B1(new_n1104), .B2(new_n780), .C1(new_n777), .C2(new_n1105), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1101), .B(new_n1106), .C1(G137), .C2(new_n840), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1002), .A2(G159), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n794), .A2(G294), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1109), .A2(new_n391), .A3(new_n786), .A4(new_n854), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n779), .A2(G283), .B1(new_n847), .B2(G97), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n758), .B2(new_n781), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n1110), .B(new_n1112), .C1(G107), .C2(new_n840), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1107), .A2(new_n1108), .B1(new_n1054), .B2(new_n1113), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n755), .B1(new_n319), .B2(new_n834), .C1(new_n1114), .C2(new_n770), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n904), .A2(new_n920), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(new_n896), .B2(new_n898), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n901), .A2(new_n903), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n902), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n882), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n920), .B1(new_n1120), .B2(new_n904), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n765), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1115), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1124), .B1(new_n1125), .B2(new_n754), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1097), .A2(new_n1126), .ZN(G378));
  XOR2_X1   g0927(.A(new_n1072), .B(KEYINPUT122), .Z(new_n1128));
  NAND2_X1  g0928(.A1(new_n1096), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n726), .A2(new_n880), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n1120), .B2(new_n904), .ZN(new_n1131));
  OAI21_X1  g0931(.A(G330), .B1(new_n1131), .B2(KEYINPUT40), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n427), .A2(new_n884), .ZN(new_n1133));
  XOR2_X1   g0933(.A(new_n450), .B(new_n1133), .Z(new_n1134));
  XNOR2_X1  g0934(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1134), .B(new_n1135), .ZN(new_n1136));
  NOR3_X1   g0936(.A1(new_n1132), .A2(new_n905), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1136), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n873), .B1(new_n910), .B2(new_n906), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n881), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1085), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1138), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1122), .A2(new_n930), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n1137), .A2(new_n1142), .B1(new_n1143), .B2(new_n919), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1136), .B1(new_n1132), .B2(new_n905), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1139), .A2(new_n1141), .A3(new_n1138), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1145), .A2(new_n932), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1129), .A2(new_n1148), .A3(KEYINPUT57), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1096), .A2(new_n1128), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1149), .B(new_n696), .C1(KEYINPUT57), .C2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n755), .B1(G50), .B2(new_n834), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n515), .A2(new_n291), .ZN(new_n1153));
  AOI211_X1 g0953(.A(G50), .B(new_n1153), .C1(new_n310), .C2(new_n518), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n775), .A2(new_n498), .B1(new_n397), .B2(new_n781), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(G116), .B2(new_n779), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n990), .A2(new_n847), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1153), .B1(new_n202), .B2(new_n788), .C1(new_n380), .C2(new_n784), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(G283), .B2(new_n794), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1003), .A2(new_n1156), .A3(new_n1157), .A4(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT58), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1154), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(G125), .A2(new_n779), .B1(new_n774), .B2(G132), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n1104), .B2(new_n781), .ZN(new_n1164));
  INV_X1    g0964(.A(G137), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n777), .A2(new_n1165), .B1(new_n784), .B2(new_n1105), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n423), .B2(new_n801), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n794), .A2(G124), .ZN(new_n1170));
  AOI211_X1 g0970(.A(G33), .B(G41), .C1(new_n836), .C2(G159), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1162), .B1(new_n1161), .B2(new_n1160), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1152), .B1(new_n1174), .B2(new_n767), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n1138), .B2(new_n765), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT121), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n1148), .B2(new_n754), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1151), .A2(new_n1178), .ZN(G375));
  NAND2_X1  g0979(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n915), .A2(new_n764), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n839), .A2(new_n1105), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n780), .A2(new_n1100), .B1(new_n329), .B2(new_n784), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n781), .A2(new_n1165), .B1(new_n423), .B2(new_n777), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n291), .B1(new_n788), .B2(new_n202), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT123), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(G128), .B2(new_n794), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1185), .B(new_n1188), .C1(new_n201), .C2(new_n801), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n840), .A2(G116), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n780), .A2(new_n571), .B1(new_n397), .B2(new_n777), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(G283), .B2(new_n1028), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n391), .B1(new_n788), .B2(new_n380), .C1(new_n498), .C2(new_n784), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(G303), .B2(new_n794), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1026), .A2(new_n1190), .A3(new_n1192), .A4(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n770), .B1(new_n1189), .B2(new_n1195), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n756), .B(new_n1196), .C1(new_n203), .C2(new_n833), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1180), .A2(new_n754), .B1(new_n1181), .B2(new_n1197), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1081), .A2(new_n973), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n1072), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1198), .B1(new_n1199), .B2(new_n1202), .ZN(G381));
  OR2_X1    g1003(.A1(G393), .A2(G396), .ZN(new_n1204));
  OR4_X1    g1004(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1204), .ZN(new_n1205));
  OR4_X1    g1005(.A1(G387), .A2(new_n1205), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1006(.A(G378), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n681), .A2(G213), .ZN(new_n1208));
  XOR2_X1   g1008(.A(new_n1208), .B(KEYINPUT124), .Z(new_n1209));
  NAND2_X1  g1009(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  OAI211_X1 g1010(.A(G407), .B(G213), .C1(G375), .C2(new_n1210), .ZN(G409));
  INV_X1    g1011(.A(KEYINPUT126), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n987), .B2(new_n1012), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n987), .A2(new_n1212), .A3(new_n1012), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(G393), .A2(G396), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(G390), .A2(new_n1204), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1204), .A2(new_n1216), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1218), .A2(new_n1048), .A3(new_n1069), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1214), .A2(new_n1215), .A3(new_n1217), .A4(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1217), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1215), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1221), .B1(new_n1222), .B2(new_n1213), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1220), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT61), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1200), .A2(KEYINPUT60), .A3(new_n1072), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n696), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1082), .A2(KEYINPUT60), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1227), .B1(new_n1201), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1198), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n832), .B(new_n860), .C1(new_n1229), .C2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1202), .B1(KEYINPUT60), .B2(new_n1082), .ZN(new_n1232));
  OAI211_X1 g1032(.A(G384), .B(new_n1198), .C1(new_n1232), .C2(new_n1227), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1209), .A2(G2897), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1234), .B(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1148), .A2(new_n754), .ZN(new_n1237));
  AND2_X1   g1037(.A1(new_n1237), .A2(new_n1176), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n973), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1150), .A2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(G378), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1145), .A2(new_n932), .A3(new_n1146), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n932), .B1(new_n1146), .B2(new_n1145), .ZN(new_n1243));
  OAI21_X1  g1043(.A(KEYINPUT57), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1072), .B(KEYINPUT122), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(new_n1125), .B2(new_n1081), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n696), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT57), .B1(new_n1129), .B2(new_n1148), .ZN(new_n1248));
  OAI211_X1 g1048(.A(G378), .B(new_n1178), .C1(new_n1247), .C2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(KEYINPUT125), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT125), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1151), .A2(new_n1251), .A3(G378), .A4(new_n1178), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1241), .B1(new_n1250), .B2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1236), .B1(new_n1253), .B2(new_n1209), .ZN(new_n1254));
  NOR3_X1   g1054(.A1(new_n1253), .A2(new_n1209), .A3(new_n1234), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT62), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1225), .B(new_n1254), .C1(new_n1255), .C2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1250), .A2(new_n1252), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1241), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1209), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1234), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1260), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1263), .A2(KEYINPUT62), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1224), .B1(new_n1257), .B2(new_n1264), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1254), .A2(new_n1225), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT63), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1263), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1224), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1255), .A2(KEYINPUT63), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1266), .A2(new_n1268), .A3(new_n1269), .A4(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1265), .A2(new_n1271), .ZN(G405));
  AOI22_X1  g1072(.A1(new_n1262), .A2(KEYINPUT127), .B1(G375), .B2(new_n1207), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1258), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1262), .A2(KEYINPUT127), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1273), .B(new_n1258), .C1(KEYINPUT127), .C2(new_n1262), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(new_n1278), .B(new_n1269), .ZN(G402));
endmodule


