

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U552 ( .A(KEYINPUT17), .ZN(n518) );
  NOR2_X1 U553 ( .A1(n529), .A2(n528), .ZN(G164) );
  NAND2_X2 U554 ( .A1(n687), .A2(n757), .ZN(n739) );
  NOR2_X1 U555 ( .A1(G164), .A2(G1384), .ZN(n686) );
  NOR2_X1 U556 ( .A1(n693), .A2(n692), .ZN(n710) );
  XNOR2_X1 U557 ( .A(n716), .B(n715), .ZN(n734) );
  OR2_X1 U558 ( .A1(n755), .A2(KEYINPUT33), .ZN(n516) );
  NAND2_X1 U559 ( .A1(n908), .A2(n814), .ZN(n517) );
  NOR2_X1 U560 ( .A1(n739), .A2(n844), .ZN(n694) );
  NOR2_X1 U561 ( .A1(n698), .A2(n697), .ZN(n699) );
  INV_X1 U562 ( .A(KEYINPUT28), .ZN(n711) );
  INV_X1 U563 ( .A(KEYINPUT29), .ZN(n715) );
  NOR2_X1 U564 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U565 ( .A1(n748), .A2(n747), .ZN(n775) );
  NOR2_X1 U566 ( .A1(n771), .A2(n517), .ZN(n772) );
  NAND2_X1 U567 ( .A1(n881), .A2(G138), .ZN(n520) );
  NOR2_X1 U568 ( .A1(G651), .A2(n637), .ZN(n650) );
  NOR2_X2 U569 ( .A1(G2105), .A2(G2104), .ZN(n519) );
  XNOR2_X2 U570 ( .A(n519), .B(n518), .ZN(n881) );
  XOR2_X1 U571 ( .A(n520), .B(KEYINPUT85), .Z(n522) );
  INV_X1 U572 ( .A(G2105), .ZN(n524) );
  AND2_X1 U573 ( .A1(n524), .A2(G2104), .ZN(n880) );
  NAND2_X1 U574 ( .A1(n880), .A2(G102), .ZN(n521) );
  NAND2_X1 U575 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U576 ( .A(n523), .B(KEYINPUT86), .ZN(n529) );
  AND2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n884) );
  NAND2_X1 U578 ( .A1(G114), .A2(n884), .ZN(n526) );
  NOR2_X1 U579 ( .A1(G2104), .A2(n524), .ZN(n885) );
  NAND2_X1 U580 ( .A1(G126), .A2(n885), .ZN(n525) );
  NAND2_X1 U581 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U582 ( .A(KEYINPUT84), .B(n527), .ZN(n528) );
  XOR2_X1 U583 ( .A(G2446), .B(G2430), .Z(n531) );
  XNOR2_X1 U584 ( .A(G2451), .B(G2454), .ZN(n530) );
  XNOR2_X1 U585 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U586 ( .A(n532), .B(G2427), .Z(n534) );
  XNOR2_X1 U587 ( .A(G1341), .B(G1348), .ZN(n533) );
  XNOR2_X1 U588 ( .A(n534), .B(n533), .ZN(n538) );
  XOR2_X1 U589 ( .A(G2443), .B(KEYINPUT100), .Z(n536) );
  XNOR2_X1 U590 ( .A(G2438), .B(G2435), .ZN(n535) );
  XNOR2_X1 U591 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U592 ( .A(n538), .B(n537), .Z(n539) );
  AND2_X1 U593 ( .A1(G14), .A2(n539), .ZN(G401) );
  XNOR2_X1 U594 ( .A(G543), .B(KEYINPUT0), .ZN(n540) );
  XNOR2_X1 U595 ( .A(n540), .B(KEYINPUT65), .ZN(n637) );
  NAND2_X1 U596 ( .A1(G52), .A2(n650), .ZN(n541) );
  XOR2_X1 U597 ( .A(KEYINPUT66), .B(n541), .Z(n550) );
  NOR2_X1 U598 ( .A1(G651), .A2(G543), .ZN(n644) );
  NAND2_X1 U599 ( .A1(G90), .A2(n644), .ZN(n543) );
  INV_X1 U600 ( .A(G651), .ZN(n545) );
  NOR2_X1 U601 ( .A1(n637), .A2(n545), .ZN(n645) );
  NAND2_X1 U602 ( .A1(G77), .A2(n645), .ZN(n542) );
  NAND2_X1 U603 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U604 ( .A(n544), .B(KEYINPUT9), .ZN(n548) );
  NOR2_X1 U605 ( .A1(G543), .A2(n545), .ZN(n546) );
  XOR2_X1 U606 ( .A(KEYINPUT1), .B(n546), .Z(n643) );
  NAND2_X1 U607 ( .A1(G64), .A2(n643), .ZN(n547) );
  NAND2_X1 U608 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U609 ( .A1(n550), .A2(n549), .ZN(G171) );
  INV_X1 U610 ( .A(G171), .ZN(G301) );
  AND2_X1 U611 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U612 ( .A(G57), .ZN(G237) );
  INV_X1 U613 ( .A(G132), .ZN(G219) );
  NAND2_X1 U614 ( .A1(G65), .A2(n643), .ZN(n552) );
  NAND2_X1 U615 ( .A1(G53), .A2(n650), .ZN(n551) );
  NAND2_X1 U616 ( .A1(n552), .A2(n551), .ZN(n556) );
  NAND2_X1 U617 ( .A1(G91), .A2(n644), .ZN(n554) );
  NAND2_X1 U618 ( .A1(G78), .A2(n645), .ZN(n553) );
  NAND2_X1 U619 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U620 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U621 ( .A(n557), .B(KEYINPUT67), .Z(n709) );
  INV_X1 U622 ( .A(n709), .ZN(G299) );
  NAND2_X1 U623 ( .A1(n643), .A2(G63), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(KEYINPUT76), .ZN(n560) );
  NAND2_X1 U625 ( .A1(G51), .A2(n650), .ZN(n559) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(KEYINPUT6), .B(n561), .ZN(n568) );
  NAND2_X1 U628 ( .A1(n644), .A2(G89), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(KEYINPUT4), .ZN(n564) );
  NAND2_X1 U630 ( .A1(G76), .A2(n645), .ZN(n563) );
  NAND2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(KEYINPUT75), .B(n565), .ZN(n566) );
  XNOR2_X1 U633 ( .A(KEYINPUT5), .B(n566), .ZN(n567) );
  NOR2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U635 ( .A(KEYINPUT7), .B(n569), .Z(G168) );
  XOR2_X1 U636 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U637 ( .A1(G7), .A2(G661), .ZN(n570) );
  XOR2_X1 U638 ( .A(n570), .B(KEYINPUT10), .Z(n907) );
  NAND2_X1 U639 ( .A1(n907), .A2(G567), .ZN(n571) );
  XOR2_X1 U640 ( .A(KEYINPUT11), .B(n571), .Z(G234) );
  NAND2_X1 U641 ( .A1(n645), .A2(G68), .ZN(n572) );
  XNOR2_X1 U642 ( .A(KEYINPUT70), .B(n572), .ZN(n575) );
  NAND2_X1 U643 ( .A1(n644), .A2(G81), .ZN(n573) );
  XNOR2_X1 U644 ( .A(KEYINPUT12), .B(n573), .ZN(n574) );
  NAND2_X1 U645 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U646 ( .A(KEYINPUT13), .B(n576), .ZN(n580) );
  XOR2_X1 U647 ( .A(KEYINPUT14), .B(KEYINPUT69), .Z(n578) );
  NAND2_X1 U648 ( .A1(G56), .A2(n643), .ZN(n577) );
  XNOR2_X1 U649 ( .A(n578), .B(n577), .ZN(n579) );
  NAND2_X1 U650 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U651 ( .A(n581), .B(KEYINPUT71), .ZN(n583) );
  NAND2_X1 U652 ( .A1(G43), .A2(n650), .ZN(n582) );
  NAND2_X1 U653 ( .A1(n583), .A2(n582), .ZN(n698) );
  INV_X1 U654 ( .A(n698), .ZN(n925) );
  XNOR2_X1 U655 ( .A(G860), .B(KEYINPUT72), .ZN(n597) );
  NAND2_X1 U656 ( .A1(n925), .A2(n597), .ZN(G153) );
  NAND2_X1 U657 ( .A1(G79), .A2(n645), .ZN(n585) );
  NAND2_X1 U658 ( .A1(G54), .A2(n650), .ZN(n584) );
  NAND2_X1 U659 ( .A1(n585), .A2(n584), .ZN(n590) );
  NAND2_X1 U660 ( .A1(G92), .A2(n644), .ZN(n587) );
  NAND2_X1 U661 ( .A1(G66), .A2(n643), .ZN(n586) );
  NAND2_X1 U662 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U663 ( .A(KEYINPUT73), .B(n588), .Z(n589) );
  NOR2_X1 U664 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U665 ( .A(KEYINPUT15), .B(n591), .ZN(n915) );
  INV_X1 U666 ( .A(G868), .ZN(n662) );
  NAND2_X1 U667 ( .A1(n915), .A2(n662), .ZN(n592) );
  XNOR2_X1 U668 ( .A(n592), .B(KEYINPUT74), .ZN(n594) );
  NAND2_X1 U669 ( .A1(G868), .A2(G301), .ZN(n593) );
  NAND2_X1 U670 ( .A1(n594), .A2(n593), .ZN(G284) );
  NAND2_X1 U671 ( .A1(G286), .A2(G868), .ZN(n596) );
  NAND2_X1 U672 ( .A1(G299), .A2(n662), .ZN(n595) );
  NAND2_X1 U673 ( .A1(n596), .A2(n595), .ZN(G297) );
  INV_X1 U674 ( .A(G559), .ZN(n598) );
  NOR2_X1 U675 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U676 ( .A1(n915), .A2(n599), .ZN(n600) );
  XOR2_X1 U677 ( .A(KEYINPUT16), .B(n600), .Z(G148) );
  NOR2_X1 U678 ( .A1(G868), .A2(n698), .ZN(n601) );
  XOR2_X1 U679 ( .A(KEYINPUT77), .B(n601), .Z(n604) );
  INV_X1 U680 ( .A(n915), .ZN(n896) );
  NAND2_X1 U681 ( .A1(G868), .A2(n896), .ZN(n602) );
  NOR2_X1 U682 ( .A1(G559), .A2(n602), .ZN(n603) );
  NOR2_X1 U683 ( .A1(n604), .A2(n603), .ZN(G282) );
  NAND2_X1 U684 ( .A1(G123), .A2(n885), .ZN(n605) );
  XNOR2_X1 U685 ( .A(n605), .B(KEYINPUT18), .ZN(n607) );
  NAND2_X1 U686 ( .A1(n884), .A2(G111), .ZN(n606) );
  NAND2_X1 U687 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U688 ( .A1(G99), .A2(n880), .ZN(n609) );
  NAND2_X1 U689 ( .A1(G135), .A2(n881), .ZN(n608) );
  NAND2_X1 U690 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U691 ( .A1(n611), .A2(n610), .ZN(n996) );
  XNOR2_X1 U692 ( .A(n996), .B(G2096), .ZN(n612) );
  INV_X1 U693 ( .A(G2100), .ZN(n829) );
  NAND2_X1 U694 ( .A1(n612), .A2(n829), .ZN(G156) );
  NAND2_X1 U695 ( .A1(G559), .A2(n896), .ZN(n613) );
  XOR2_X1 U696 ( .A(n925), .B(n613), .Z(n660) );
  NOR2_X1 U697 ( .A1(n660), .A2(G860), .ZN(n620) );
  NAND2_X1 U698 ( .A1(G93), .A2(n644), .ZN(n615) );
  NAND2_X1 U699 ( .A1(G80), .A2(n645), .ZN(n614) );
  NAND2_X1 U700 ( .A1(n615), .A2(n614), .ZN(n619) );
  NAND2_X1 U701 ( .A1(G67), .A2(n643), .ZN(n617) );
  NAND2_X1 U702 ( .A1(G55), .A2(n650), .ZN(n616) );
  NAND2_X1 U703 ( .A1(n617), .A2(n616), .ZN(n618) );
  OR2_X1 U704 ( .A1(n619), .A2(n618), .ZN(n663) );
  XOR2_X1 U705 ( .A(n620), .B(n663), .Z(G145) );
  NAND2_X1 U706 ( .A1(G88), .A2(n644), .ZN(n622) );
  NAND2_X1 U707 ( .A1(G75), .A2(n645), .ZN(n621) );
  NAND2_X1 U708 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U709 ( .A1(G62), .A2(n643), .ZN(n624) );
  NAND2_X1 U710 ( .A1(G50), .A2(n650), .ZN(n623) );
  NAND2_X1 U711 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U712 ( .A1(n626), .A2(n625), .ZN(G166) );
  INV_X1 U713 ( .A(G166), .ZN(G303) );
  XOR2_X1 U714 ( .A(KEYINPUT2), .B(KEYINPUT79), .Z(n628) );
  NAND2_X1 U715 ( .A1(G73), .A2(n645), .ZN(n627) );
  XNOR2_X1 U716 ( .A(n628), .B(n627), .ZN(n635) );
  NAND2_X1 U717 ( .A1(G86), .A2(n644), .ZN(n630) );
  NAND2_X1 U718 ( .A1(G61), .A2(n643), .ZN(n629) );
  NAND2_X1 U719 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U720 ( .A1(n650), .A2(G48), .ZN(n631) );
  XOR2_X1 U721 ( .A(KEYINPUT80), .B(n631), .Z(n632) );
  NOR2_X1 U722 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U723 ( .A1(n635), .A2(n634), .ZN(G305) );
  NAND2_X1 U724 ( .A1(G49), .A2(n650), .ZN(n636) );
  XNOR2_X1 U725 ( .A(n636), .B(KEYINPUT78), .ZN(n642) );
  NAND2_X1 U726 ( .A1(G87), .A2(n637), .ZN(n639) );
  NAND2_X1 U727 ( .A1(G74), .A2(G651), .ZN(n638) );
  NAND2_X1 U728 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U729 ( .A1(n643), .A2(n640), .ZN(n641) );
  NAND2_X1 U730 ( .A1(n642), .A2(n641), .ZN(G288) );
  AND2_X1 U731 ( .A1(n643), .A2(G60), .ZN(n649) );
  NAND2_X1 U732 ( .A1(G85), .A2(n644), .ZN(n647) );
  NAND2_X1 U733 ( .A1(G72), .A2(n645), .ZN(n646) );
  NAND2_X1 U734 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U735 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U736 ( .A1(n650), .A2(G47), .ZN(n651) );
  NAND2_X1 U737 ( .A1(n652), .A2(n651), .ZN(G290) );
  XOR2_X1 U738 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n654) );
  XOR2_X1 U739 ( .A(G303), .B(KEYINPUT19), .Z(n653) );
  XNOR2_X1 U740 ( .A(n654), .B(n653), .ZN(n657) );
  XOR2_X1 U741 ( .A(G299), .B(G305), .Z(n655) );
  XNOR2_X1 U742 ( .A(n655), .B(G288), .ZN(n656) );
  XNOR2_X1 U743 ( .A(n657), .B(n656), .ZN(n659) );
  XOR2_X1 U744 ( .A(G290), .B(n663), .Z(n658) );
  XNOR2_X1 U745 ( .A(n659), .B(n658), .ZN(n895) );
  XNOR2_X1 U746 ( .A(n895), .B(n660), .ZN(n661) );
  NOR2_X1 U747 ( .A1(n662), .A2(n661), .ZN(n665) );
  NOR2_X1 U748 ( .A1(G868), .A2(n663), .ZN(n664) );
  NOR2_X1 U749 ( .A1(n665), .A2(n664), .ZN(G295) );
  NAND2_X1 U750 ( .A1(G2084), .A2(G2078), .ZN(n666) );
  XOR2_X1 U751 ( .A(KEYINPUT20), .B(n666), .Z(n667) );
  NAND2_X1 U752 ( .A1(G2090), .A2(n667), .ZN(n668) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n668), .ZN(n669) );
  NAND2_X1 U754 ( .A1(n669), .A2(G2072), .ZN(n670) );
  XOR2_X1 U755 ( .A(KEYINPUT83), .B(n670), .Z(G158) );
  XNOR2_X1 U756 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U757 ( .A(KEYINPUT68), .B(G82), .Z(G220) );
  NOR2_X1 U758 ( .A1(G220), .A2(G219), .ZN(n671) );
  XOR2_X1 U759 ( .A(KEYINPUT22), .B(n671), .Z(n672) );
  NOR2_X1 U760 ( .A1(G218), .A2(n672), .ZN(n673) );
  NAND2_X1 U761 ( .A1(G96), .A2(n673), .ZN(n826) );
  NAND2_X1 U762 ( .A1(n826), .A2(G2106), .ZN(n677) );
  NAND2_X1 U763 ( .A1(G120), .A2(G108), .ZN(n674) );
  NOR2_X1 U764 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U765 ( .A1(G69), .A2(n675), .ZN(n827) );
  NAND2_X1 U766 ( .A1(n827), .A2(G567), .ZN(n676) );
  NAND2_X1 U767 ( .A1(n677), .A2(n676), .ZN(n828) );
  NAND2_X1 U768 ( .A1(G661), .A2(G483), .ZN(n678) );
  NOR2_X1 U769 ( .A1(n828), .A2(n678), .ZN(n825) );
  NAND2_X1 U770 ( .A1(n825), .A2(G36), .ZN(G176) );
  NAND2_X1 U771 ( .A1(n881), .A2(G137), .ZN(n681) );
  NAND2_X1 U772 ( .A1(G101), .A2(n880), .ZN(n679) );
  XOR2_X1 U773 ( .A(KEYINPUT23), .B(n679), .Z(n680) );
  NAND2_X1 U774 ( .A1(n681), .A2(n680), .ZN(n685) );
  NAND2_X1 U775 ( .A1(G113), .A2(n884), .ZN(n683) );
  NAND2_X1 U776 ( .A1(G125), .A2(n885), .ZN(n682) );
  NAND2_X1 U777 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U778 ( .A1(n685), .A2(n684), .ZN(G160) );
  NAND2_X1 U779 ( .A1(G160), .A2(G40), .ZN(n758) );
  INV_X1 U780 ( .A(n758), .ZN(n687) );
  XNOR2_X1 U781 ( .A(n686), .B(KEYINPUT64), .ZN(n757) );
  INV_X1 U782 ( .A(KEYINPUT94), .ZN(n688) );
  XNOR2_X2 U783 ( .A(n739), .B(n688), .ZN(n700) );
  XNOR2_X1 U784 ( .A(G2078), .B(KEYINPUT25), .ZN(n970) );
  NAND2_X1 U785 ( .A1(n700), .A2(n970), .ZN(n690) );
  INV_X1 U786 ( .A(G1961), .ZN(n840) );
  NAND2_X1 U787 ( .A1(n840), .A2(n739), .ZN(n689) );
  NAND2_X1 U788 ( .A1(n690), .A2(n689), .ZN(n720) );
  NAND2_X1 U789 ( .A1(n720), .A2(G171), .ZN(n732) );
  NAND2_X1 U790 ( .A1(n700), .A2(G2072), .ZN(n691) );
  XNOR2_X1 U791 ( .A(n691), .B(KEYINPUT27), .ZN(n693) );
  INV_X1 U792 ( .A(G1956), .ZN(n843) );
  NOR2_X1 U793 ( .A1(n700), .A2(n843), .ZN(n692) );
  NAND2_X1 U794 ( .A1(n709), .A2(n710), .ZN(n708) );
  INV_X1 U795 ( .A(G1996), .ZN(n844) );
  XOR2_X1 U796 ( .A(n694), .B(KEYINPUT26), .Z(n696) );
  NAND2_X1 U797 ( .A1(n739), .A2(G1341), .ZN(n695) );
  NAND2_X1 U798 ( .A1(n696), .A2(n695), .ZN(n697) );
  OR2_X1 U799 ( .A1(n896), .A2(n699), .ZN(n706) );
  NAND2_X1 U800 ( .A1(n896), .A2(n699), .ZN(n704) );
  NAND2_X1 U801 ( .A1(G2067), .A2(n700), .ZN(n702) );
  NAND2_X1 U802 ( .A1(G1348), .A2(n739), .ZN(n701) );
  NAND2_X1 U803 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U804 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U805 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U806 ( .A1(n708), .A2(n707), .ZN(n714) );
  NOR2_X1 U807 ( .A1(n710), .A2(n709), .ZN(n712) );
  XNOR2_X1 U808 ( .A(n712), .B(n711), .ZN(n713) );
  NAND2_X1 U809 ( .A1(n714), .A2(n713), .ZN(n716) );
  NAND2_X1 U810 ( .A1(n732), .A2(n734), .ZN(n725) );
  NOR2_X1 U811 ( .A1(G2084), .A2(n739), .ZN(n729) );
  NAND2_X1 U812 ( .A1(G8), .A2(n739), .ZN(n781) );
  NOR2_X1 U813 ( .A1(G1966), .A2(n781), .ZN(n726) );
  NOR2_X1 U814 ( .A1(n729), .A2(n726), .ZN(n717) );
  NAND2_X1 U815 ( .A1(G8), .A2(n717), .ZN(n718) );
  XNOR2_X1 U816 ( .A(KEYINPUT30), .B(n718), .ZN(n719) );
  NOR2_X1 U817 ( .A1(G168), .A2(n719), .ZN(n722) );
  NOR2_X1 U818 ( .A1(G171), .A2(n720), .ZN(n721) );
  NOR2_X1 U819 ( .A1(n722), .A2(n721), .ZN(n724) );
  XNOR2_X1 U820 ( .A(KEYINPUT31), .B(KEYINPUT95), .ZN(n723) );
  XNOR2_X1 U821 ( .A(n724), .B(n723), .ZN(n735) );
  AND2_X1 U822 ( .A1(n725), .A2(n735), .ZN(n727) );
  XNOR2_X1 U823 ( .A(n728), .B(KEYINPUT96), .ZN(n731) );
  NAND2_X1 U824 ( .A1(n729), .A2(G8), .ZN(n730) );
  NAND2_X1 U825 ( .A1(n731), .A2(n730), .ZN(n748) );
  AND2_X1 U826 ( .A1(n732), .A2(G286), .ZN(n733) );
  NAND2_X1 U827 ( .A1(n734), .A2(n733), .ZN(n738) );
  INV_X1 U828 ( .A(G286), .ZN(n736) );
  OR2_X1 U829 ( .A1(n736), .A2(n735), .ZN(n737) );
  AND2_X1 U830 ( .A1(n738), .A2(n737), .ZN(n744) );
  NOR2_X1 U831 ( .A1(G1971), .A2(n781), .ZN(n741) );
  NOR2_X1 U832 ( .A1(G2090), .A2(n739), .ZN(n740) );
  NOR2_X1 U833 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U834 ( .A1(n742), .A2(G303), .ZN(n743) );
  NAND2_X1 U835 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U836 ( .A1(n745), .A2(G8), .ZN(n746) );
  XNOR2_X1 U837 ( .A(n746), .B(KEYINPUT32), .ZN(n747) );
  NOR2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n918) );
  NOR2_X1 U839 ( .A1(G1971), .A2(G303), .ZN(n749) );
  NOR2_X1 U840 ( .A1(n918), .A2(n749), .ZN(n750) );
  NAND2_X1 U841 ( .A1(n775), .A2(n750), .ZN(n751) );
  XNOR2_X1 U842 ( .A(KEYINPUT97), .B(n751), .ZN(n754) );
  NAND2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n920) );
  INV_X1 U844 ( .A(n920), .ZN(n752) );
  OR2_X1 U845 ( .A1(n781), .A2(n752), .ZN(n753) );
  NOR2_X1 U846 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U847 ( .A1(n918), .A2(KEYINPUT33), .ZN(n756) );
  NOR2_X1 U848 ( .A1(n756), .A2(n781), .ZN(n771) );
  XOR2_X1 U849 ( .A(G1981), .B(G305), .Z(n908) );
  NOR2_X1 U850 ( .A1(n758), .A2(n757), .ZN(n818) );
  NAND2_X1 U851 ( .A1(G104), .A2(n880), .ZN(n760) );
  NAND2_X1 U852 ( .A1(G140), .A2(n881), .ZN(n759) );
  NAND2_X1 U853 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U854 ( .A(KEYINPUT34), .B(n761), .ZN(n768) );
  XNOR2_X1 U855 ( .A(KEYINPUT35), .B(KEYINPUT88), .ZN(n766) );
  NAND2_X1 U856 ( .A1(n884), .A2(G116), .ZN(n764) );
  NAND2_X1 U857 ( .A1(n885), .A2(G128), .ZN(n762) );
  XOR2_X1 U858 ( .A(KEYINPUT87), .B(n762), .Z(n763) );
  NAND2_X1 U859 ( .A1(n764), .A2(n763), .ZN(n765) );
  XOR2_X1 U860 ( .A(n766), .B(n765), .Z(n767) );
  NOR2_X1 U861 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U862 ( .A(n769), .B(KEYINPUT36), .Z(n770) );
  XNOR2_X1 U863 ( .A(KEYINPUT89), .B(n770), .ZN(n862) );
  XNOR2_X1 U864 ( .A(KEYINPUT37), .B(G2067), .ZN(n816) );
  NOR2_X1 U865 ( .A1(n862), .A2(n816), .ZN(n994) );
  NAND2_X1 U866 ( .A1(n818), .A2(n994), .ZN(n814) );
  NAND2_X1 U867 ( .A1(n516), .A2(n772), .ZN(n786) );
  NOR2_X1 U868 ( .A1(G2090), .A2(G303), .ZN(n773) );
  NAND2_X1 U869 ( .A1(G8), .A2(n773), .ZN(n774) );
  NAND2_X1 U870 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U871 ( .A(n776), .B(KEYINPUT98), .ZN(n777) );
  NAND2_X1 U872 ( .A1(n777), .A2(n781), .ZN(n783) );
  NOR2_X1 U873 ( .A1(G1981), .A2(G305), .ZN(n778) );
  XNOR2_X1 U874 ( .A(n778), .B(KEYINPUT93), .ZN(n779) );
  XNOR2_X1 U875 ( .A(KEYINPUT24), .B(n779), .ZN(n780) );
  OR2_X1 U876 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U877 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U878 ( .A1(n814), .A2(n784), .ZN(n785) );
  NAND2_X1 U879 ( .A1(n786), .A2(n785), .ZN(n808) );
  NAND2_X1 U880 ( .A1(n880), .A2(G105), .ZN(n787) );
  XNOR2_X1 U881 ( .A(n787), .B(KEYINPUT38), .ZN(n789) );
  NAND2_X1 U882 ( .A1(G117), .A2(n884), .ZN(n788) );
  NAND2_X1 U883 ( .A1(n789), .A2(n788), .ZN(n792) );
  NAND2_X1 U884 ( .A1(G129), .A2(n885), .ZN(n790) );
  XNOR2_X1 U885 ( .A(KEYINPUT91), .B(n790), .ZN(n791) );
  NOR2_X1 U886 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U887 ( .A(n793), .B(KEYINPUT92), .ZN(n795) );
  NAND2_X1 U888 ( .A1(G141), .A2(n881), .ZN(n794) );
  NAND2_X1 U889 ( .A1(n795), .A2(n794), .ZN(n874) );
  NAND2_X1 U890 ( .A1(n874), .A2(G1996), .ZN(n804) );
  NAND2_X1 U891 ( .A1(G131), .A2(n881), .ZN(n797) );
  NAND2_X1 U892 ( .A1(G119), .A2(n885), .ZN(n796) );
  NAND2_X1 U893 ( .A1(n797), .A2(n796), .ZN(n801) );
  NAND2_X1 U894 ( .A1(G95), .A2(n880), .ZN(n799) );
  NAND2_X1 U895 ( .A1(G107), .A2(n884), .ZN(n798) );
  NAND2_X1 U896 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U897 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U898 ( .A(KEYINPUT90), .B(n802), .Z(n860) );
  NAND2_X1 U899 ( .A1(n860), .A2(G1991), .ZN(n803) );
  NAND2_X1 U900 ( .A1(n804), .A2(n803), .ZN(n993) );
  INV_X1 U901 ( .A(n993), .ZN(n805) );
  XOR2_X1 U902 ( .A(G1986), .B(G290), .Z(n912) );
  NAND2_X1 U903 ( .A1(n805), .A2(n912), .ZN(n806) );
  NAND2_X1 U904 ( .A1(n806), .A2(n818), .ZN(n807) );
  NAND2_X1 U905 ( .A1(n808), .A2(n807), .ZN(n821) );
  NOR2_X1 U906 ( .A1(G1996), .A2(n874), .ZN(n1008) );
  NOR2_X1 U907 ( .A1(G1991), .A2(n860), .ZN(n1000) );
  NOR2_X1 U908 ( .A1(G1986), .A2(G290), .ZN(n809) );
  NOR2_X1 U909 ( .A1(n1000), .A2(n809), .ZN(n810) );
  XOR2_X1 U910 ( .A(KEYINPUT99), .B(n810), .Z(n811) );
  NOR2_X1 U911 ( .A1(n993), .A2(n811), .ZN(n812) );
  NOR2_X1 U912 ( .A1(n1008), .A2(n812), .ZN(n813) );
  XNOR2_X1 U913 ( .A(n813), .B(KEYINPUT39), .ZN(n815) );
  NAND2_X1 U914 ( .A1(n815), .A2(n814), .ZN(n817) );
  NAND2_X1 U915 ( .A1(n862), .A2(n816), .ZN(n997) );
  NAND2_X1 U916 ( .A1(n817), .A2(n997), .ZN(n819) );
  NAND2_X1 U917 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U918 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U919 ( .A(n822), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n907), .ZN(G217) );
  AND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n823) );
  NAND2_X1 U922 ( .A1(G661), .A2(n823), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U924 ( .A1(n825), .A2(n824), .ZN(G188) );
  XOR2_X1 U925 ( .A(G108), .B(KEYINPUT108), .Z(G238) );
  INV_X1 U927 ( .A(G120), .ZN(G236) );
  INV_X1 U928 ( .A(G96), .ZN(G221) );
  NOR2_X1 U929 ( .A1(n827), .A2(n826), .ZN(G325) );
  INV_X1 U930 ( .A(G325), .ZN(G261) );
  INV_X1 U931 ( .A(n828), .ZN(G319) );
  XNOR2_X1 U932 ( .A(n829), .B(KEYINPUT43), .ZN(n831) );
  XNOR2_X1 U933 ( .A(KEYINPUT42), .B(G2678), .ZN(n830) );
  XNOR2_X1 U934 ( .A(n831), .B(n830), .ZN(n835) );
  XOR2_X1 U935 ( .A(KEYINPUT101), .B(G2090), .Z(n833) );
  XNOR2_X1 U936 ( .A(G2067), .B(G2072), .ZN(n832) );
  XNOR2_X1 U937 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U938 ( .A(n835), .B(n834), .Z(n837) );
  XNOR2_X1 U939 ( .A(KEYINPUT102), .B(G2096), .ZN(n836) );
  XNOR2_X1 U940 ( .A(n837), .B(n836), .ZN(n839) );
  XOR2_X1 U941 ( .A(G2084), .B(G2078), .Z(n838) );
  XNOR2_X1 U942 ( .A(n839), .B(n838), .ZN(G227) );
  XNOR2_X1 U943 ( .A(G1971), .B(n840), .ZN(n842) );
  XNOR2_X1 U944 ( .A(G1986), .B(G1966), .ZN(n841) );
  XNOR2_X1 U945 ( .A(n842), .B(n841), .ZN(n848) );
  XNOR2_X1 U946 ( .A(G1976), .B(n843), .ZN(n846) );
  XOR2_X1 U947 ( .A(n844), .B(G1991), .Z(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U949 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U950 ( .A(KEYINPUT103), .B(G2474), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(n852) );
  XOR2_X1 U952 ( .A(G1981), .B(KEYINPUT41), .Z(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(G229) );
  NAND2_X1 U954 ( .A1(G124), .A2(n885), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n853), .B(KEYINPUT44), .ZN(n855) );
  NAND2_X1 U956 ( .A1(n884), .A2(G112), .ZN(n854) );
  NAND2_X1 U957 ( .A1(n855), .A2(n854), .ZN(n859) );
  NAND2_X1 U958 ( .A1(G100), .A2(n880), .ZN(n857) );
  NAND2_X1 U959 ( .A1(G136), .A2(n881), .ZN(n856) );
  NAND2_X1 U960 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U961 ( .A1(n859), .A2(n858), .ZN(G162) );
  XOR2_X1 U962 ( .A(G160), .B(n860), .Z(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U964 ( .A(KEYINPUT106), .B(KEYINPUT48), .Z(n864) );
  XNOR2_X1 U965 ( .A(KEYINPUT46), .B(KEYINPUT104), .ZN(n863) );
  XNOR2_X1 U966 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U967 ( .A(n866), .B(n865), .Z(n878) );
  NAND2_X1 U968 ( .A1(G118), .A2(n884), .ZN(n868) );
  NAND2_X1 U969 ( .A1(G130), .A2(n885), .ZN(n867) );
  NAND2_X1 U970 ( .A1(n868), .A2(n867), .ZN(n873) );
  NAND2_X1 U971 ( .A1(G106), .A2(n880), .ZN(n870) );
  NAND2_X1 U972 ( .A1(G142), .A2(n881), .ZN(n869) );
  NAND2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U974 ( .A(n871), .B(KEYINPUT45), .Z(n872) );
  NOR2_X1 U975 ( .A1(n873), .A2(n872), .ZN(n875) );
  XNOR2_X1 U976 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U977 ( .A(G164), .B(n876), .ZN(n877) );
  XNOR2_X1 U978 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U979 ( .A(n879), .B(n996), .Z(n893) );
  NAND2_X1 U980 ( .A1(G103), .A2(n880), .ZN(n883) );
  NAND2_X1 U981 ( .A1(G139), .A2(n881), .ZN(n882) );
  NAND2_X1 U982 ( .A1(n883), .A2(n882), .ZN(n890) );
  NAND2_X1 U983 ( .A1(G115), .A2(n884), .ZN(n887) );
  NAND2_X1 U984 ( .A1(G127), .A2(n885), .ZN(n886) );
  NAND2_X1 U985 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U986 ( .A(KEYINPUT47), .B(n888), .Z(n889) );
  NOR2_X1 U987 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U988 ( .A(KEYINPUT105), .B(n891), .Z(n1003) );
  XNOR2_X1 U989 ( .A(n1003), .B(G162), .ZN(n892) );
  XNOR2_X1 U990 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U991 ( .A1(G37), .A2(n894), .ZN(G395) );
  XOR2_X1 U992 ( .A(n895), .B(G286), .Z(n898) );
  XOR2_X1 U993 ( .A(G301), .B(n896), .Z(n897) );
  XNOR2_X1 U994 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U995 ( .A(n899), .B(n925), .Z(n900) );
  NOR2_X1 U996 ( .A1(G37), .A2(n900), .ZN(G397) );
  NOR2_X1 U997 ( .A1(G227), .A2(G229), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n901), .B(KEYINPUT49), .ZN(n902) );
  NOR2_X1 U999 ( .A1(G401), .A2(n902), .ZN(n903) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n903), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(KEYINPUT107), .B(n904), .ZN(n906) );
  NOR2_X1 U1002 ( .A1(G395), .A2(G397), .ZN(n905) );
  NAND2_X1 U1003 ( .A1(n906), .A2(n905), .ZN(G225) );
  INV_X1 U1004 ( .A(G225), .ZN(G308) );
  INV_X1 U1005 ( .A(G69), .ZN(G235) );
  INV_X1 U1006 ( .A(n907), .ZN(G223) );
  XNOR2_X1 U1007 ( .A(G1966), .B(G168), .ZN(n909) );
  NAND2_X1 U1008 ( .A1(n909), .A2(n908), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(n910), .B(KEYINPUT115), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(KEYINPUT57), .B(n911), .ZN(n934) );
  XOR2_X1 U1011 ( .A(G299), .B(G1956), .Z(n913) );
  NAND2_X1 U1012 ( .A1(n913), .A2(n912), .ZN(n931) );
  XNOR2_X1 U1013 ( .A(G1971), .B(KEYINPUT118), .ZN(n914) );
  XOR2_X1 U1014 ( .A(n914), .B(G166), .Z(n917) );
  XNOR2_X1 U1015 ( .A(G1348), .B(n915), .ZN(n916) );
  NOR2_X1 U1016 ( .A1(n917), .A2(n916), .ZN(n929) );
  INV_X1 U1017 ( .A(n918), .ZN(n919) );
  NAND2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1019 ( .A(n921), .B(KEYINPUT117), .ZN(n924) );
  XOR2_X1 U1020 ( .A(G301), .B(G1961), .Z(n922) );
  XNOR2_X1 U1021 ( .A(n922), .B(KEYINPUT116), .ZN(n923) );
  NAND2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n927) );
  XOR2_X1 U1023 ( .A(G1341), .B(n925), .Z(n926) );
  NOR2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1027 ( .A(KEYINPUT119), .B(n932), .ZN(n933) );
  NOR2_X1 U1028 ( .A1(n934), .A2(n933), .ZN(n936) );
  XOR2_X1 U1029 ( .A(KEYINPUT56), .B(G16), .Z(n935) );
  NOR2_X1 U1030 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1031 ( .A(KEYINPUT120), .B(n937), .Z(n991) );
  XOR2_X1 U1032 ( .A(G1961), .B(G5), .Z(n961) );
  XOR2_X1 U1033 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n944) );
  XNOR2_X1 U1034 ( .A(G1971), .B(G22), .ZN(n939) );
  XNOR2_X1 U1035 ( .A(G23), .B(G1976), .ZN(n938) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n942) );
  XOR2_X1 U1037 ( .A(G1986), .B(KEYINPUT124), .Z(n940) );
  XNOR2_X1 U1038 ( .A(G24), .B(n940), .ZN(n941) );
  NAND2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1040 ( .A(n944), .B(n943), .ZN(n959) );
  XNOR2_X1 U1041 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n954) );
  XOR2_X1 U1042 ( .A(G20), .B(G1956), .Z(n948) );
  XNOR2_X1 U1043 ( .A(G1341), .B(G19), .ZN(n946) );
  XNOR2_X1 U1044 ( .A(G1981), .B(G6), .ZN(n945) );
  NOR2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1047 ( .A(KEYINPUT121), .B(n949), .ZN(n952) );
  XNOR2_X1 U1048 ( .A(G1348), .B(KEYINPUT59), .ZN(n950) );
  XNOR2_X1 U1049 ( .A(n950), .B(G4), .ZN(n951) );
  NAND2_X1 U1050 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1051 ( .A(n954), .B(n953), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(G21), .B(G1966), .ZN(n955) );
  NOR2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1054 ( .A(n957), .B(KEYINPUT123), .ZN(n958) );
  NOR2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(n962), .B(KEYINPUT61), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(n963), .B(KEYINPUT126), .ZN(n964) );
  NOR2_X1 U1059 ( .A1(G16), .A2(n964), .ZN(n989) );
  XNOR2_X1 U1060 ( .A(G29), .B(KEYINPUT113), .ZN(n985) );
  XNOR2_X1 U1061 ( .A(KEYINPUT55), .B(KEYINPUT109), .ZN(n1015) );
  XNOR2_X1 U1062 ( .A(KEYINPUT54), .B(G34), .ZN(n965) );
  XNOR2_X1 U1063 ( .A(n965), .B(KEYINPUT111), .ZN(n966) );
  XNOR2_X1 U1064 ( .A(G2084), .B(n966), .ZN(n981) );
  XNOR2_X1 U1065 ( .A(G2090), .B(G35), .ZN(n979) );
  XOR2_X1 U1066 ( .A(G1991), .B(G25), .Z(n967) );
  NAND2_X1 U1067 ( .A1(n967), .A2(G28), .ZN(n976) );
  XNOR2_X1 U1068 ( .A(G2067), .B(G26), .ZN(n969) );
  XNOR2_X1 U1069 ( .A(G33), .B(G2072), .ZN(n968) );
  NOR2_X1 U1070 ( .A1(n969), .A2(n968), .ZN(n974) );
  XOR2_X1 U1071 ( .A(n970), .B(G27), .Z(n972) );
  XNOR2_X1 U1072 ( .A(G1996), .B(G32), .ZN(n971) );
  NOR2_X1 U1073 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1074 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1075 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1076 ( .A(KEYINPUT53), .B(n977), .ZN(n978) );
  NOR2_X1 U1077 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1078 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1079 ( .A(n982), .B(KEYINPUT112), .ZN(n983) );
  XNOR2_X1 U1080 ( .A(n1015), .B(n983), .ZN(n984) );
  NAND2_X1 U1081 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1082 ( .A(KEYINPUT114), .B(n986), .ZN(n987) );
  NAND2_X1 U1083 ( .A1(n987), .A2(G11), .ZN(n988) );
  NOR2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1086 ( .A(n992), .B(KEYINPUT127), .ZN(n1020) );
  NOR2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n1002) );
  XOR2_X1 U1088 ( .A(G2084), .B(G160), .Z(n995) );
  NOR2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n998) );
  NAND2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1013) );
  XOR2_X1 U1093 ( .A(G2072), .B(n1003), .Z(n1005) );
  XOR2_X1 U1094 ( .A(G164), .B(G2078), .Z(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1096 ( .A(KEYINPUT50), .B(n1006), .ZN(n1011) );
  XOR2_X1 U1097 ( .A(G2090), .B(G162), .Z(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1099 ( .A(KEYINPUT51), .B(n1009), .Z(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(n1014), .B(KEYINPUT52), .ZN(n1016) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(KEYINPUT110), .B(n1017), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(G29), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1021), .ZN(G150) );
  INV_X1 U1108 ( .A(G150), .ZN(G311) );
endmodule

