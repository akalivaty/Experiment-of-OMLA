//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 0 0 1 1 0 0 1 1 0 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n547, new_n549, new_n550, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n562,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n592, new_n593, new_n596, new_n598,
    new_n599, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n462), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n462), .A2(new_n464), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n465), .A2(new_n471), .ZN(G160));
  NAND2_X1  g047(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n477), .A2(KEYINPUT66), .A3(G136), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n479));
  INV_X1    g054(.A(G136), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n479), .B1(new_n469), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n476), .A2(new_n464), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n485));
  AND4_X1   g060(.A1(new_n478), .A2(new_n481), .A3(new_n483), .A4(new_n485), .ZN(G162));
  NAND4_X1  g061(.A1(new_n473), .A2(new_n475), .A3(G138), .A4(new_n464), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n462), .A2(new_n489), .A3(G138), .A4(new_n464), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G114), .C2(new_n464), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n473), .A2(new_n475), .A3(G126), .A4(G2105), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT67), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT67), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n491), .A2(new_n498), .A3(new_n495), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n508), .A2(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  NAND3_X1  g091(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n517));
  XOR2_X1   g092(.A(new_n517), .B(KEYINPUT68), .Z(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  INV_X1    g095(.A(G51), .ZN(new_n521));
  INV_X1    g096(.A(G89), .ZN(new_n522));
  OAI221_X1 g097(.A(new_n520), .B1(new_n512), .B2(new_n521), .C1(new_n510), .C2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n518), .A2(new_n523), .ZN(G168));
  AOI22_X1  g099(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n507), .ZN(new_n526));
  INV_X1    g101(.A(G90), .ZN(new_n527));
  INV_X1    g102(.A(G52), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n510), .A2(new_n527), .B1(new_n512), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n526), .A2(new_n529), .ZN(G171));
  XOR2_X1   g105(.A(KEYINPUT71), .B(G81), .Z(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G43), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n510), .A2(new_n532), .B1(new_n512), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(G68), .A2(G543), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n502), .A2(new_n504), .ZN(new_n536));
  INV_X1    g111(.A(G56), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT69), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g115(.A(G651), .B1(new_n538), .B2(new_n539), .ZN(new_n541));
  OR3_X1    g116(.A1(new_n540), .A2(new_n541), .A3(KEYINPUT70), .ZN(new_n542));
  OAI21_X1  g117(.A(KEYINPUT70), .B1(new_n540), .B2(new_n541), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n534), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT72), .ZN(G153));
  AND3_X1   g121(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G36), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n547), .A2(new_n550), .ZN(G188));
  NAND3_X1  g126(.A1(new_n509), .A2(G53), .A3(G543), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT9), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n505), .A2(new_n509), .ZN(new_n554));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n536), .B2(new_n556), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n554), .A2(G91), .B1(new_n557), .B2(G651), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n553), .A2(new_n558), .ZN(G299));
  INV_X1    g134(.A(G171), .ZN(G301));
  INV_X1    g135(.A(G168), .ZN(G286));
  NAND2_X1  g136(.A1(new_n554), .A2(G87), .ZN(new_n562));
  INV_X1    g137(.A(new_n512), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G49), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n562), .A2(new_n564), .A3(new_n565), .ZN(G288));
  NAND2_X1  g141(.A1(new_n554), .A2(G86), .ZN(new_n567));
  NAND2_X1  g142(.A1(G73), .A2(G543), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT73), .ZN(new_n569));
  AND3_X1   g144(.A1(new_n502), .A2(new_n504), .A3(G61), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n563), .A2(G48), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n567), .A2(new_n571), .A3(new_n572), .ZN(G305));
  AOI22_X1  g148(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n574), .A2(new_n507), .ZN(new_n575));
  XOR2_X1   g150(.A(KEYINPUT74), .B(G85), .Z(new_n576));
  INV_X1    g151(.A(G47), .ZN(new_n577));
  OAI22_X1  g152(.A1(new_n510), .A2(new_n576), .B1(new_n512), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT75), .ZN(G290));
  NAND2_X1  g155(.A1(G301), .A2(G868), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n505), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G54), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n582), .A2(new_n507), .B1(new_n583), .B2(new_n512), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT76), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n554), .A2(G92), .ZN(new_n586));
  XOR2_X1   g161(.A(new_n586), .B(KEYINPUT10), .Z(new_n587));
  NAND2_X1  g162(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n581), .B1(new_n589), .B2(G868), .ZN(G284));
  OAI21_X1  g165(.A(new_n581), .B1(new_n589), .B2(G868), .ZN(G321));
  NAND2_X1  g166(.A1(G286), .A2(G868), .ZN(new_n592));
  INV_X1    g167(.A(G299), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(G868), .B2(new_n593), .ZN(G297));
  XOR2_X1   g169(.A(G297), .B(KEYINPUT77), .Z(G280));
  INV_X1    g170(.A(G559), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n589), .B1(new_n596), .B2(G860), .ZN(G148));
  NAND2_X1  g172(.A1(new_n589), .A2(new_n596), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G868), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(G868), .B2(new_n544), .ZN(G323));
  XNOR2_X1  g175(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g176(.A1(new_n477), .A2(G135), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT78), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n482), .A2(G123), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n464), .A2(G111), .ZN(new_n605));
  OAI21_X1  g180(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n606));
  OAI211_X1 g181(.A(new_n603), .B(new_n604), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(G2096), .Z(new_n610));
  NAND2_X1  g185(.A1(new_n462), .A2(new_n467), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(G2100), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n610), .A2(new_n614), .ZN(G156));
  INV_X1    g190(.A(G14), .ZN(new_n616));
  XNOR2_X1  g191(.A(G2427), .B(G2430), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT82), .ZN(new_n618));
  XOR2_X1   g193(.A(KEYINPUT81), .B(G2438), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(KEYINPUT15), .B(G2435), .Z(new_n621));
  OR2_X1    g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n622), .A2(KEYINPUT14), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2443), .B(G2446), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2451), .B(G2454), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n624), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n628), .A2(new_n630), .ZN(new_n632));
  AND2_X1   g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G1341), .B(G1348), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n616), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n631), .A2(new_n632), .ZN(new_n636));
  INV_X1    g211(.A(new_n634), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT83), .Z(G401));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2067), .B(G2678), .Z(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n642), .A2(new_n643), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(new_n646), .A3(KEYINPUT17), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2096), .B(G2100), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT86), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n649), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT84), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n644), .B2(new_n648), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n652), .B(new_n655), .ZN(G227));
  XNOR2_X1  g231(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1956), .B(G2474), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT87), .ZN(new_n660));
  XOR2_X1   g235(.A(G1961), .B(G1966), .Z(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n664), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n660), .A2(new_n661), .ZN(new_n667));
  AOI22_X1  g242(.A1(new_n665), .A2(KEYINPUT20), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n666), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(new_n662), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n668), .B(new_n670), .C1(KEYINPUT20), .C2(new_n665), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(G1991), .Z(new_n672));
  INV_X1    g247(.A(G1996), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n672), .B(G1996), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n678), .A2(new_n675), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n658), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n675), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n674), .A2(new_n676), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n681), .A2(new_n682), .A3(new_n657), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(G229));
  AND2_X1   g259(.A1(KEYINPUT89), .A2(G16), .ZN(new_n685));
  NOR2_X1   g260(.A1(KEYINPUT89), .A2(G16), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G22), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G166), .B2(new_n688), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(G1971), .Z(new_n691));
  MUX2_X1   g266(.A(G6), .B(G305), .S(G16), .Z(new_n692));
  XOR2_X1   g267(.A(KEYINPUT32), .B(G1981), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(G16), .A2(G23), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT90), .ZN(new_n696));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(G288), .B2(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT33), .B(G1976), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT91), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n698), .B(new_n700), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n691), .A2(new_n694), .A3(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT92), .B(KEYINPUT34), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  MUX2_X1   g279(.A(G24), .B(G290), .S(new_n687), .Z(new_n705));
  INV_X1    g280(.A(G1986), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G25), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n477), .A2(G131), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n482), .A2(G119), .ZN(new_n711));
  OR3_X1    g286(.A1(KEYINPUT88), .A2(G95), .A3(G2105), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n464), .A2(G107), .ZN(new_n713));
  OAI21_X1  g288(.A(KEYINPUT88), .B1(G95), .B2(G2105), .ZN(new_n714));
  NAND4_X1  g289(.A1(new_n712), .A2(new_n713), .A3(G2104), .A4(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n710), .A2(new_n711), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n709), .B1(new_n717), .B2(new_n708), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT35), .B(G1991), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n704), .A2(new_n707), .A3(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT36), .Z(new_n722));
  NAND2_X1  g297(.A1(new_n482), .A2(G129), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT96), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n467), .A2(G105), .ZN(new_n725));
  NAND3_X1  g300(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT26), .ZN(new_n727));
  AOI211_X1 g302(.A(new_n725), .B(new_n727), .C1(G141), .C2(new_n477), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G29), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT97), .ZN(new_n732));
  INV_X1    g307(.A(G32), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n732), .B1(new_n708), .B2(new_n733), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT27), .B(G1996), .Z(new_n735));
  NOR2_X1   g310(.A1(new_n589), .A2(new_n697), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G4), .B2(new_n697), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n734), .A2(new_n735), .B1(G1348), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(G168), .A2(G16), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G16), .B2(G21), .ZN(new_n741));
  INV_X1    g316(.A(G1966), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT100), .Z(new_n744));
  NAND2_X1  g319(.A1(G162), .A2(G29), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G29), .B2(G35), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT101), .B(KEYINPUT29), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(G2090), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n744), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n708), .A2(G27), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G164), .B2(new_n708), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n752), .A2(G2078), .ZN(new_n753));
  INV_X1    g328(.A(G1348), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n737), .A2(new_n754), .B1(G2078), .B2(new_n752), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n739), .A2(new_n750), .A3(new_n753), .A4(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT31), .B(G11), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT99), .B(KEYINPUT30), .Z(new_n758));
  NOR2_X1   g333(.A1(new_n758), .A2(G28), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(G28), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(new_n708), .ZN(new_n761));
  OAI221_X1 g336(.A(new_n757), .B1(new_n759), .B2(new_n761), .C1(new_n609), .C2(new_n708), .ZN(new_n762));
  NOR2_X1   g337(.A1(G5), .A2(G16), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G171), .B2(G16), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(G1961), .Z(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n742), .B2(new_n741), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(G34), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n768), .A2(KEYINPUT24), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n768), .A2(KEYINPUT24), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n708), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G160), .B2(new_n708), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT95), .Z(new_n773));
  INV_X1    g348(.A(G2084), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n708), .A2(G26), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n482), .A2(G128), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n477), .A2(G140), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n464), .A2(G116), .ZN(new_n778));
  OAI21_X1  g353(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n776), .B(new_n777), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n775), .B1(new_n780), .B2(G29), .ZN(new_n781));
  MUX2_X1   g356(.A(new_n775), .B(new_n781), .S(KEYINPUT28), .Z(new_n782));
  INV_X1    g357(.A(G2067), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n773), .A2(new_n774), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  INV_X1    g360(.A(new_n773), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(G2084), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n708), .A2(G33), .ZN(new_n788));
  AOI21_X1  g363(.A(KEYINPUT25), .B1(new_n467), .B2(G103), .ZN(new_n789));
  AND3_X1   g364(.A1(new_n467), .A2(KEYINPUT25), .A3(G103), .ZN(new_n790));
  INV_X1    g365(.A(G139), .ZN(new_n791));
  OAI22_X1  g366(.A1(new_n789), .A2(new_n790), .B1(new_n469), .B2(new_n791), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n793), .A2(new_n464), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n794), .A2(KEYINPUT93), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(KEYINPUT93), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n792), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n788), .B1(new_n797), .B2(new_n708), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT94), .B(G2072), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n767), .A2(new_n784), .A3(new_n787), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n688), .A2(G19), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n544), .B2(new_n688), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1341), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n756), .A2(new_n801), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n688), .A2(G20), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT23), .Z(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G299), .B2(G16), .ZN(new_n808));
  INV_X1    g383(.A(G1956), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n748), .B2(G2090), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n811), .A2(KEYINPUT102), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n734), .A2(new_n735), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT98), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n811), .A2(KEYINPUT102), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n805), .A2(new_n812), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n722), .A2(new_n816), .ZN(G311));
  INV_X1    g392(.A(G311), .ZN(G150));
  NAND2_X1  g393(.A1(new_n505), .A2(G67), .ZN(new_n819));
  NAND2_X1  g394(.A1(G80), .A2(G543), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n507), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(KEYINPUT104), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(KEYINPUT104), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n554), .A2(G93), .B1(new_n563), .B2(G55), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT105), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(G860), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT37), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n588), .A2(new_n596), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT106), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT39), .ZN(new_n833));
  INV_X1    g408(.A(new_n544), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n827), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n544), .A2(new_n825), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n837), .B(new_n838), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n833), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(new_n828), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n833), .A2(new_n839), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n830), .B1(new_n841), .B2(new_n842), .ZN(G145));
  NAND2_X1  g418(.A1(new_n477), .A2(G142), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n464), .A2(G118), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(G130), .B2(new_n482), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(new_n612), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n716), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT108), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT107), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n797), .A2(new_n852), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n797), .A2(new_n852), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(new_n853), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n780), .B(new_n496), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n730), .B(new_n856), .ZN(new_n857));
  MUX2_X1   g432(.A(new_n853), .B(new_n855), .S(new_n857), .Z(new_n858));
  OR2_X1    g433(.A1(new_n851), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n850), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n609), .B(G160), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(G162), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n862), .A2(KEYINPUT110), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(KEYINPUT110), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n859), .B(new_n860), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n851), .B(new_n858), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(new_n862), .ZN(new_n867));
  XOR2_X1   g442(.A(KEYINPUT109), .B(G37), .Z(new_n868));
  NAND3_X1  g443(.A1(new_n865), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g445(.A(new_n837), .B(new_n598), .Z(new_n871));
  NAND2_X1  g446(.A1(new_n589), .A2(G299), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n588), .A2(new_n593), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n588), .B(G299), .ZN(new_n876));
  XOR2_X1   g451(.A(KEYINPUT111), .B(KEYINPUT41), .Z(new_n877));
  AND2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n876), .A2(KEYINPUT41), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n875), .B1(new_n871), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(KEYINPUT42), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT42), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n875), .B(new_n883), .C1(new_n871), .C2(new_n880), .ZN(new_n884));
  XNOR2_X1  g459(.A(G290), .B(G288), .ZN(new_n885));
  XOR2_X1   g460(.A(G303), .B(G305), .Z(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n882), .A2(new_n884), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n888), .B1(new_n882), .B2(new_n884), .ZN(new_n890));
  OAI21_X1  g465(.A(G868), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n827), .A2(G868), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(G295));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n892), .ZN(G331));
  INV_X1    g469(.A(KEYINPUT43), .ZN(new_n895));
  XNOR2_X1  g470(.A(G171), .B(KEYINPUT112), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(G286), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n837), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n897), .A2(new_n835), .A3(new_n836), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n874), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n899), .B(new_n900), .C1(new_n878), .C2(new_n879), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n902), .A2(new_n888), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n868), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n874), .A2(KEYINPUT41), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n874), .A2(new_n877), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n906), .A2(new_n899), .A3(new_n900), .A4(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n888), .B1(new_n902), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT113), .B1(new_n905), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n909), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT113), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n911), .A2(new_n912), .A3(new_n868), .A4(new_n904), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n895), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(G37), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n904), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n888), .B1(new_n902), .B2(new_n903), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT44), .B1(new_n914), .B2(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n911), .A2(new_n895), .A3(new_n868), .A4(new_n904), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n921), .B1(new_n918), .B2(new_n895), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n920), .A2(new_n924), .ZN(G397));
  AOI22_X1  g500(.A1(new_n477), .A2(G137), .B1(G101), .B2(new_n467), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n926), .B(G40), .C1(new_n464), .C2(new_n463), .ZN(new_n927));
  AOI21_X1  g502(.A(G1384), .B1(new_n491), .B2(new_n495), .ZN(new_n928));
  NOR3_X1   g503(.A1(new_n927), .A2(new_n928), .A3(KEYINPUT45), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n780), .B(new_n783), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n930), .B1(new_n730), .B2(new_n931), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n929), .A2(KEYINPUT46), .A3(new_n673), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT46), .B1(new_n929), .B2(new_n673), .ZN(new_n934));
  NOR3_X1   g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n935), .B(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n730), .A2(G1996), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n729), .A2(new_n673), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n931), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n717), .A2(new_n719), .ZN(new_n941));
  OAI22_X1  g516(.A1(new_n940), .A2(new_n941), .B1(G2067), .B2(new_n780), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n929), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT48), .ZN(new_n944));
  NOR2_X1   g519(.A1(G290), .A2(G1986), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n944), .B1(new_n946), .B2(new_n930), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n945), .A2(KEYINPUT48), .A3(new_n929), .ZN(new_n948));
  XOR2_X1   g523(.A(new_n716), .B(new_n719), .Z(new_n949));
  NOR2_X1   g524(.A1(new_n940), .A2(new_n949), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n947), .B(new_n948), .C1(new_n950), .C2(new_n930), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n937), .A2(new_n943), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G1384), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n497), .A2(new_n953), .A3(new_n499), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT50), .ZN(new_n955));
  XNOR2_X1  g530(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n928), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n927), .B1(new_n958), .B2(KEYINPUT115), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT115), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n928), .A2(new_n960), .A3(new_n957), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n955), .A2(new_n959), .A3(new_n774), .A4(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n928), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT45), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n927), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n953), .A4(new_n499), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n742), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n962), .A2(new_n968), .A3(G168), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT51), .ZN(new_n970));
  AND2_X1   g545(.A1(KEYINPUT123), .A2(G8), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n962), .A2(new_n968), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n973), .A2(G8), .A3(G286), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n970), .B1(new_n969), .B2(new_n971), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT62), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n976), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT62), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n978), .A2(new_n979), .A3(new_n974), .A4(new_n972), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n953), .ZN(new_n981));
  INV_X1    g556(.A(G40), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n465), .A2(new_n471), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n984), .B1(new_n964), .B2(new_n954), .ZN(new_n985));
  INV_X1    g560(.A(G2078), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT53), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n955), .A2(new_n961), .A3(new_n959), .ZN(new_n988));
  XNOR2_X1  g563(.A(KEYINPUT124), .B(G1961), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n987), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n965), .A2(KEYINPUT53), .A3(new_n986), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n966), .ZN(new_n993));
  AOI21_X1  g568(.A(G301), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n977), .A2(new_n980), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G8), .ZN(new_n996));
  AOI211_X1 g571(.A(new_n996), .B(G286), .C1(new_n962), .C2(new_n968), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT63), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n927), .B1(new_n963), .B2(new_n956), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT50), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n497), .A2(new_n1001), .A3(new_n953), .A4(new_n499), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n809), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n927), .B1(KEYINPUT45), .B2(new_n928), .ZN(new_n1005));
  XNOR2_X1  g580(.A(KEYINPUT56), .B(G2072), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n497), .A2(new_n953), .A3(new_n499), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1005), .B(new_n1006), .C1(new_n1007), .C2(KEYINPUT45), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1004), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n553), .A2(new_n558), .A3(KEYINPUT57), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT121), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n553), .A2(new_n558), .A3(KEYINPUT121), .A4(KEYINPUT57), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n557), .A2(G651), .ZN(new_n1015));
  INV_X1    g590(.A(G91), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1015), .B1(new_n1016), .B2(new_n510), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT120), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT120), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n558), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1018), .A2(new_n1020), .A3(new_n553), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT57), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1014), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1009), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1004), .A2(new_n1024), .A3(new_n1008), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n589), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n983), .A2(new_n928), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(G2067), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1030), .B1(new_n988), .B2(new_n754), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1026), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT59), .ZN(new_n1033));
  XOR2_X1   g608(.A(KEYINPUT58), .B(G1341), .Z(new_n1034));
  NAND2_X1  g609(.A1(new_n1029), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1036), .B1(new_n985), .B2(new_n673), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n544), .A2(KEYINPUT122), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1033), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n673), .B(new_n1005), .C1(new_n1007), .C2(KEYINPUT45), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n1035), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1038), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(KEYINPUT59), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1039), .A2(new_n1043), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1004), .A2(new_n1024), .A3(new_n1008), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1024), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT61), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT61), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1026), .A2(new_n1048), .A3(new_n1027), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1044), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1031), .A2(KEYINPUT60), .A3(new_n588), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n588), .B1(new_n1031), .B2(KEYINPUT60), .ZN(new_n1052));
  OAI22_X1  g627(.A1(new_n1051), .A2(new_n1052), .B1(KEYINPUT60), .B2(new_n1031), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1032), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  XOR2_X1   g629(.A(G171), .B(KEYINPUT54), .Z(new_n1055));
  AND3_X1   g630(.A1(new_n990), .A2(new_n993), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n992), .A2(new_n981), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1055), .B1(new_n990), .B2(new_n1057), .ZN(new_n1058));
  OAI22_X1  g633(.A1(new_n1056), .A2(new_n1058), .B1(new_n976), .B2(new_n975), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n995), .B(new_n999), .C1(new_n1054), .C2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1029), .A2(G8), .ZN(new_n1061));
  INV_X1    g636(.A(new_n571), .ZN(new_n1062));
  INV_X1    g637(.A(G86), .ZN(new_n1063));
  INV_X1    g638(.A(G48), .ZN(new_n1064));
  OAI22_X1  g639(.A1(new_n510), .A2(new_n1063), .B1(new_n512), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(G1981), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G1981), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n567), .A2(new_n1067), .A3(new_n571), .A4(new_n572), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1061), .B1(new_n1070), .B2(KEYINPUT49), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(new_n1070), .B2(KEYINPUT49), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT49), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1069), .A2(KEYINPUT116), .A3(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1071), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1071), .A2(new_n1073), .A3(KEYINPUT117), .A4(new_n1075), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n1081));
  INV_X1    g656(.A(G288), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1081), .B1(new_n1082), .B2(G1976), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1061), .B1(G1976), .B2(new_n1082), .ZN(new_n1084));
  MUX2_X1   g659(.A(new_n1081), .B(new_n1083), .S(new_n1084), .Z(new_n1085));
  AND2_X1   g660(.A1(new_n1080), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n1087));
  NAND2_X1  g662(.A1(G303), .A2(G8), .ZN(new_n1088));
  XOR2_X1   g663(.A(new_n1088), .B(KEYINPUT55), .Z(new_n1089));
  OR2_X1    g664(.A1(new_n985), .A2(G1971), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(G2090), .B2(new_n1003), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1089), .B1(new_n1091), .B2(G8), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1086), .B1(new_n1087), .B2(new_n1092), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1092), .A2(new_n1087), .ZN(new_n1094));
  OR2_X1    g669(.A1(new_n988), .A2(G2090), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n996), .B1(new_n1095), .B2(new_n1090), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1096), .A2(new_n1089), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1093), .A2(new_n1094), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1060), .A2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(G288), .A2(G1976), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1080), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1101), .A2(KEYINPUT118), .A3(new_n1068), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1061), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT118), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1100), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1105), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1068), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1104), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1102), .A2(new_n1103), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1080), .A2(new_n1085), .A3(new_n997), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1096), .A2(new_n1089), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT63), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1086), .A2(new_n1097), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1109), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1099), .A2(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g691(.A(G290), .B(new_n706), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n930), .B1(new_n950), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT125), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1114), .B1(new_n1060), .B2(new_n1098), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT125), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1121), .A2(new_n1122), .A3(new_n1118), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n952), .B1(new_n1120), .B2(new_n1123), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g699(.A1(G227), .A2(new_n460), .ZN(new_n1126));
  INV_X1    g700(.A(new_n1126), .ZN(new_n1127));
  AOI21_X1  g701(.A(new_n1127), .B1(new_n635), .B2(new_n638), .ZN(new_n1128));
  NAND3_X1  g702(.A1(new_n1128), .A2(new_n683), .A3(new_n680), .ZN(new_n1129));
  NAND2_X1  g703(.A1(new_n1129), .A2(KEYINPUT127), .ZN(new_n1130));
  INV_X1    g704(.A(KEYINPUT127), .ZN(new_n1131));
  NAND4_X1  g705(.A1(new_n1128), .A2(new_n680), .A3(new_n1131), .A4(new_n683), .ZN(new_n1132));
  NAND4_X1  g706(.A1(new_n1130), .A2(new_n869), .A3(new_n922), .A4(new_n1132), .ZN(G225));
  INV_X1    g707(.A(G225), .ZN(G308));
endmodule


