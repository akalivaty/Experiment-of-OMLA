//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 1 0 1 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 1 0 1 1 0 0 0 1 1 0 0 0 1 0 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n861, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n991, new_n992;
  AOI21_X1  g000(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT69), .ZN(new_n203));
  OR2_X1    g002(.A1(G197gat), .A2(G204gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205));
  AND3_X1   g004(.A1(new_n204), .A2(KEYINPUT68), .A3(new_n205), .ZN(new_n206));
  AOI21_X1  g005(.A(KEYINPUT68), .B1(new_n204), .B2(new_n205), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n203), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G211gat), .B(G218gat), .Z(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n209), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n203), .B(new_n211), .C1(new_n206), .C2(new_n207), .ZN(new_n212));
  AND2_X1   g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT24), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(G183gat), .A3(G190gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n218), .A2(KEYINPUT23), .ZN(new_n219));
  OR2_X1    g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(KEYINPUT24), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n218), .A2(KEYINPUT23), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n217), .A2(new_n219), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT25), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n225), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT27), .B(G183gat), .ZN(new_n228));
  INV_X1    g027(.A(G190gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT28), .ZN(new_n232));
  AOI22_X1  g031(.A1(new_n231), .A2(new_n232), .B1(G183gat), .B2(G190gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n234), .B(KEYINPUT26), .ZN(new_n235));
  AOI22_X1  g034(.A1(new_n216), .A2(new_n235), .B1(new_n230), .B2(KEYINPUT28), .ZN(new_n236));
  AOI22_X1  g035(.A1(new_n226), .A2(new_n227), .B1(new_n233), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G226gat), .A2(G233gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(KEYINPUT70), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n239), .A2(KEYINPUT29), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n237), .A2(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n213), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n210), .A2(new_n212), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n241), .B(new_n246), .C1(new_n237), .C2(new_n243), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G64gat), .B(G92gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT71), .ZN(new_n250));
  XNOR2_X1  g049(.A(G8gat), .B(G36gat), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n250), .B(new_n251), .Z(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n248), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n245), .A2(new_n252), .A3(new_n247), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n254), .A2(new_n255), .A3(KEYINPUT30), .ZN(new_n256));
  OR3_X1    g055(.A1(new_n248), .A2(KEYINPUT30), .A3(new_n253), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(G225gat), .A2(G233gat), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G155gat), .A2(G162gat), .ZN(new_n261));
  OR2_X1    g060(.A1(new_n261), .A2(KEYINPUT72), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(KEYINPUT72), .ZN(new_n263));
  INV_X1    g062(.A(G155gat), .ZN(new_n264));
  INV_X1    g063(.A(G162gat), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n262), .A2(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(G148gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G141gat), .ZN(new_n268));
  INV_X1    g067(.A(G141gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(G148gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT73), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n268), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(KEYINPUT72), .A2(KEYINPUT2), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G141gat), .B(G148gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n275), .A2(new_n271), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n266), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(KEYINPUT74), .B(G162gat), .Z(new_n278));
  OAI21_X1  g077(.A(KEYINPUT2), .B1(new_n278), .B2(new_n264), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n265), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n275), .B1(new_n280), .B2(new_n261), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT66), .ZN(new_n283));
  INV_X1    g082(.A(G120gat), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n283), .B1(new_n284), .B2(G113gat), .ZN(new_n285));
  INV_X1    g084(.A(G113gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n286), .A2(KEYINPUT66), .A3(G120gat), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n285), .B(new_n287), .C1(new_n286), .C2(G120gat), .ZN(new_n288));
  INV_X1    g087(.A(G134gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G127gat), .ZN(new_n290));
  INV_X1    g089(.A(G127gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(G134gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT1), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n290), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n286), .A2(G120gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n284), .A2(G113gat), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n293), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT65), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(new_n291), .B2(G134gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n289), .A2(KEYINPUT65), .A3(G127gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(new_n300), .A3(new_n292), .ZN(new_n301));
  AOI22_X1  g100(.A1(new_n288), .A2(new_n294), .B1(new_n297), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n277), .A2(new_n282), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n260), .B1(new_n304), .B2(KEYINPUT4), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n277), .A2(new_n282), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT3), .ZN(new_n307));
  INV_X1    g106(.A(new_n302), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT3), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n277), .A2(new_n282), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n307), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT75), .B(KEYINPUT4), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n303), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n305), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT5), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n306), .A2(new_n308), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(new_n303), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n315), .B1(new_n317), .B2(new_n260), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n260), .A2(KEYINPUT5), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n303), .A2(KEYINPUT4), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n268), .A2(new_n270), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT73), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n323), .A2(new_n273), .A3(new_n272), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n324), .A2(new_n266), .B1(new_n279), .B2(new_n281), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n302), .B1(new_n325), .B2(new_n309), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n321), .B1(new_n326), .B2(new_n307), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n304), .A2(new_n312), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n320), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G1gat), .B(G29gat), .ZN(new_n331));
  INV_X1    g130(.A(G85gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT0), .B(G57gat), .ZN(new_n334));
  XOR2_X1   g133(.A(new_n333), .B(new_n334), .Z(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n330), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT6), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT76), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT77), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT76), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n337), .A2(new_n342), .A3(new_n338), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n319), .A2(new_n330), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n335), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n340), .A2(new_n341), .A3(new_n343), .A4(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(KEYINPUT6), .A3(new_n335), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n339), .A2(KEYINPUT76), .B1(new_n344), .B2(new_n335), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n341), .B1(new_n349), .B2(new_n343), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n258), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n226), .A2(new_n227), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n233), .A2(new_n236), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n308), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(G227gat), .ZN(new_n355));
  INV_X1    g154(.A(G233gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n237), .A2(new_n302), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n354), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT34), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n354), .A2(new_n359), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(new_n357), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT32), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT33), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  XOR2_X1   g166(.A(G15gat), .B(G43gat), .Z(new_n368));
  XNOR2_X1  g167(.A(G71gat), .B(G99gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n368), .B(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n365), .A2(new_n367), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT67), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n366), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n373), .B1(new_n372), .B2(new_n370), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n364), .A2(KEYINPUT32), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n362), .A2(new_n371), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n358), .B1(new_n354), .B2(new_n359), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT32), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n370), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n377), .A2(KEYINPUT33), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n375), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n361), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  XOR2_X1   g182(.A(KEYINPUT31), .B(G50gat), .Z(new_n384));
  XNOR2_X1  g183(.A(new_n384), .B(KEYINPUT78), .ZN(new_n385));
  XNOR2_X1  g184(.A(G78gat), .B(G106gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(KEYINPUT79), .ZN(new_n388));
  XNOR2_X1  g187(.A(KEYINPUT83), .B(G22gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(G228gat), .A2(G233gat), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT29), .B1(new_n210), .B2(new_n212), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n306), .B1(new_n391), .B2(KEYINPUT3), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT81), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n390), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n310), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n213), .B(KEYINPUT82), .C1(new_n395), .C2(KEYINPUT29), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT82), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT29), .B1(new_n325), .B2(new_n309), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n397), .B1(new_n398), .B2(new_n246), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  OAI211_X1 g199(.A(KEYINPUT81), .B(new_n306), .C1(new_n391), .C2(KEYINPUT3), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n394), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT80), .B1(new_n398), .B2(new_n246), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n392), .ZN(new_n404));
  NOR3_X1   g203(.A1(new_n398), .A2(KEYINPUT80), .A3(new_n246), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n390), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n389), .B1(new_n402), .B2(new_n406), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n402), .A2(new_n406), .A3(new_n389), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT84), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n402), .A2(new_n406), .A3(new_n389), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT84), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n388), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  AND2_X1   g212(.A1(new_n411), .A2(new_n387), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n402), .A2(new_n406), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(G22gat), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n383), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT35), .B1(new_n351), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT87), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g220(.A(KEYINPUT87), .B(KEYINPUT35), .C1(new_n351), .C2(new_n418), .ZN(new_n422));
  INV_X1    g221(.A(new_n258), .ZN(new_n423));
  XOR2_X1   g222(.A(KEYINPUT86), .B(KEYINPUT35), .Z(new_n424));
  NOR2_X1   g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n345), .A2(new_n338), .A3(new_n337), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n347), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n428), .A2(new_n418), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n421), .A2(new_n422), .A3(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n402), .A2(new_n406), .A3(new_n409), .A4(new_n389), .ZN(new_n432));
  INV_X1    g231(.A(new_n415), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n412), .B(new_n432), .C1(new_n389), .C2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n388), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n414), .A2(new_n416), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n256), .A2(new_n257), .A3(new_n345), .ZN(new_n439));
  INV_X1    g238(.A(new_n321), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n311), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n441), .A2(new_n328), .A3(new_n260), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT85), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT85), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n441), .A2(new_n444), .A3(new_n328), .A4(new_n260), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT39), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n316), .A2(new_n303), .A3(new_n259), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n443), .A2(KEYINPUT39), .A3(new_n445), .A4(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n336), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT40), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n448), .A2(KEYINPUT40), .A3(new_n336), .A4(new_n450), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n439), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n255), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n248), .A2(KEYINPUT37), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT37), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n245), .A2(new_n458), .A3(new_n247), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n457), .A2(new_n459), .A3(new_n253), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n456), .B1(new_n460), .B2(KEYINPUT38), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT38), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n457), .A2(new_n459), .A3(new_n462), .A4(new_n253), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n461), .A2(new_n347), .A3(new_n426), .A4(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n438), .A2(new_n455), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n376), .A2(new_n382), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT36), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n466), .B(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n349), .A2(new_n343), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT77), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n471), .A2(new_n347), .A3(new_n346), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n438), .B1(new_n472), .B2(new_n258), .ZN(new_n473));
  OR2_X1    g272(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n431), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n476), .A2(KEYINPUT89), .ZN(new_n477));
  INV_X1    g276(.A(G29gat), .ZN(new_n478));
  INV_X1    g277(.A(G36gat), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT14), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n482), .A2(new_n478), .A3(new_n479), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n483), .A2(KEYINPUT89), .A3(new_n476), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(G50gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(G43gat), .ZN(new_n487));
  INV_X1    g286(.A(G43gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(G50gat), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n487), .A2(new_n489), .A3(KEYINPUT15), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT15), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n488), .A2(G50gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n486), .A2(G43gat), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n496), .A2(KEYINPUT90), .A3(new_n490), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT90), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n498), .B(new_n493), .C1(new_n494), .C2(new_n495), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT92), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n483), .A2(new_n476), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT91), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n483), .A2(KEYINPUT91), .A3(new_n476), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n480), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n500), .A2(new_n501), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n501), .B1(new_n500), .B2(new_n506), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n492), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT17), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OR2_X1    g310(.A1(G15gat), .A2(G22gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(G15gat), .A2(G22gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(G1gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT16), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n512), .A2(new_n515), .A3(new_n513), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(G8gat), .B1(new_n518), .B2(KEYINPUT93), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n517), .B(new_n518), .C1(KEYINPUT93), .C2(G8gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g322(.A(KEYINPUT17), .B(new_n492), .C1(new_n507), .C2(new_n508), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n511), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(G229gat), .A2(G233gat), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n521), .A2(KEYINPUT94), .A3(new_n522), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT94), .B1(new_n521), .B2(new_n522), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(new_n509), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n525), .A2(KEYINPUT18), .A3(new_n526), .A4(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n526), .B(KEYINPUT13), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n530), .A2(new_n509), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n500), .A2(new_n506), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT92), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n500), .A2(new_n501), .A3(new_n506), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n491), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n539), .A2(new_n529), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n534), .B1(new_n535), .B2(new_n540), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n532), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n525), .A2(new_n526), .A3(new_n531), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT18), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT95), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n547));
  XNOR2_X1  g346(.A(G113gat), .B(G141gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G169gat), .B(G197gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(KEYINPUT12), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n542), .B(new_n545), .C1(new_n546), .C2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n532), .A2(new_n546), .A3(new_n541), .ZN(new_n554));
  INV_X1    g353(.A(new_n552), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n532), .A2(new_n541), .ZN(new_n556));
  AOI22_X1  g355(.A1(new_n509), .A2(new_n510), .B1(new_n522), .B2(new_n521), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n540), .B1(new_n557), .B2(new_n524), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT18), .B1(new_n558), .B2(new_n526), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n554), .B(new_n555), .C1(new_n556), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n553), .A2(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(G183gat), .B(G211gat), .Z(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n562), .B(new_n563), .Z(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(G57gat), .B(G64gat), .Z(new_n566));
  INV_X1    g365(.A(G71gat), .ZN(new_n567));
  INV_X1    g366(.A(G78gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G71gat), .A2(G78gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT9), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n566), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G57gat), .B(G64gat), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n570), .B(new_n569), .C1(new_n575), .C2(new_n572), .ZN(new_n576));
  AND2_X1   g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT21), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n529), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT96), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT96), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n529), .A2(new_n581), .A3(new_n578), .ZN(new_n582));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n580), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n584), .B1(new_n580), .B2(new_n582), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n577), .A2(KEYINPUT21), .ZN(new_n588));
  XOR2_X1   g387(.A(G127gat), .B(G155gat), .Z(new_n589));
  XOR2_X1   g388(.A(new_n588), .B(new_n589), .Z(new_n590));
  NOR3_X1   g389(.A1(new_n586), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n590), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n580), .A2(new_n582), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(new_n583), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n592), .B1(new_n594), .B2(new_n585), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n565), .B1(new_n591), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n590), .B1(new_n586), .B2(new_n587), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n594), .A2(new_n585), .A3(new_n592), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n597), .A2(new_n598), .A3(new_n564), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G190gat), .B(G218gat), .Z(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT98), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G134gat), .B(G162gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G85gat), .A2(G92gat), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT7), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G99gat), .A2(G106gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(KEYINPUT8), .ZN(new_n615));
  INV_X1    g414(.A(G92gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n332), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n614), .ZN(new_n619));
  NOR2_X1   g418(.A1(G99gat), .A2(G106gat), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT97), .ZN(new_n621));
  NOR3_X1   g420(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(G99gat), .ZN(new_n623));
  INV_X1    g422(.A(G106gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(KEYINPUT97), .B1(new_n625), .B2(new_n614), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n613), .B(new_n618), .C1(new_n622), .C2(new_n626), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n615), .A2(new_n611), .A3(new_n617), .A4(new_n612), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n621), .B1(new_n619), .B2(new_n620), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n625), .A2(KEYINPUT97), .A3(new_n614), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n511), .A2(new_n524), .A3(new_n632), .ZN(new_n633));
  AND3_X1   g432(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n634));
  INV_X1    g433(.A(new_n632), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n634), .B1(new_n509), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n602), .A2(new_n603), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n608), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n637), .A2(new_n639), .A3(new_n608), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(KEYINPUT99), .B1(new_n600), .B2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n642), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n645), .A2(new_n640), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT99), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n596), .A2(new_n646), .A3(new_n647), .A4(new_n599), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n635), .A2(KEYINPUT10), .A3(new_n577), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT100), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n622), .A2(new_n626), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n651), .B1(new_n652), .B2(new_n628), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n632), .A2(new_n653), .A3(new_n577), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n574), .A2(new_n576), .ZN(new_n655));
  OAI211_X1 g454(.A(new_n627), .B(new_n631), .C1(new_n655), .C2(new_n651), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT10), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT101), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n660));
  AOI211_X1 g459(.A(new_n660), .B(KEYINPUT10), .C1(new_n654), .C2(new_n656), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n650), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(G230gat), .A2(G233gat), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n663), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n654), .A2(new_n665), .A3(new_n656), .ZN(new_n666));
  XNOR2_X1  g465(.A(G120gat), .B(G148gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(G176gat), .B(G204gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n664), .A2(new_n666), .A3(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n670), .B1(new_n664), .B2(new_n666), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n649), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n475), .A2(new_n561), .A3(new_n676), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n677), .A2(KEYINPUT102), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(KEYINPUT102), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n472), .A2(KEYINPUT103), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n472), .A2(KEYINPUT103), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g484(.A(KEYINPUT16), .B(G8gat), .Z(new_n686));
  INV_X1    g485(.A(new_n679), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n677), .A2(KEYINPUT102), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n423), .B(new_n686), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT42), .ZN(new_n690));
  OAI21_X1  g489(.A(KEYINPUT104), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n258), .B1(new_n678), .B2(new_n679), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n692), .A2(new_n693), .A3(KEYINPUT42), .A4(new_n686), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(G8gat), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT42), .B1(new_n692), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n689), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n695), .A2(new_n698), .ZN(G1325gat));
  AOI21_X1  g498(.A(G15gat), .B1(new_n680), .B2(new_n383), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n466), .B(KEYINPUT36), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n701), .A2(G15gat), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n700), .B1(new_n680), .B2(new_n702), .ZN(G1326gat));
  INV_X1    g502(.A(new_n438), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n680), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(KEYINPUT43), .B(G22gat), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1327gat));
  NAND2_X1  g506(.A1(new_n475), .A2(new_n561), .ZN(new_n708));
  INV_X1    g507(.A(new_n600), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(new_n675), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n643), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT105), .Z(new_n712));
  NOR2_X1   g511(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n713), .A2(new_n478), .A3(new_n683), .ZN(new_n714));
  XOR2_X1   g513(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n469), .A2(new_n473), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n429), .B1(new_n419), .B2(new_n420), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n717), .B1(new_n718), .B2(new_n422), .ZN(new_n719));
  OAI21_X1  g518(.A(KEYINPUT44), .B1(new_n719), .B2(new_n646), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n475), .A2(new_n721), .A3(new_n643), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(new_n561), .A3(new_n710), .ZN(new_n724));
  INV_X1    g523(.A(new_n683), .ZN(new_n725));
  OAI21_X1  g524(.A(G29gat), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n716), .A2(new_n726), .ZN(G1328gat));
  NAND3_X1  g526(.A1(new_n713), .A2(new_n479), .A3(new_n423), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n728), .B(KEYINPUT46), .Z(new_n729));
  OAI21_X1  g528(.A(G36gat), .B1(new_n724), .B2(new_n258), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(G1329gat));
  OAI21_X1  g530(.A(G43gat), .B1(new_n724), .B2(new_n468), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n713), .A2(new_n488), .A3(new_n383), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT47), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n732), .A2(KEYINPUT47), .A3(new_n733), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(G1330gat));
  OAI21_X1  g537(.A(G50gat), .B1(new_n724), .B2(new_n438), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n438), .A2(G50gat), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT107), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n713), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT48), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n739), .A2(KEYINPUT48), .A3(new_n742), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(G1331gat));
  INV_X1    g546(.A(new_n649), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n561), .A2(new_n674), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n475), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n683), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g552(.A1(new_n750), .A2(new_n258), .ZN(new_n754));
  NOR2_X1   g553(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n755));
  AND2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(new_n754), .B2(new_n755), .ZN(G1333gat));
  OAI21_X1  g557(.A(new_n567), .B1(new_n750), .B2(new_n466), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n701), .A2(G71gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(new_n750), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1334gat));
  NOR2_X1   g562(.A1(new_n750), .A2(new_n438), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(new_n568), .ZN(G1335gat));
  NOR2_X1   g564(.A1(new_n709), .A2(new_n561), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n767), .A2(new_n674), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n769), .B1(new_n720), .B2(new_n722), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(G85gat), .B1(new_n771), .B2(new_n725), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n475), .A2(KEYINPUT51), .A3(new_n643), .A4(new_n766), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n646), .B1(new_n431), .B2(new_n474), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n776), .A2(KEYINPUT109), .A3(KEYINPUT51), .A4(new_n766), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT110), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n776), .A2(new_n766), .ZN(new_n781));
  AOI22_X1  g580(.A1(new_n778), .A2(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n775), .A2(KEYINPUT110), .A3(new_n777), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n683), .A2(new_n332), .A3(new_n675), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n772), .B1(new_n784), .B2(new_n785), .ZN(G1336gat));
  NAND3_X1  g585(.A1(new_n423), .A2(new_n675), .A3(new_n616), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n781), .A2(new_n780), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n787), .B1(new_n778), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n616), .B1(new_n770), .B2(new_n423), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT52), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n721), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n719), .A2(KEYINPUT44), .A3(new_n646), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n423), .B(new_n768), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT111), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n770), .A2(new_n796), .A3(new_n423), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n795), .A2(G92gat), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n787), .B1(new_n782), .B2(new_n783), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n791), .B1(new_n800), .B2(new_n801), .ZN(G1337gat));
  OAI21_X1  g601(.A(G99gat), .B1(new_n771), .B2(new_n468), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n383), .A2(new_n623), .A3(new_n675), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n803), .B1(new_n784), .B2(new_n804), .ZN(G1338gat));
  NAND3_X1  g604(.A1(new_n704), .A2(new_n624), .A3(new_n675), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n778), .B2(new_n788), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n624), .B1(new_n770), .B2(new_n704), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT53), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n806), .B1(new_n782), .B2(new_n783), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n808), .A2(KEYINPUT53), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(G1339gat));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n665), .B(new_n650), .C1(new_n659), .C2(new_n661), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n664), .A2(KEYINPUT54), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n662), .A2(new_n816), .A3(new_n663), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n815), .A2(KEYINPUT55), .A3(new_n669), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n671), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n817), .A2(new_n669), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT55), .B1(new_n820), .B2(new_n815), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n819), .A2(new_n821), .A3(new_n646), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n545), .A2(new_n541), .A3(new_n532), .A4(new_n552), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n558), .A2(new_n526), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n535), .A2(new_n540), .A3(new_n534), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n551), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n813), .B1(new_n822), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n664), .A2(KEYINPUT54), .A3(new_n814), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n817), .A2(new_n669), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n833), .A2(new_n643), .A3(new_n671), .A4(new_n818), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n834), .A2(KEYINPUT112), .A3(new_n827), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n819), .A2(new_n821), .ZN(new_n836));
  AOI22_X1  g635(.A1(new_n836), .A2(new_n561), .B1(new_n675), .B2(new_n828), .ZN(new_n837));
  OAI22_X1  g636(.A1(new_n829), .A2(new_n835), .B1(new_n837), .B2(new_n643), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n600), .ZN(new_n839));
  INV_X1    g638(.A(new_n561), .ZN(new_n840));
  AND4_X1   g639(.A1(new_n840), .A2(new_n644), .A3(new_n648), .A4(new_n674), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(KEYINPUT113), .A3(new_n438), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT113), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n841), .B1(new_n838), .B2(new_n600), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n845), .B1(new_n846), .B2(new_n704), .ZN(new_n847));
  AND3_X1   g646(.A1(new_n844), .A2(new_n383), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n725), .A2(new_n423), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(G113gat), .B1(new_n850), .B2(new_n840), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n846), .A2(new_n725), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n418), .A2(new_n423), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n286), .A3(new_n561), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n851), .A2(new_n856), .ZN(G1340gat));
  OAI21_X1  g656(.A(G120gat), .B1(new_n850), .B2(new_n674), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n855), .A2(new_n284), .A3(new_n675), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1341gat));
  NOR3_X1   g659(.A1(new_n850), .A2(new_n291), .A3(new_n600), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n855), .A2(KEYINPUT114), .A3(new_n709), .ZN(new_n862));
  AOI21_X1  g661(.A(KEYINPUT114), .B1(new_n855), .B2(new_n709), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(G127gat), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n861), .B1(new_n862), .B2(new_n864), .ZN(G1342gat));
  OAI21_X1  g664(.A(G134gat), .B1(new_n850), .B2(new_n646), .ZN(new_n866));
  AND4_X1   g665(.A1(new_n289), .A2(new_n852), .A3(new_n643), .A4(new_n853), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(KEYINPUT56), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT115), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n866), .A2(new_n868), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(G1343gat));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n874), .B1(new_n846), .B2(new_n438), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT116), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n836), .A2(new_n813), .A3(new_n643), .A4(new_n828), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT112), .B1(new_n834), .B2(new_n827), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n880), .B1(new_n831), .B2(new_n832), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n820), .A2(KEYINPUT117), .A3(new_n815), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(new_n830), .A3(new_n882), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n818), .A2(new_n671), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n883), .A2(new_n561), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n828), .A2(new_n675), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n643), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n879), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI211_X1 g688(.A(KEYINPUT118), .B(new_n643), .C1(new_n885), .C2(new_n886), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n600), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n842), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n438), .A2(new_n874), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT116), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n895), .B(new_n874), .C1(new_n846), .C2(new_n438), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n876), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n725), .A2(new_n423), .A3(new_n701), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(G141gat), .B1(new_n899), .B2(new_n840), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n701), .A2(new_n438), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n423), .B1(new_n901), .B2(KEYINPUT119), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n852), .B(new_n902), .C1(KEYINPUT119), .C2(new_n901), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n269), .A3(new_n561), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n900), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(KEYINPUT58), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT58), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n900), .A2(new_n908), .A3(new_n905), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(G1344gat));
  NAND3_X1  g709(.A1(new_n897), .A2(new_n675), .A3(new_n898), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n267), .A2(KEYINPUT59), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT120), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n911), .A2(new_n915), .A3(new_n912), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n874), .B1(new_n843), .B2(new_n704), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n834), .A2(new_n827), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n600), .B1(new_n887), .B2(new_n918), .ZN(new_n919));
  AOI211_X1 g718(.A(KEYINPUT57), .B(new_n438), .C1(new_n919), .C2(new_n842), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n921), .A2(new_n675), .A3(new_n898), .ZN(new_n922));
  OAI21_X1  g721(.A(KEYINPUT59), .B1(new_n922), .B2(new_n267), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n914), .A2(new_n916), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n904), .A2(new_n267), .A3(new_n675), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1345gat));
  NOR3_X1   g725(.A1(new_n899), .A2(new_n264), .A3(new_n600), .ZN(new_n927));
  AOI21_X1  g726(.A(G155gat), .B1(new_n904), .B2(new_n709), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n927), .A2(new_n928), .ZN(G1346gat));
  NAND3_X1  g728(.A1(new_n904), .A2(new_n278), .A3(new_n643), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT121), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n931), .B1(new_n899), .B2(new_n646), .ZN(new_n932));
  INV_X1    g731(.A(new_n278), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n899), .A2(new_n931), .A3(new_n646), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n930), .B1(new_n934), .B2(new_n935), .ZN(G1347gat));
  NOR2_X1   g735(.A1(new_n683), .A2(new_n258), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n844), .A2(new_n847), .A3(new_n383), .A4(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(G169gat), .B1(new_n938), .B2(new_n840), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n846), .A2(new_n683), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n418), .A2(new_n258), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OR2_X1    g741(.A1(new_n840), .A2(G169gat), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n939), .B1(new_n942), .B2(new_n943), .ZN(G1348gat));
  NAND2_X1  g743(.A1(new_n675), .A2(G176gat), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n938), .A2(new_n945), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n946), .A2(KEYINPUT122), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n946), .A2(KEYINPUT122), .ZN(new_n948));
  INV_X1    g747(.A(new_n942), .ZN(new_n949));
  AOI21_X1  g748(.A(G176gat), .B1(new_n949), .B2(new_n675), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n947), .A2(new_n948), .A3(new_n950), .ZN(G1349gat));
  OAI21_X1  g750(.A(G183gat), .B1(new_n938), .B2(new_n600), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n949), .A2(new_n228), .A3(new_n709), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g754(.A1(new_n949), .A2(new_n229), .A3(new_n643), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n848), .A2(new_n643), .A3(new_n937), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT61), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n957), .A2(new_n958), .A3(G190gat), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n958), .B1(new_n957), .B2(G190gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(G1351gat));
  NAND2_X1  g760(.A1(new_n901), .A2(new_n423), .ZN(new_n962));
  XOR2_X1   g761(.A(new_n962), .B(KEYINPUT123), .Z(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(new_n940), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT124), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n964), .B(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(G197gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n966), .A2(new_n967), .A3(new_n561), .ZN(new_n968));
  OR3_X1    g767(.A1(new_n917), .A2(KEYINPUT125), .A3(new_n920), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n683), .A2(new_n258), .A3(new_n701), .ZN(new_n970));
  OAI21_X1  g769(.A(KEYINPUT125), .B1(new_n917), .B2(new_n920), .ZN(new_n971));
  AND3_X1   g770(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n972), .A2(new_n561), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n968), .B1(new_n973), .B2(new_n967), .ZN(G1352gat));
  XNOR2_X1  g773(.A(KEYINPUT126), .B(G204gat), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n964), .A2(new_n674), .A3(new_n975), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n976), .B(KEYINPUT62), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n972), .A2(new_n675), .ZN(new_n978));
  INV_X1    g777(.A(new_n975), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(G1353gat));
  INV_X1    g779(.A(G211gat), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n970), .A2(new_n709), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n981), .B1(new_n921), .B2(new_n982), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT127), .ZN(new_n984));
  OR3_X1    g783(.A1(new_n983), .A2(new_n984), .A3(KEYINPUT63), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n984), .B1(new_n983), .B2(KEYINPUT63), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n983), .A2(KEYINPUT63), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n966), .A2(new_n981), .A3(new_n709), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n988), .A2(new_n989), .ZN(G1354gat));
  AOI21_X1  g789(.A(G218gat), .B1(new_n966), .B2(new_n643), .ZN(new_n991));
  AND2_X1   g790(.A1(new_n643), .A2(G218gat), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n991), .B1(new_n972), .B2(new_n992), .ZN(G1355gat));
endmodule


