//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 1 0 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n525, new_n526, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n549, new_n551, new_n552, new_n553,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n600, new_n603, new_n605,
    new_n606, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1219, new_n1220, new_n1221;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT65), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT66), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT67), .B(G69), .Z(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT68), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G101), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n467), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n466), .B1(new_n462), .B2(new_n474), .ZN(G160));
  OAI21_X1  g050(.A(G2104), .B1(new_n462), .B2(G112), .ZN(new_n476));
  INV_X1    g051(.A(G100), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(new_n462), .ZN(new_n478));
  XOR2_X1   g053(.A(new_n478), .B(KEYINPUT69), .Z(new_n479));
  NOR2_X1   g054(.A1(new_n472), .A2(new_n462), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n472), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NAND2_X1  g060(.A1(G114), .A2(G2104), .ZN(new_n486));
  INV_X1    g061(.A(G126), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n486), .B1(new_n472), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n468), .A2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G102), .ZN(new_n491));
  AND2_X1   g066(.A1(KEYINPUT70), .A2(G138), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n469), .A2(new_n471), .A3(new_n492), .A4(new_n462), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n463), .A2(KEYINPUT4), .A3(new_n462), .A4(new_n492), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n489), .A2(new_n491), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT71), .B1(new_n501), .B2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(new_n499), .A3(G543), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n500), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  OR3_X1    g082(.A1(new_n506), .A2(KEYINPUT72), .A3(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n509), .A2(G543), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n511), .A2(G88), .B1(G50), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g088(.A(KEYINPUT72), .B1(new_n506), .B2(new_n507), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n508), .A2(new_n513), .A3(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  NAND2_X1  g091(.A1(new_n511), .A2(G89), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT7), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n519), .A2(KEYINPUT7), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n512), .A2(G51), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n517), .A2(new_n518), .A3(new_n522), .ZN(G286));
  INV_X1    g098(.A(G286), .ZN(G168));
  XNOR2_X1  g099(.A(KEYINPUT73), .B(G52), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n512), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G90), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n527), .B2(new_n510), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n507), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n529), .A2(new_n532), .ZN(G301));
  INV_X1    g108(.A(G301), .ZN(G171));
  NAND3_X1  g109(.A1(new_n509), .A2(G43), .A3(G543), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n536), .B1(new_n511), .B2(G81), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT74), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n502), .A2(new_n504), .ZN(new_n539));
  INV_X1    g114(.A(new_n500), .ZN(new_n540));
  AND3_X1   g115(.A1(new_n539), .A2(G56), .A3(new_n540), .ZN(new_n541));
  AND2_X1   g116(.A1(G68), .A2(G543), .ZN(new_n542));
  OAI211_X1 g117(.A(new_n538), .B(G651), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n542), .B1(new_n505), .B2(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(KEYINPUT74), .B1(new_n544), .B2(new_n507), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n537), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT75), .ZN(G188));
  INV_X1    g129(.A(KEYINPUT9), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n512), .A2(new_n555), .A3(G53), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n509), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  OAI21_X1  g133(.A(KEYINPUT9), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n511), .A2(G91), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n505), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n560), .B(new_n561), .C1(new_n507), .C2(new_n562), .ZN(G299));
  NAND2_X1  g138(.A1(new_n512), .A2(G49), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n505), .A2(G87), .A3(new_n509), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(G288));
  AND3_X1   g142(.A1(new_n539), .A2(G61), .A3(new_n540), .ZN(new_n568));
  NAND2_X1  g143(.A1(G73), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n539), .A2(G86), .A3(new_n509), .A4(new_n540), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n509), .A2(G48), .A3(G543), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n571), .A2(new_n575), .ZN(G305));
  INV_X1    g151(.A(G85), .ZN(new_n577));
  INV_X1    g152(.A(G47), .ZN(new_n578));
  OAI22_X1  g153(.A1(new_n510), .A2(new_n577), .B1(new_n578), .B2(new_n557), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n505), .A2(G60), .ZN(new_n580));
  NAND2_X1  g155(.A1(G72), .A2(G543), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n507), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OR3_X1    g157(.A1(new_n579), .A2(new_n582), .A3(KEYINPUT76), .ZN(new_n583));
  OAI21_X1  g158(.A(KEYINPUT76), .B1(new_n579), .B2(new_n582), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  INV_X1    g161(.A(G92), .ZN(new_n587));
  OAI21_X1  g162(.A(KEYINPUT10), .B1(new_n510), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT10), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n505), .A2(new_n589), .A3(G92), .A4(new_n509), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n512), .A2(G54), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n505), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n593), .B2(new_n507), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT77), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n586), .B1(new_n596), .B2(G868), .ZN(G284));
  OAI21_X1  g172(.A(new_n586), .B1(new_n596), .B2(G868), .ZN(G321));
  NAND2_X1  g173(.A1(G286), .A2(G868), .ZN(new_n599));
  INV_X1    g174(.A(G299), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(G868), .ZN(G280));
  XOR2_X1   g176(.A(G280), .B(KEYINPUT78), .Z(G297));
  XOR2_X1   g177(.A(KEYINPUT79), .B(G559), .Z(new_n603));
  OAI21_X1  g178(.A(new_n596), .B1(G860), .B2(new_n603), .ZN(G148));
  NAND2_X1  g179(.A1(new_n596), .A2(new_n603), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G868), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g182(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g183(.A1(new_n482), .A2(G135), .ZN(new_n609));
  OR2_X1    g184(.A1(G99), .A2(G2105), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n610), .B(G2104), .C1(G111), .C2(new_n462), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(G123), .B2(new_n480), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(G2096), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(KEYINPUT12), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT12), .ZN(new_n617));
  NAND4_X1  g192(.A1(new_n617), .A2(new_n462), .A3(KEYINPUT3), .A4(G2104), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2100), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n614), .A2(new_n621), .ZN(G156));
  XNOR2_X1  g197(.A(G2427), .B(G2430), .ZN(new_n623));
  OR2_X1    g198(.A1(KEYINPUT15), .A2(G2435), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT80), .ZN(new_n625));
  NAND2_X1  g200(.A1(KEYINPUT15), .A2(G2435), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(G2438), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n625), .B1(new_n624), .B2(new_n626), .ZN(new_n630));
  NOR3_X1   g205(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n624), .A2(new_n626), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(KEYINPUT80), .ZN(new_n633));
  AOI21_X1  g208(.A(G2438), .B1(new_n633), .B2(new_n627), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n623), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n629), .B1(new_n628), .B2(new_n630), .ZN(new_n636));
  INV_X1    g211(.A(new_n623), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n633), .A2(G2438), .A3(new_n627), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  INV_X1    g220(.A(new_n643), .ZN(new_n646));
  NAND4_X1  g221(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n639), .A4(new_n646), .ZN(new_n647));
  AND3_X1   g222(.A1(new_n644), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n645), .B1(new_n644), .B2(new_n647), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G1341), .B(G1348), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT83), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n650), .A2(KEYINPUT83), .A3(new_n652), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(G14), .ZN(new_n658));
  OAI21_X1  g233(.A(KEYINPUT82), .B1(new_n650), .B2(new_n652), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT82), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n660), .B(new_n651), .C1(new_n648), .C2(new_n649), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n658), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n657), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G401));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n665), .B1(new_n668), .B2(KEYINPUT18), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G2096), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(G2100), .Z(new_n671));
  AND2_X1   g246(.A1(new_n668), .A2(KEYINPUT17), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n666), .A2(new_n667), .ZN(new_n673));
  AOI21_X1  g248(.A(KEYINPUT18), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n671), .B(new_n674), .ZN(G227));
  XNOR2_X1  g250(.A(KEYINPUT84), .B(G1986), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  OR2_X1    g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n681), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n683), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n679), .A2(new_n682), .A3(new_n684), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n687), .B(new_n688), .C1(new_n686), .C2(new_n685), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n691), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  INV_X1    g269(.A(G1981), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  AND3_X1   g272(.A1(new_n692), .A2(new_n693), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n697), .B1(new_n692), .B2(new_n693), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n677), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n692), .A2(new_n693), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(new_n696), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n692), .A2(new_n693), .A3(new_n697), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n702), .A2(new_n676), .A3(new_n703), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n700), .A2(new_n704), .ZN(G229));
  AND2_X1   g280(.A1(KEYINPUT85), .A2(G29), .ZN(new_n706));
  NOR2_X1   g281(.A1(KEYINPUT85), .A2(G29), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n497), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n708), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G27), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n712), .A2(KEYINPUT96), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(KEYINPUT96), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G2078), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n713), .A2(G2078), .A3(new_n714), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT92), .B(G34), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT24), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n721), .A2(new_n710), .A3(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n723), .A2(KEYINPUT93), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G29), .B2(G160), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(KEYINPUT93), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G2084), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT95), .B(KEYINPUT31), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G11), .ZN(new_n731));
  OR2_X1    g306(.A1(G16), .A2(G21), .ZN(new_n732));
  INV_X1    g307(.A(G16), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(G286), .B2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G1966), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n731), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n717), .A2(new_n718), .A3(new_n729), .A4(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(G29), .A2(G33), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n490), .A2(G103), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT25), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(G115), .A2(G2104), .ZN(new_n742));
  INV_X1    g317(.A(G127), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n472), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G2105), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n482), .A2(G139), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n741), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n738), .B1(new_n748), .B2(G29), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n749), .A2(G2072), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n727), .A2(new_n728), .ZN(new_n751));
  INV_X1    g326(.A(G29), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT30), .B(G28), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n613), .A2(new_n708), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI221_X1 g329(.A(new_n754), .B1(new_n749), .B2(G2072), .C1(new_n734), .C2(new_n735), .ZN(new_n755));
  NOR4_X1   g330(.A1(new_n737), .A2(new_n750), .A3(new_n751), .A4(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n752), .A2(G32), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n482), .A2(G141), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n480), .A2(G129), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n490), .A2(G105), .ZN(new_n760));
  NAND3_X1  g335(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT26), .Z(new_n762));
  NAND4_X1  g337(.A1(new_n758), .A2(new_n759), .A3(new_n760), .A4(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n757), .B1(new_n764), .B2(new_n752), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT94), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT27), .B(G1996), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n733), .A2(G5), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G171), .B2(new_n733), .ZN(new_n770));
  INV_X1    g345(.A(G1961), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n756), .A2(new_n768), .A3(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT97), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n756), .A2(KEYINPUT97), .A3(new_n768), .A4(new_n772), .ZN(new_n776));
  NOR2_X1   g351(.A1(G4), .A2(G16), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n596), .B2(G16), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1348), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT98), .B(KEYINPUT23), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n733), .A2(G20), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G299), .B2(G16), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(G1956), .Z(new_n784));
  NOR2_X1   g359(.A1(new_n779), .A2(new_n784), .ZN(new_n785));
  AND3_X1   g360(.A1(new_n775), .A2(new_n776), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n710), .A2(KEYINPUT28), .A3(G26), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n463), .A2(G128), .A3(G2105), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n463), .A2(G140), .A3(new_n462), .ZN(new_n789));
  OR2_X1    g364(.A1(G104), .A2(G2105), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n790), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n791));
  AND3_X1   g366(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n787), .B1(new_n792), .B2(new_n752), .ZN(new_n793));
  AOI21_X1  g368(.A(KEYINPUT28), .B1(new_n710), .B2(G26), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT91), .ZN(new_n796));
  INV_X1    g371(.A(G2067), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT36), .ZN(new_n799));
  NOR2_X1   g374(.A1(G16), .A2(G22), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G166), .B2(G16), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT89), .B(G1971), .Z(new_n802));
  XOR2_X1   g377(.A(new_n801), .B(new_n802), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n505), .A2(G61), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n507), .B1(new_n804), .B2(new_n569), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n805), .A2(new_n574), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(G16), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT32), .ZN(new_n808));
  NOR2_X1   g383(.A1(G6), .A2(G16), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n807), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n808), .B1(new_n807), .B2(new_n810), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n695), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n813), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n815), .A2(G1981), .A3(new_n811), .ZN(new_n816));
  NOR2_X1   g391(.A1(G16), .A2(G23), .ZN(new_n817));
  INV_X1    g392(.A(G288), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(G16), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT33), .B(G1976), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  AND3_X1   g396(.A1(new_n814), .A2(new_n816), .A3(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT90), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n803), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n801), .B(new_n802), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n814), .A2(new_n816), .A3(new_n821), .ZN(new_n826));
  OAI21_X1  g401(.A(KEYINPUT90), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT34), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT34), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n824), .A2(new_n830), .A3(new_n827), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n710), .A2(G25), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n463), .A2(G119), .A3(G2105), .ZN(new_n834));
  INV_X1    g409(.A(G107), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n468), .B1(new_n835), .B2(G2105), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT86), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(G95), .B2(G2105), .ZN(new_n838));
  INV_X1    g413(.A(G95), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n839), .A2(new_n462), .A3(KEYINPUT86), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n836), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n463), .A2(new_n462), .ZN(new_n842));
  INV_X1    g417(.A(G131), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n834), .B(new_n841), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(KEYINPUT87), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n482), .A2(G131), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT87), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n846), .A2(new_n834), .A3(new_n847), .A4(new_n841), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n833), .B1(new_n850), .B2(new_n710), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT88), .ZN(new_n852));
  XNOR2_X1  g427(.A(KEYINPUT35), .B(G1991), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n733), .A2(G24), .ZN(new_n855));
  INV_X1    g430(.A(G290), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n855), .B1(new_n856), .B2(new_n733), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n857), .A2(G1986), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(G1986), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n854), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n799), .B1(new_n832), .B2(new_n861), .ZN(new_n862));
  AOI211_X1 g437(.A(KEYINPUT36), .B(new_n860), .C1(new_n829), .C2(new_n831), .ZN(new_n863));
  OAI211_X1 g438(.A(new_n786), .B(new_n798), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n733), .A2(G19), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n865), .B1(new_n547), .B2(new_n733), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(G1341), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n710), .A2(G35), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n868), .B1(G162), .B2(new_n710), .ZN(new_n869));
  XNOR2_X1  g444(.A(KEYINPUT29), .B(G2090), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  NOR3_X1   g446(.A1(new_n864), .A2(new_n867), .A3(new_n871), .ZN(G311));
  NAND3_X1  g447(.A1(new_n775), .A2(new_n776), .A3(new_n785), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n832), .A2(new_n861), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(KEYINPUT36), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n832), .A2(new_n799), .A3(new_n861), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n873), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n867), .ZN(new_n878));
  INV_X1    g453(.A(new_n871), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .A4(new_n798), .ZN(G150));
  XNOR2_X1  g455(.A(KEYINPUT99), .B(G55), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n512), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(G93), .ZN(new_n883));
  AOI22_X1  g458(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n884));
  OAI221_X1 g459(.A(new_n882), .B1(new_n510), .B2(new_n883), .C1(new_n884), .C2(new_n507), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(G860), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n886), .B(KEYINPUT37), .Z(new_n887));
  NAND2_X1  g462(.A1(new_n596), .A2(G559), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT39), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n882), .B1(new_n883), .B2(new_n510), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n884), .A2(new_n507), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n546), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n885), .A2(new_n537), .A3(new_n545), .A4(new_n543), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  XOR2_X1   g470(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n889), .B(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n887), .B1(new_n898), .B2(G860), .ZN(G145));
  INV_X1    g474(.A(G37), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n495), .A2(new_n496), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  AOI22_X1  g477(.A1(new_n488), .A2(G2105), .B1(G102), .B2(new_n490), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n486), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n906), .B1(new_n463), .B2(G126), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n491), .B1(new_n907), .B2(new_n462), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n792), .B1(new_n908), .B2(new_n901), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n905), .A2(new_n909), .A3(new_n747), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n747), .B1(new_n905), .B2(new_n909), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n763), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n905), .A2(new_n909), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n748), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n905), .A2(new_n909), .A3(new_n747), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(new_n764), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n480), .A2(G130), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n482), .A2(G142), .ZN(new_n919));
  OR2_X1    g494(.A1(G106), .A2(G2105), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n920), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT101), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n619), .B(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n845), .A2(new_n848), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n924), .B1(new_n845), .B2(new_n848), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n922), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n924), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n849), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n922), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n931), .A3(new_n925), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT102), .B1(new_n917), .B2(new_n933), .ZN(new_n934));
  NOR3_X1   g509(.A1(new_n926), .A2(new_n927), .A3(new_n922), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n931), .B1(new_n930), .B2(new_n925), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT102), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n937), .A2(new_n938), .A3(new_n916), .A4(new_n912), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n934), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n917), .A2(new_n933), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n613), .B(G160), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(new_n484), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n940), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT103), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n934), .A2(new_n939), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(new_n941), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n946), .B1(new_n934), .B2(new_n939), .ZN(new_n949));
  OAI211_X1 g524(.A(KEYINPUT104), .B(new_n943), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n940), .A2(KEYINPUT103), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n952), .A2(new_n941), .A3(new_n947), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT104), .B1(new_n953), .B2(new_n943), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n900), .B(new_n945), .C1(new_n951), .C2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT40), .ZN(G395));
  NAND3_X1  g531(.A1(new_n605), .A2(new_n894), .A3(new_n893), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n596), .A2(new_n603), .A3(new_n895), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n600), .A2(new_n595), .ZN(new_n959));
  OAI21_X1  g534(.A(G299), .B1(new_n594), .B2(new_n591), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n959), .A2(KEYINPUT41), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT41), .B1(new_n959), .B2(new_n960), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n957), .A2(new_n958), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n957), .A2(new_n958), .ZN(new_n965));
  INV_X1    g540(.A(new_n959), .ZN(new_n966));
  INV_X1    g541(.A(new_n960), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AOI22_X1  g543(.A1(new_n964), .A2(KEYINPUT105), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n965), .A2(KEYINPUT105), .A3(new_n968), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n970), .A2(KEYINPUT107), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(G305), .A2(new_n818), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n806), .A2(G288), .ZN(new_n974));
  AOI21_X1  g549(.A(G290), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(G290), .A2(new_n973), .A3(new_n974), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(G166), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n977), .ZN(new_n979));
  OAI21_X1  g554(.A(G303), .B1(new_n979), .B2(new_n975), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n981), .B(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT107), .ZN(new_n984));
  INV_X1    g559(.A(new_n971), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n984), .B1(new_n969), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n972), .A2(new_n983), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n983), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n988), .A2(KEYINPUT107), .A3(new_n970), .A4(new_n971), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n987), .A2(G868), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT108), .B1(new_n892), .B2(G868), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT108), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n992), .B1(new_n993), .B2(new_n990), .ZN(G295));
  OAI21_X1  g569(.A(new_n992), .B1(new_n993), .B2(new_n990), .ZN(G331));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT109), .ZN(new_n997));
  NAND3_X1  g572(.A1(G286), .A2(new_n532), .A3(new_n529), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n512), .A2(G51), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n521), .A2(new_n520), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n999), .A2(new_n518), .A3(new_n1000), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n1001), .B(new_n517), .C1(new_n531), .C2(new_n528), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n997), .B1(new_n895), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n895), .A2(new_n1003), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n893), .A2(new_n894), .A3(new_n998), .A4(new_n1002), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1004), .B1(new_n1007), .B2(new_n997), .ZN(new_n1008));
  OR2_X1    g583(.A1(new_n961), .A2(new_n962), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n996), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n968), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT109), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n963), .B(KEYINPUT110), .C1(new_n1012), .C2(new_n1004), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1010), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n981), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT43), .ZN(new_n1017));
  AOI22_X1  g592(.A1(new_n1008), .A2(new_n968), .B1(new_n963), .B2(new_n1007), .ZN(new_n1018));
  AOI21_X1  g593(.A(G37), .B1(new_n1018), .B2(new_n981), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1008), .A2(new_n968), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n963), .A2(new_n1007), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n981), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n900), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1018), .A2(new_n981), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT43), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT44), .B1(new_n1020), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  AOI211_X1 g604(.A(KEYINPUT111), .B(KEYINPUT44), .C1(new_n1020), .C2(new_n1026), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n1024), .A2(new_n1025), .A3(KEYINPUT43), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1024), .B1(new_n1015), .B2(new_n1014), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT44), .B1(new_n1032), .B2(new_n1017), .ZN(new_n1033));
  OAI22_X1  g608(.A1(new_n1029), .A2(new_n1030), .B1(new_n1031), .B2(new_n1033), .ZN(G397));
  INV_X1    g609(.A(G1384), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(new_n908), .B2(new_n901), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT45), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(G160), .A2(G40), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  OR3_X1    g616(.A1(new_n1041), .A2(G290), .A3(G1986), .ZN(new_n1042));
  NAND3_X1  g617(.A1(G290), .A2(G1986), .A3(new_n1040), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n1044), .B(KEYINPUT112), .ZN(new_n1045));
  INV_X1    g620(.A(G1996), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n764), .A2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n904), .B(new_n797), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n763), .A2(G1996), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n849), .A2(new_n853), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n849), .A2(new_n853), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(new_n1041), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1045), .A2(new_n1054), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n474), .A2(new_n462), .ZN(new_n1056));
  INV_X1    g631(.A(G40), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1056), .A2(new_n1057), .A3(new_n466), .ZN(new_n1058));
  OAI211_X1 g633(.A(KEYINPUT45), .B(new_n1035), .C1(new_n908), .C2(new_n901), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1038), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(new_n1061), .A3(new_n735), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT50), .B1(new_n497), .B2(new_n1035), .ZN(new_n1063));
  OAI211_X1 g638(.A(KEYINPUT50), .B(new_n1035), .C1(new_n908), .C2(new_n901), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n728), .B(new_n1058), .C1(new_n1063), .C2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1062), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1061), .B1(new_n1060), .B2(new_n735), .ZN(new_n1068));
  OAI21_X1  g643(.A(G8), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT51), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(G286), .A2(G8), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1069), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1060), .A2(new_n735), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT118), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1077), .A2(new_n1066), .A3(new_n1062), .ZN(new_n1078));
  OAI211_X1 g653(.A(G8), .B(new_n1072), .C1(new_n1078), .C2(G286), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1075), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1078), .A2(G8), .A3(G286), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  XNOR2_X1  g658(.A(KEYINPUT113), .B(G1971), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1060), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT114), .ZN(new_n1086));
  INV_X1    g661(.A(G2090), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1087), .B(new_n1058), .C1(new_n1063), .C2(new_n1065), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT114), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1060), .A2(new_n1089), .A3(new_n1084), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1086), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(G303), .A2(G8), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT55), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT55), .ZN(new_n1094));
  NAND3_X1  g669(.A1(G303), .A2(new_n1094), .A3(G8), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1091), .A2(new_n1097), .A3(G8), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT49), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n695), .B1(new_n571), .B2(new_n575), .ZN(new_n1100));
  XNOR2_X1  g675(.A(KEYINPUT115), .B(G1981), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n805), .A2(new_n574), .A3(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1099), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(G8), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1036), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1104), .B1(new_n1105), .B2(new_n1058), .ZN(new_n1106));
  OAI21_X1  g681(.A(G1981), .B1(new_n805), .B2(new_n574), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1107), .B(KEYINPUT49), .C1(G305), .C2(new_n1101), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1103), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n564), .A2(new_n565), .A3(G1976), .A4(new_n566), .ZN(new_n1110));
  INV_X1    g685(.A(G1976), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT52), .B1(G288), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1106), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  OAI211_X1 g688(.A(G8), .B(new_n1110), .C1(new_n1039), .C2(new_n1036), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT52), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1109), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(G8), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1116), .B1(new_n1118), .B2(new_n1096), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1098), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT45), .B1(new_n497), .B2(new_n1035), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1059), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1123), .A2(KEYINPUT53), .A3(new_n716), .A4(new_n1058), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n1060), .B2(G2078), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1058), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n771), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1124), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(G171), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1124), .A2(new_n1126), .A3(new_n1128), .A4(G301), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1132), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT54), .B1(new_n1134), .B2(KEYINPUT123), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1120), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1130), .A2(KEYINPUT54), .A3(new_n1132), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT124), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT124), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1130), .A2(new_n1139), .A3(KEYINPUT54), .A4(new_n1132), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1083), .A2(new_n1136), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT125), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(G299), .B(KEYINPUT57), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(KEYINPUT56), .B(G2072), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1123), .A2(new_n1058), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1127), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1146), .B(new_n1148), .C1(G1956), .C2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1148), .B1(new_n1149), .B2(G1956), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n1145), .ZN(new_n1152));
  XOR2_X1   g727(.A(new_n1152), .B(KEYINPUT119), .Z(new_n1153));
  NAND2_X1  g728(.A1(new_n1105), .A2(new_n1058), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1154), .A2(G2067), .ZN(new_n1155));
  INV_X1    g730(.A(G1348), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1155), .B1(new_n1156), .B2(new_n1127), .ZN(new_n1157));
  NOR3_X1   g732(.A1(new_n1157), .A2(new_n594), .A3(new_n591), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1150), .B1(new_n1153), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT61), .B1(new_n1151), .B2(new_n1145), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(new_n1150), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1157), .A2(KEYINPUT121), .A3(KEYINPUT60), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n595), .B1(new_n1157), .B2(KEYINPUT60), .ZN(new_n1163));
  AOI21_X1  g738(.A(KEYINPUT121), .B1(new_n1157), .B2(KEYINPUT60), .ZN(new_n1164));
  OR3_X1    g739(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT120), .ZN(new_n1166));
  XOR2_X1   g741(.A(KEYINPUT58), .B(G1341), .Z(new_n1167));
  NAND2_X1  g742(.A1(new_n1154), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1168), .B1(new_n1060), .B2(G1996), .ZN(new_n1169));
  AOI211_X1 g744(.A(new_n1166), .B(KEYINPUT59), .C1(new_n1169), .C2(new_n547), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n547), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT59), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1171), .B1(KEYINPUT120), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1170), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1163), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1161), .A2(new_n1165), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1159), .A2(new_n1177), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1083), .A2(new_n1136), .A3(new_n1141), .A4(KEYINPUT125), .ZN(new_n1179));
  AND3_X1   g754(.A1(new_n1144), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1083), .A2(KEYINPUT62), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1120), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT62), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1081), .A2(new_n1183), .A3(new_n1082), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1130), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1181), .A2(new_n1182), .A3(new_n1184), .A4(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1116), .B(KEYINPUT116), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1097), .B1(new_n1091), .B2(G8), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1078), .A2(G8), .A3(G168), .ZN(new_n1189));
  NOR3_X1   g764(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1190), .A2(KEYINPUT63), .A3(new_n1098), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT63), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1192), .B1(new_n1120), .B2(new_n1189), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1109), .A2(new_n1111), .A3(new_n818), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n1102), .B(KEYINPUT117), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  AOI22_X1  g771(.A1(new_n1191), .A2(new_n1193), .B1(new_n1106), .B2(new_n1196), .ZN(new_n1197));
  OR2_X1    g772(.A1(new_n1187), .A2(new_n1098), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1186), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1055), .B1(new_n1180), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1041), .B1(new_n764), .B2(new_n1048), .ZN(new_n1201));
  AND3_X1   g776(.A1(new_n1040), .A2(KEYINPUT46), .A3(new_n1046), .ZN(new_n1202));
  AOI21_X1  g777(.A(KEYINPUT46), .B1(new_n1040), .B2(new_n1046), .ZN(new_n1203));
  NOR3_X1   g778(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1204), .B(KEYINPUT47), .ZN(new_n1205));
  XOR2_X1   g780(.A(new_n1042), .B(KEYINPUT48), .Z(new_n1206));
  NOR2_X1   g781(.A1(new_n1206), .A2(new_n1054), .ZN(new_n1207));
  INV_X1    g782(.A(new_n1052), .ZN(new_n1208));
  OAI22_X1  g783(.A1(new_n1050), .A2(new_n1208), .B1(G2067), .B2(new_n904), .ZN(new_n1209));
  AOI211_X1 g784(.A(new_n1205), .B(new_n1207), .C1(new_n1040), .C2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1200), .A2(new_n1210), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g786(.A(G227), .B1(new_n657), .B2(new_n662), .ZN(new_n1213));
  AOI21_X1  g787(.A(new_n460), .B1(new_n700), .B2(new_n704), .ZN(new_n1214));
  AOI21_X1  g788(.A(KEYINPUT126), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g789(.A(new_n1215), .B1(new_n1020), .B2(new_n1026), .ZN(new_n1216));
  NAND3_X1  g790(.A1(new_n1213), .A2(new_n1214), .A3(KEYINPUT126), .ZN(new_n1217));
  NAND3_X1  g791(.A1(new_n1216), .A2(new_n955), .A3(new_n1217), .ZN(G225));
  NAND2_X1  g792(.A1(G225), .A2(KEYINPUT127), .ZN(new_n1219));
  INV_X1    g793(.A(KEYINPUT127), .ZN(new_n1220));
  NAND4_X1  g794(.A1(new_n1216), .A2(new_n955), .A3(new_n1220), .A4(new_n1217), .ZN(new_n1221));
  NAND2_X1  g795(.A1(new_n1219), .A2(new_n1221), .ZN(G308));
endmodule


