

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586;

  XNOR2_X1 U321 ( .A(n445), .B(n444), .ZN(n563) );
  XNOR2_X1 U322 ( .A(n391), .B(n390), .ZN(n553) );
  XOR2_X1 U323 ( .A(G43GAT), .B(KEYINPUT8), .Z(n289) );
  XOR2_X1 U324 ( .A(G92GAT), .B(KEYINPUT77), .Z(n290) );
  INV_X1 U325 ( .A(KEYINPUT96), .ZN(n455) );
  XNOR2_X1 U326 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U327 ( .A(n344), .B(n343), .ZN(n347) );
  XNOR2_X1 U328 ( .A(n326), .B(G204GAT), .ZN(n329) );
  OR2_X1 U329 ( .A1(n348), .A2(n349), .ZN(n351) );
  NOR2_X1 U330 ( .A1(n419), .A2(n418), .ZN(n420) );
  XNOR2_X1 U331 ( .A(n329), .B(n389), .ZN(n330) );
  XNOR2_X1 U332 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U333 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U334 ( .A(n334), .B(n333), .ZN(n337) );
  XNOR2_X1 U335 ( .A(n356), .B(n355), .ZN(n573) );
  NOR2_X1 U336 ( .A1(n568), .A2(n563), .ZN(n557) );
  XOR2_X1 U337 ( .A(KEYINPUT91), .B(n457), .Z(n540) );
  XNOR2_X1 U338 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n447) );
  XNOR2_X1 U339 ( .A(n448), .B(n447), .ZN(G1351GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n292) );
  XNOR2_X1 U341 ( .A(G169GAT), .B(KEYINPUT66), .ZN(n291) );
  XNOR2_X1 U342 ( .A(n292), .B(n291), .ZN(n301) );
  XOR2_X1 U343 ( .A(G183GAT), .B(KEYINPUT17), .Z(n294) );
  XNOR2_X1 U344 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n293) );
  XNOR2_X1 U345 ( .A(n294), .B(n293), .ZN(n332) );
  XOR2_X1 U346 ( .A(G120GAT), .B(n332), .Z(n299) );
  XOR2_X1 U347 ( .A(KEYINPUT0), .B(KEYINPUT83), .Z(n296) );
  XNOR2_X1 U348 ( .A(KEYINPUT82), .B(G127GAT), .ZN(n295) );
  XNOR2_X1 U349 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U350 ( .A(G113GAT), .B(n297), .Z(n437) );
  XNOR2_X1 U351 ( .A(G15GAT), .B(n437), .ZN(n298) );
  XNOR2_X1 U352 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U353 ( .A(n301), .B(n300), .ZN(n309) );
  NAND2_X1 U354 ( .A1(G227GAT), .A2(G233GAT), .ZN(n307) );
  XOR2_X1 U355 ( .A(G176GAT), .B(G71GAT), .Z(n303) );
  XNOR2_X1 U356 ( .A(G43GAT), .B(G190GAT), .ZN(n302) );
  XNOR2_X1 U357 ( .A(n303), .B(n302), .ZN(n305) );
  XOR2_X1 U358 ( .A(G134GAT), .B(G99GAT), .Z(n304) );
  XNOR2_X1 U359 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U361 ( .A(n309), .B(n308), .ZN(n521) );
  XOR2_X1 U362 ( .A(KEYINPUT86), .B(KEYINPUT23), .Z(n311) );
  NAND2_X1 U363 ( .A1(G228GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U364 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U365 ( .A(n312), .B(KEYINPUT24), .Z(n321) );
  XNOR2_X1 U366 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n313) );
  XNOR2_X1 U367 ( .A(n313), .B(KEYINPUT2), .ZN(n314) );
  XOR2_X1 U368 ( .A(n314), .B(KEYINPUT85), .Z(n316) );
  XNOR2_X1 U369 ( .A(G141GAT), .B(G148GAT), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n316), .B(n315), .ZN(n436) );
  XOR2_X1 U371 ( .A(KEYINPUT22), .B(G106GAT), .Z(n318) );
  XNOR2_X1 U372 ( .A(G22GAT), .B(G218GAT), .ZN(n317) );
  XNOR2_X1 U373 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U374 ( .A(n436), .B(n319), .ZN(n320) );
  XNOR2_X1 U375 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U376 ( .A(G204GAT), .B(G78GAT), .Z(n352) );
  XOR2_X1 U377 ( .A(n322), .B(n352), .Z(n325) );
  XOR2_X1 U378 ( .A(G50GAT), .B(G162GAT), .Z(n387) );
  XNOR2_X1 U379 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n323) );
  XNOR2_X1 U380 ( .A(n323), .B(G211GAT), .ZN(n335) );
  XNOR2_X1 U381 ( .A(n387), .B(n335), .ZN(n324) );
  XNOR2_X1 U382 ( .A(n325), .B(n324), .ZN(n460) );
  XOR2_X1 U383 ( .A(G169GAT), .B(G8GAT), .Z(n364) );
  XOR2_X1 U384 ( .A(G176GAT), .B(G64GAT), .Z(n345) );
  XOR2_X1 U385 ( .A(n345), .B(KEYINPUT92), .Z(n326) );
  INV_X1 U386 ( .A(G36GAT), .ZN(n474) );
  XNOR2_X1 U387 ( .A(G190GAT), .B(G218GAT), .ZN(n327) );
  XNOR2_X1 U388 ( .A(n290), .B(n327), .ZN(n328) );
  XNOR2_X1 U389 ( .A(n474), .B(n328), .ZN(n389) );
  XNOR2_X1 U390 ( .A(n364), .B(n330), .ZN(n334) );
  AND2_X1 U391 ( .A1(G226GAT), .A2(G233GAT), .ZN(n331) );
  INV_X1 U392 ( .A(n335), .ZN(n336) );
  XNOR2_X1 U393 ( .A(n337), .B(n336), .ZN(n512) );
  XOR2_X1 U394 ( .A(KEYINPUT46), .B(KEYINPUT109), .Z(n374) );
  XOR2_X1 U395 ( .A(KEYINPUT74), .B(G92GAT), .Z(n339) );
  XNOR2_X1 U396 ( .A(G148GAT), .B(G85GAT), .ZN(n338) );
  XNOR2_X1 U397 ( .A(n339), .B(n338), .ZN(n356) );
  XNOR2_X1 U398 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n340) );
  XNOR2_X1 U399 ( .A(n340), .B(KEYINPUT73), .ZN(n394) );
  INV_X1 U400 ( .A(n394), .ZN(n348) );
  XOR2_X1 U401 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n344) );
  NAND2_X1 U402 ( .A1(G230GAT), .A2(G233GAT), .ZN(n342) );
  INV_X1 U403 ( .A(KEYINPUT32), .ZN(n341) );
  XOR2_X1 U404 ( .A(G120GAT), .B(G57GAT), .Z(n425) );
  XNOR2_X1 U405 ( .A(n425), .B(n345), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n349) );
  NAND2_X1 U407 ( .A1(n348), .A2(n349), .ZN(n350) );
  NAND2_X1 U408 ( .A1(n351), .A2(n350), .ZN(n354) );
  XOR2_X1 U409 ( .A(G99GAT), .B(G106GAT), .Z(n386) );
  XNOR2_X1 U410 ( .A(n352), .B(n386), .ZN(n353) );
  XNOR2_X1 U411 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U412 ( .A(KEYINPUT41), .B(n573), .ZN(n527) );
  XOR2_X1 U413 ( .A(G113GAT), .B(G36GAT), .Z(n358) );
  XNOR2_X1 U414 ( .A(G29GAT), .B(G50GAT), .ZN(n357) );
  XNOR2_X1 U415 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U416 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n360) );
  XNOR2_X1 U417 ( .A(G197GAT), .B(G141GAT), .ZN(n359) );
  XNOR2_X1 U418 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U419 ( .A(n362), .B(n361), .ZN(n372) );
  XNOR2_X1 U420 ( .A(G15GAT), .B(G22GAT), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n363), .B(G1GAT), .ZN(n395) );
  XOR2_X1 U422 ( .A(n364), .B(n395), .Z(n366) );
  NAND2_X1 U423 ( .A1(G229GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U425 ( .A(n367), .B(KEYINPUT70), .Z(n370) );
  XNOR2_X1 U426 ( .A(KEYINPUT72), .B(KEYINPUT7), .ZN(n368) );
  XNOR2_X1 U427 ( .A(n289), .B(n368), .ZN(n376) );
  XNOR2_X1 U428 ( .A(n376), .B(KEYINPUT71), .ZN(n369) );
  XNOR2_X1 U429 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n372), .B(n371), .ZN(n470) );
  NAND2_X1 U431 ( .A1(n527), .A2(n470), .ZN(n373) );
  XNOR2_X1 U432 ( .A(n374), .B(n373), .ZN(n411) );
  XNOR2_X1 U433 ( .A(G29GAT), .B(G134GAT), .ZN(n375) );
  XNOR2_X1 U434 ( .A(n375), .B(G85GAT), .ZN(n429) );
  XNOR2_X1 U435 ( .A(n376), .B(n429), .ZN(n381) );
  XNOR2_X1 U436 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(n378) );
  AND2_X1 U437 ( .A1(G232GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U438 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U439 ( .A(n379), .B(KEYINPUT9), .Z(n380) );
  XNOR2_X1 U440 ( .A(n381), .B(n380), .ZN(n385) );
  XOR2_X1 U441 ( .A(KEYINPUT75), .B(KEYINPUT68), .Z(n383) );
  XNOR2_X1 U442 ( .A(KEYINPUT76), .B(KEYINPUT65), .ZN(n382) );
  XOR2_X1 U443 ( .A(n383), .B(n382), .Z(n384) );
  XNOR2_X1 U444 ( .A(n385), .B(n384), .ZN(n391) );
  XNOR2_X1 U445 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U446 ( .A(KEYINPUT14), .B(KEYINPUT79), .Z(n393) );
  XNOR2_X1 U447 ( .A(KEYINPUT80), .B(KEYINPUT15), .ZN(n392) );
  XNOR2_X1 U448 ( .A(n393), .B(n392), .ZN(n401) );
  XNOR2_X1 U449 ( .A(n395), .B(n394), .ZN(n399) );
  XOR2_X1 U450 ( .A(KEYINPUT81), .B(KEYINPUT12), .Z(n397) );
  XNOR2_X1 U451 ( .A(G57GAT), .B(G64GAT), .ZN(n396) );
  XNOR2_X1 U452 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U453 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U454 ( .A(n401), .B(n400), .ZN(n409) );
  NAND2_X1 U455 ( .A1(G231GAT), .A2(G233GAT), .ZN(n407) );
  XOR2_X1 U456 ( .A(G78GAT), .B(G211GAT), .Z(n403) );
  XNOR2_X1 U457 ( .A(G8GAT), .B(G155GAT), .ZN(n402) );
  XNOR2_X1 U458 ( .A(n403), .B(n402), .ZN(n405) );
  XOR2_X1 U459 ( .A(G127GAT), .B(G183GAT), .Z(n404) );
  XNOR2_X1 U460 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U461 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U462 ( .A(n409), .B(n408), .ZN(n475) );
  NOR2_X1 U463 ( .A1(n553), .A2(n475), .ZN(n410) );
  NAND2_X1 U464 ( .A1(n411), .A2(n410), .ZN(n412) );
  XNOR2_X1 U465 ( .A(n412), .B(KEYINPUT47), .ZN(n413) );
  XNOR2_X1 U466 ( .A(n413), .B(KEYINPUT110), .ZN(n419) );
  XNOR2_X1 U467 ( .A(KEYINPUT78), .B(n553), .ZN(n535) );
  XNOR2_X1 U468 ( .A(KEYINPUT36), .B(n535), .ZN(n582) );
  NAND2_X1 U469 ( .A1(n582), .A2(n475), .ZN(n415) );
  XNOR2_X1 U470 ( .A(KEYINPUT67), .B(KEYINPUT45), .ZN(n414) );
  XNOR2_X1 U471 ( .A(n415), .B(n414), .ZN(n417) );
  INV_X1 U472 ( .A(n470), .ZN(n568) );
  AND2_X1 U473 ( .A1(n573), .A2(n568), .ZN(n416) );
  AND2_X1 U474 ( .A1(n417), .A2(n416), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n420), .B(KEYINPUT48), .ZN(n539) );
  NOR2_X1 U476 ( .A1(n512), .A2(n539), .ZN(n421) );
  XNOR2_X1 U477 ( .A(n421), .B(KEYINPUT54), .ZN(n440) );
  XOR2_X1 U478 ( .A(KEYINPUT90), .B(KEYINPUT4), .Z(n423) );
  XNOR2_X1 U479 ( .A(G1GAT), .B(G162GAT), .ZN(n422) );
  XNOR2_X1 U480 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U481 ( .A(n425), .B(n424), .Z(n427) );
  NAND2_X1 U482 ( .A1(G225GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U484 ( .A(n428), .B(KEYINPUT5), .Z(n431) );
  XNOR2_X1 U485 ( .A(n429), .B(KEYINPUT1), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U487 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n433) );
  XNOR2_X1 U488 ( .A(KEYINPUT87), .B(KEYINPUT6), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U490 ( .A(n435), .B(n434), .Z(n439) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n457) );
  NAND2_X1 U493 ( .A1(n440), .A2(n540), .ZN(n441) );
  XNOR2_X1 U494 ( .A(n441), .B(KEYINPUT64), .ZN(n565) );
  NOR2_X1 U495 ( .A1(n460), .A2(n565), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n442), .B(KEYINPUT55), .ZN(n443) );
  NOR2_X1 U497 ( .A1(n521), .A2(n443), .ZN(n445) );
  INV_X1 U498 ( .A(KEYINPUT120), .ZN(n444) );
  INV_X1 U499 ( .A(n563), .ZN(n446) );
  NAND2_X1 U500 ( .A1(n446), .A2(n535), .ZN(n448) );
  XOR2_X1 U501 ( .A(KEYINPUT95), .B(KEYINPUT26), .Z(n450) );
  NAND2_X1 U502 ( .A1(n460), .A2(n521), .ZN(n449) );
  XNOR2_X1 U503 ( .A(n450), .B(n449), .ZN(n566) );
  XOR2_X1 U504 ( .A(KEYINPUT27), .B(KEYINPUT93), .Z(n451) );
  XNOR2_X1 U505 ( .A(n512), .B(n451), .ZN(n462) );
  NOR2_X1 U506 ( .A1(n566), .A2(n462), .ZN(n542) );
  NOR2_X1 U507 ( .A1(n521), .A2(n512), .ZN(n452) );
  NOR2_X1 U508 ( .A1(n452), .A2(n460), .ZN(n453) );
  XOR2_X1 U509 ( .A(KEYINPUT25), .B(n453), .Z(n454) );
  NOR2_X1 U510 ( .A1(n542), .A2(n454), .ZN(n456) );
  XNOR2_X1 U511 ( .A(n456), .B(n455), .ZN(n458) );
  NAND2_X1 U512 ( .A1(n458), .A2(n457), .ZN(n459) );
  XOR2_X1 U513 ( .A(KEYINPUT97), .B(n459), .Z(n467) );
  XNOR2_X1 U514 ( .A(n460), .B(KEYINPUT69), .ZN(n461) );
  XNOR2_X1 U515 ( .A(n461), .B(KEYINPUT28), .ZN(n518) );
  INV_X1 U516 ( .A(n462), .ZN(n463) );
  NAND2_X1 U517 ( .A1(n518), .A2(n463), .ZN(n464) );
  NOR2_X1 U518 ( .A1(n540), .A2(n464), .ZN(n523) );
  XNOR2_X1 U519 ( .A(n523), .B(KEYINPUT94), .ZN(n465) );
  NAND2_X1 U520 ( .A1(n465), .A2(n521), .ZN(n466) );
  NAND2_X1 U521 ( .A1(n467), .A2(n466), .ZN(n477) );
  NAND2_X1 U522 ( .A1(n477), .A2(n582), .ZN(n468) );
  NOR2_X1 U523 ( .A1(n468), .A2(n475), .ZN(n469) );
  XNOR2_X1 U524 ( .A(n469), .B(KEYINPUT37), .ZN(n510) );
  NAND2_X1 U525 ( .A1(n470), .A2(n573), .ZN(n480) );
  NOR2_X1 U526 ( .A1(n510), .A2(n480), .ZN(n471) );
  XOR2_X1 U527 ( .A(KEYINPUT38), .B(n471), .Z(n494) );
  NOR2_X1 U528 ( .A1(n494), .A2(n512), .ZN(n472) );
  XNOR2_X1 U529 ( .A(n472), .B(KEYINPUT100), .ZN(n473) );
  XNOR2_X1 U530 ( .A(n474), .B(n473), .ZN(G1329GAT) );
  INV_X1 U531 ( .A(n475), .ZN(n579) );
  NOR2_X1 U532 ( .A1(n535), .A2(n579), .ZN(n476) );
  XNOR2_X1 U533 ( .A(KEYINPUT16), .B(n476), .ZN(n478) );
  NAND2_X1 U534 ( .A1(n478), .A2(n477), .ZN(n479) );
  XNOR2_X1 U535 ( .A(n479), .B(KEYINPUT98), .ZN(n496) );
  OR2_X1 U536 ( .A1(n496), .A2(n480), .ZN(n487) );
  NOR2_X1 U537 ( .A1(n540), .A2(n487), .ZN(n481) );
  XOR2_X1 U538 ( .A(n481), .B(KEYINPUT34), .Z(n482) );
  XNOR2_X1 U539 ( .A(G1GAT), .B(n482), .ZN(G1324GAT) );
  NOR2_X1 U540 ( .A1(n512), .A2(n487), .ZN(n483) );
  XOR2_X1 U541 ( .A(G8GAT), .B(n483), .Z(G1325GAT) );
  NOR2_X1 U542 ( .A1(n521), .A2(n487), .ZN(n485) );
  XNOR2_X1 U543 ( .A(KEYINPUT99), .B(KEYINPUT35), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U545 ( .A(G15GAT), .B(n486), .Z(G1326GAT) );
  NOR2_X1 U546 ( .A1(n518), .A2(n487), .ZN(n488) );
  XOR2_X1 U547 ( .A(G22GAT), .B(n488), .Z(G1327GAT) );
  XNOR2_X1 U548 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n490) );
  NOR2_X1 U549 ( .A1(n540), .A2(n494), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(G1328GAT) );
  NOR2_X1 U551 ( .A1(n494), .A2(n521), .ZN(n492) );
  XNOR2_X1 U552 ( .A(KEYINPUT101), .B(KEYINPUT40), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U554 ( .A(G43GAT), .B(n493), .ZN(G1330GAT) );
  NOR2_X1 U555 ( .A1(n518), .A2(n494), .ZN(n495) );
  XOR2_X1 U556 ( .A(G50GAT), .B(n495), .Z(G1331GAT) );
  XNOR2_X1 U557 ( .A(KEYINPUT102), .B(KEYINPUT42), .ZN(n500) );
  NAND2_X1 U558 ( .A1(n527), .A2(n568), .ZN(n509) );
  OR2_X1 U559 ( .A1(n496), .A2(n509), .ZN(n505) );
  NOR2_X1 U560 ( .A1(n540), .A2(n505), .ZN(n498) );
  XNOR2_X1 U561 ( .A(G57GAT), .B(KEYINPUT103), .ZN(n497) );
  XNOR2_X1 U562 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n500), .B(n499), .ZN(G1332GAT) );
  NOR2_X1 U564 ( .A1(n512), .A2(n505), .ZN(n501) );
  XOR2_X1 U565 ( .A(KEYINPUT104), .B(n501), .Z(n502) );
  XNOR2_X1 U566 ( .A(G64GAT), .B(n502), .ZN(G1333GAT) );
  NOR2_X1 U567 ( .A1(n521), .A2(n505), .ZN(n504) );
  XNOR2_X1 U568 ( .A(G71GAT), .B(KEYINPUT105), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n504), .B(n503), .ZN(G1334GAT) );
  NOR2_X1 U570 ( .A1(n518), .A2(n505), .ZN(n507) );
  XNOR2_X1 U571 ( .A(KEYINPUT43), .B(KEYINPUT106), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U573 ( .A(G78GAT), .B(n508), .ZN(G1335GAT) );
  OR2_X1 U574 ( .A1(n510), .A2(n509), .ZN(n517) );
  NOR2_X1 U575 ( .A1(n540), .A2(n517), .ZN(n511) );
  XOR2_X1 U576 ( .A(G85GAT), .B(n511), .Z(G1336GAT) );
  NOR2_X1 U577 ( .A1(n512), .A2(n517), .ZN(n514) );
  XNOR2_X1 U578 ( .A(G92GAT), .B(KEYINPUT107), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(G1337GAT) );
  NOR2_X1 U580 ( .A1(n521), .A2(n517), .ZN(n515) );
  XOR2_X1 U581 ( .A(KEYINPUT108), .B(n515), .Z(n516) );
  XNOR2_X1 U582 ( .A(G99GAT), .B(n516), .ZN(G1338GAT) );
  NOR2_X1 U583 ( .A1(n518), .A2(n517), .ZN(n519) );
  XOR2_X1 U584 ( .A(KEYINPUT44), .B(n519), .Z(n520) );
  XNOR2_X1 U585 ( .A(G106GAT), .B(n520), .ZN(G1339GAT) );
  NOR2_X1 U586 ( .A1(n521), .A2(n539), .ZN(n522) );
  NAND2_X1 U587 ( .A1(n523), .A2(n522), .ZN(n534) );
  NOR2_X1 U588 ( .A1(n568), .A2(n534), .ZN(n524) );
  XOR2_X1 U589 ( .A(G113GAT), .B(n524), .Z(G1340GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n526) );
  XNOR2_X1 U591 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(n529) );
  INV_X1 U593 ( .A(n527), .ZN(n559) );
  NOR2_X1 U594 ( .A1(n559), .A2(n534), .ZN(n528) );
  XOR2_X1 U595 ( .A(n529), .B(n528), .Z(n530) );
  XNOR2_X1 U596 ( .A(KEYINPUT111), .B(n530), .ZN(G1341GAT) );
  NOR2_X1 U597 ( .A1(n579), .A2(n534), .ZN(n532) );
  XNOR2_X1 U598 ( .A(KEYINPUT50), .B(KEYINPUT114), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U600 ( .A(G127GAT), .B(n533), .Z(G1342GAT) );
  XOR2_X1 U601 ( .A(G134GAT), .B(KEYINPUT51), .Z(n538) );
  INV_X1 U602 ( .A(n534), .ZN(n536) );
  NAND2_X1 U603 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(G1343GAT) );
  NOR2_X1 U605 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U606 ( .A1(n542), .A2(n541), .ZN(n552) );
  NOR2_X1 U607 ( .A1(n568), .A2(n552), .ZN(n544) );
  XNOR2_X1 U608 ( .A(G141GAT), .B(KEYINPUT115), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n546) );
  XNOR2_X1 U611 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n550) );
  NOR2_X1 U613 ( .A1(n559), .A2(n552), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1345GAT) );
  NOR2_X1 U617 ( .A1(n579), .A2(n552), .ZN(n551) );
  XOR2_X1 U618 ( .A(G155GAT), .B(n551), .Z(G1346GAT) );
  XOR2_X1 U619 ( .A(G162GAT), .B(KEYINPUT119), .Z(n556) );
  INV_X1 U620 ( .A(n552), .ZN(n554) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1347GAT) );
  XNOR2_X1 U623 ( .A(n557), .B(KEYINPUT121), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G169GAT), .ZN(G1348GAT) );
  NOR2_X1 U625 ( .A1(n563), .A2(n559), .ZN(n561) );
  XNOR2_X1 U626 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(n562), .ZN(G1349GAT) );
  NOR2_X1 U629 ( .A1(n579), .A2(n563), .ZN(n564) );
  XOR2_X1 U630 ( .A(G183GAT), .B(n564), .Z(G1350GAT) );
  NOR2_X1 U631 ( .A1(n565), .A2(n566), .ZN(n567) );
  XOR2_X1 U632 ( .A(KEYINPUT122), .B(n567), .Z(n581) );
  NOR2_X1 U633 ( .A1(n568), .A2(n581), .ZN(n572) );
  XOR2_X1 U634 ( .A(KEYINPUT59), .B(KEYINPUT60), .Z(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  NOR2_X1 U638 ( .A1(n581), .A2(n573), .ZN(n578) );
  XOR2_X1 U639 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n575) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(KEYINPUT124), .B(n576), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n581), .ZN(n580) );
  XOR2_X1 U645 ( .A(G211GAT), .B(n580), .Z(G1354GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n585) );
  INV_X1 U647 ( .A(n581), .ZN(n583) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

