//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 0 0 0 0 0 1 1 1 1 0 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n548, new_n550, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n599, new_n600, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1139, new_n1140, new_n1141, new_n1142;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT66), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  INV_X1    g030(.A(new_n452), .ZN(new_n456));
  AOI22_X1  g031(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n459), .A2(G101), .A3(G2104), .ZN(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(new_n459), .ZN(new_n462));
  INV_X1    g037(.A(G137), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n461), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n459), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n464), .A2(new_n467), .ZN(G160));
  OAI21_X1  g043(.A(KEYINPUT69), .B1(G100), .B2(G2105), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  NOR3_X1   g045(.A1(KEYINPUT69), .A2(G100), .A3(G2105), .ZN(new_n471));
  OAI221_X1 g046(.A(G2104), .B1(G112), .B2(new_n459), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  XOR2_X1   g047(.A(new_n472), .B(KEYINPUT70), .Z(new_n473));
  INV_X1    g048(.A(new_n462), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n473), .B1(G136), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G124), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n477));
  INV_X1    g052(.A(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(KEYINPUT3), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n477), .B1(new_n482), .B2(new_n459), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n461), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n475), .B1(new_n476), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND4_X1  g063(.A1(new_n479), .A2(new_n481), .A3(G126), .A4(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n479), .A2(new_n481), .A3(G138), .A4(new_n459), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n461), .A2(new_n496), .A3(G138), .A4(new_n459), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n493), .B1(new_n495), .B2(new_n497), .ZN(G164));
  NAND2_X1  g073(.A1(G75), .A2(G543), .ZN(new_n499));
  XOR2_X1   g074(.A(KEYINPUT5), .B(G543), .Z(new_n500));
  INV_X1    g075(.A(G62), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G651), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n507), .A2(G88), .B1(new_n509), .B2(G50), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n510), .A2(new_n511), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n503), .B1(new_n512), .B2(new_n513), .ZN(G303));
  INV_X1    g089(.A(G303), .ZN(G166));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT7), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n504), .A2(new_n505), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G51), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(G89), .ZN(new_n522));
  NAND2_X1  g097(.A1(G63), .A2(G651), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n500), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n521), .A2(new_n524), .ZN(G168));
  XNOR2_X1  g100(.A(KEYINPUT5), .B(G543), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G52), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n518), .A2(new_n526), .ZN(new_n531));
  INV_X1    g106(.A(G90), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n530), .A2(new_n519), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT72), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT72), .ZN(new_n535));
  OAI221_X1 g110(.A(new_n535), .B1(new_n531), .B2(new_n532), .C1(new_n530), .C2(new_n519), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n529), .B1(new_n534), .B2(new_n536), .ZN(G171));
  NAND2_X1  g112(.A1(G68), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G56), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n500), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n528), .B1(new_n540), .B2(KEYINPUT73), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n541), .B1(KEYINPUT73), .B2(new_n540), .ZN(new_n542));
  XNOR2_X1  g117(.A(KEYINPUT74), .B(G43), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n507), .A2(G81), .B1(new_n509), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  XOR2_X1   g124(.A(KEYINPUT75), .B(KEYINPUT8), .Z(new_n550));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n550), .B(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n548), .A2(new_n552), .ZN(G188));
  NAND2_X1  g128(.A1(new_n526), .A2(G65), .ZN(new_n554));
  INV_X1    g129(.A(G78), .ZN(new_n555));
  OAI21_X1  g130(.A(KEYINPUT76), .B1(new_n555), .B2(new_n508), .ZN(new_n556));
  OR3_X1    g131(.A1(new_n555), .A2(new_n508), .A3(KEYINPUT76), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n554), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G651), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n507), .A2(G91), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n509), .A2(G53), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n562), .A2(new_n564), .ZN(G299));
  INV_X1    g140(.A(G171), .ZN(G301));
  INV_X1    g141(.A(G168), .ZN(G286));
  OAI21_X1  g142(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT77), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n507), .A2(G87), .B1(new_n509), .B2(G49), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(G288));
  NAND3_X1  g146(.A1(new_n518), .A2(G86), .A3(new_n526), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n518), .A2(G48), .A3(G543), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n526), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n574));
  OAI211_X1 g149(.A(new_n572), .B(new_n573), .C1(new_n574), .C2(new_n528), .ZN(G305));
  AOI22_X1  g150(.A1(new_n507), .A2(G85), .B1(new_n509), .B2(G47), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n528), .B2(new_n577), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT78), .ZN(G290));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n580));
  INV_X1    g155(.A(G868), .ZN(new_n581));
  NOR2_X1   g156(.A1(G171), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n526), .A2(G66), .ZN(new_n583));
  NAND2_X1  g158(.A1(G79), .A2(G543), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT80), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n528), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(G54), .B2(new_n509), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT81), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n507), .A2(G92), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT10), .Z(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  AOI211_X1 g166(.A(new_n580), .B(new_n582), .C1(new_n591), .C2(new_n581), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n580), .B2(new_n582), .ZN(G284));
  AOI21_X1  g168(.A(new_n592), .B1(new_n580), .B2(new_n582), .ZN(G321));
  NAND2_X1  g169(.A1(G286), .A2(G868), .ZN(new_n595));
  INV_X1    g170(.A(G299), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(G868), .ZN(G297));
  OAI21_X1  g172(.A(new_n595), .B1(new_n596), .B2(G868), .ZN(G280));
  INV_X1    g173(.A(new_n591), .ZN(new_n599));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(G860), .ZN(G148));
  NAND2_X1  g176(.A1(new_n599), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g180(.A1(new_n474), .A2(G2104), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT12), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(KEYINPUT13), .Z(new_n608));
  OR2_X1    g183(.A1(new_n608), .A2(G2100), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(G2100), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n485), .A2(G123), .ZN(new_n611));
  INV_X1    g186(.A(G111), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n612), .A2(KEYINPUT82), .A3(G2105), .ZN(new_n613));
  AOI21_X1  g188(.A(KEYINPUT82), .B1(new_n612), .B2(G2105), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n474), .A2(G135), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(G2096), .Z(new_n619));
  NAND3_X1  g194(.A1(new_n609), .A2(new_n610), .A3(new_n619), .ZN(G156));
  INV_X1    g195(.A(KEYINPUT14), .ZN(new_n621));
  XNOR2_X1  g196(.A(G2427), .B(G2438), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2430), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2435), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n621), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(new_n624), .B2(new_n623), .ZN(new_n626));
  XNOR2_X1  g201(.A(G1341), .B(G1348), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT84), .ZN(new_n628));
  XOR2_X1   g203(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n626), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G2451), .B(G2454), .Z(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n631), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(G14), .A3(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(G401));
  XNOR2_X1  g213(.A(G2084), .B(G2090), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2067), .B(G2678), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  AOI21_X1  g218(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT85), .B(KEYINPUT17), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n644), .B1(new_n646), .B2(new_n642), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT86), .Z(new_n648));
  NAND3_X1  g223(.A1(new_n646), .A2(new_n642), .A3(new_n640), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT87), .ZN(new_n650));
  NOR3_X1   g225(.A1(new_n642), .A2(new_n643), .A3(new_n639), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT18), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n648), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2100), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT88), .B(G2096), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(G227));
  XOR2_X1   g231(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n657));
  XNOR2_X1  g232(.A(G1971), .B(G1976), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1956), .B(G2474), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1961), .B(G1966), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT20), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n660), .B(new_n661), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n660), .A2(new_n661), .ZN(new_n666));
  MUX2_X1   g241(.A(new_n665), .B(new_n666), .S(new_n659), .Z(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT90), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G1981), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(G1986), .ZN(new_n671));
  INV_X1    g246(.A(G1981), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n669), .B(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(G1986), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT91), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n678), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n671), .A2(new_n675), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1991), .B(G1996), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n683), .B1(new_n679), .B2(new_n681), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(G229));
  INV_X1    g262(.A(G29), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G35), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G162), .B2(new_n688), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT29), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n691), .A2(KEYINPUT107), .A3(G2090), .ZN(new_n692));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G20), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT23), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(new_n596), .B2(new_n693), .ZN(new_n696));
  INV_X1    g271(.A(G1956), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n692), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(KEYINPUT107), .B1(new_n691), .B2(G2090), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT108), .ZN(new_n702));
  MUX2_X1   g277(.A(G24), .B(G290), .S(G16), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT93), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(G1986), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n688), .A2(G25), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n485), .A2(G119), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n474), .A2(G131), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n459), .A2(G107), .ZN(new_n709));
  OAI21_X1  g284(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n707), .B(new_n708), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT92), .Z(new_n712));
  OAI21_X1  g287(.A(new_n706), .B1(new_n712), .B2(new_n688), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT35), .B(G1991), .Z(new_n714));
  XOR2_X1   g289(.A(new_n713), .B(new_n714), .Z(new_n715));
  NOR2_X1   g290(.A1(new_n705), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n693), .A2(G22), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT97), .Z(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G166), .B2(new_n693), .ZN(new_n719));
  INV_X1    g294(.A(G1971), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n693), .A2(G6), .ZN(new_n722));
  INV_X1    g297(.A(G305), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(new_n693), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT94), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT32), .B(G1981), .Z(new_n726));
  OR2_X1    g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(new_n726), .ZN(new_n728));
  NOR2_X1   g303(.A1(G16), .A2(G23), .ZN(new_n729));
  INV_X1    g304(.A(G288), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(G16), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT33), .B(G1976), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n731), .B(new_n734), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n721), .A2(new_n727), .A3(new_n728), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(KEYINPUT34), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n736), .A2(KEYINPUT34), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n716), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT98), .B(KEYINPUT36), .Z(new_n740));
  OR2_X1    g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n739), .A2(new_n740), .ZN(new_n742));
  NOR2_X1   g317(.A1(G16), .A2(G19), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n546), .B2(G16), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT101), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(G1341), .Z(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G2090), .B2(new_n691), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT31), .B(G11), .ZN(new_n748));
  INV_X1    g323(.A(G28), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n749), .A2(KEYINPUT30), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT30), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n688), .B1(new_n751), .B2(G28), .ZN(new_n752));
  OAI221_X1 g327(.A(new_n748), .B1(new_n750), .B2(new_n752), .C1(new_n618), .C2(new_n688), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n688), .A2(G33), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT102), .B(KEYINPUT25), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n758), .A2(new_n459), .ZN(new_n759));
  AOI211_X1 g334(.A(new_n757), .B(new_n759), .C1(G139), .C2(new_n474), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n754), .B1(new_n760), .B2(new_n688), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G2072), .ZN(new_n762));
  INV_X1    g337(.A(G2084), .ZN(new_n763));
  NAND2_X1  g338(.A1(G160), .A2(G29), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT103), .B(KEYINPUT24), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(G34), .Z(new_n766));
  OAI21_X1  g341(.A(new_n764), .B1(G29), .B2(new_n766), .ZN(new_n767));
  AOI211_X1 g342(.A(new_n753), .B(new_n762), .C1(new_n763), .C2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n693), .A2(G21), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G168), .B2(new_n693), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT106), .B(G1966), .Z(new_n771));
  XOR2_X1   g346(.A(new_n770), .B(new_n771), .Z(new_n772));
  NAND3_X1  g347(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT26), .Z(new_n774));
  NAND3_X1  g349(.A1(new_n459), .A2(G105), .A3(G2104), .ZN(new_n775));
  INV_X1    g350(.A(G141), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n774), .B(new_n775), .C1(new_n776), .C2(new_n462), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n485), .B2(G129), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n778), .A2(new_n688), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n688), .B2(G32), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT27), .B(G1996), .ZN(new_n781));
  NOR2_X1   g356(.A1(G27), .A2(G29), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G164), .B2(G29), .ZN(new_n783));
  OAI22_X1  g358(.A1(new_n780), .A2(new_n781), .B1(G2078), .B2(new_n783), .ZN(new_n784));
  AOI211_X1 g359(.A(new_n772), .B(new_n784), .C1(G2078), .C2(new_n783), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n780), .A2(new_n781), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT105), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n693), .A2(G5), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G171), .B2(new_n693), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G1961), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n768), .A2(new_n785), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(G4), .A2(G16), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n599), .B2(G16), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT100), .B(G1348), .Z(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT99), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n793), .B(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n767), .A2(new_n763), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT104), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n688), .A2(G26), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT28), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n485), .A2(G128), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n459), .A2(G116), .ZN(new_n802));
  OAI21_X1  g377(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n474), .A2(G140), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n800), .B1(new_n806), .B2(G29), .ZN(new_n807));
  INV_X1    g382(.A(G2067), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n798), .A2(new_n809), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n796), .B(new_n810), .C1(G1961), .C2(new_n789), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n747), .A2(new_n791), .A3(new_n811), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n702), .A2(new_n741), .A3(new_n742), .A4(new_n812), .ZN(G150));
  INV_X1    g388(.A(G150), .ZN(G311));
  INV_X1    g389(.A(G55), .ZN(new_n815));
  INV_X1    g390(.A(G93), .ZN(new_n816));
  OAI22_X1  g391(.A1(new_n815), .A2(new_n519), .B1(new_n531), .B2(new_n816), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n526), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(new_n528), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(G860), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT37), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n591), .A2(new_n600), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT38), .ZN(new_n825));
  INV_X1    g400(.A(new_n820), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n545), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n820), .B1(new_n542), .B2(new_n544), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n825), .B(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT39), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT109), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n834), .B(new_n821), .C1(new_n831), .C2(new_n830), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n832), .A2(new_n833), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n823), .B1(new_n835), .B2(new_n836), .ZN(G145));
  XOR2_X1   g412(.A(new_n618), .B(G160), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n487), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n495), .A2(new_n497), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n489), .A2(new_n492), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n806), .B(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n778), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n760), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n474), .A2(G142), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n459), .A2(G118), .ZN(new_n848));
  OAI21_X1  g423(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(G130), .B2(new_n485), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(new_n607), .Z(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(new_n711), .Z(new_n853));
  OR2_X1    g428(.A1(new_n846), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT110), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n846), .A2(new_n855), .A3(new_n853), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n855), .B1(new_n846), .B2(new_n853), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n839), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n839), .B1(new_n846), .B2(new_n853), .ZN(new_n860));
  AOI21_X1  g435(.A(G37), .B1(new_n854), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g438(.A1(new_n826), .A2(new_n581), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n602), .B(new_n829), .ZN(new_n865));
  XNOR2_X1  g440(.A(KEYINPUT111), .B(KEYINPUT41), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n588), .A2(new_n596), .A3(new_n590), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n596), .B1(new_n588), .B2(new_n590), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n591), .A2(G299), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT41), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n588), .A2(new_n596), .A3(new_n590), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n865), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n868), .A2(new_n869), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n877), .B1(new_n878), .B2(new_n865), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT42), .ZN(new_n880));
  XNOR2_X1  g455(.A(G290), .B(G166), .ZN(new_n881));
  XNOR2_X1  g456(.A(G288), .B(new_n723), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n880), .B(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n864), .B1(new_n885), .B2(new_n581), .ZN(G295));
  OAI21_X1  g461(.A(new_n864), .B1(new_n885), .B2(new_n581), .ZN(G331));
  NOR3_X1   g462(.A1(new_n827), .A2(G171), .A3(new_n828), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(G171), .B1(new_n827), .B2(new_n828), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n890), .A3(G168), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n546), .A2(new_n820), .ZN(new_n892));
  INV_X1    g467(.A(new_n828), .ZN(new_n893));
  AOI21_X1  g468(.A(G301), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(G286), .B1(new_n894), .B2(new_n888), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(KEYINPUT112), .B1(new_n876), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT112), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n875), .A2(new_n898), .A3(new_n895), .A4(new_n891), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(new_n878), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n897), .A2(new_n883), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(G37), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n899), .A2(new_n900), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n883), .B1(new_n904), .B2(new_n897), .ZN(new_n905));
  OR3_X1    g480(.A1(new_n903), .A2(new_n905), .A3(KEYINPUT43), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n878), .A2(new_n867), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(KEYINPUT41), .B2(new_n878), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n900), .B1(new_n896), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n903), .B1(new_n884), .B2(new_n910), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n906), .B(KEYINPUT44), .C1(new_n907), .C2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT43), .B1(new_n903), .B2(new_n905), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n884), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n914), .A2(new_n901), .A3(new_n907), .A4(new_n902), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT113), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT113), .ZN(new_n919));
  AOI211_X1 g494(.A(new_n919), .B(KEYINPUT44), .C1(new_n913), .C2(new_n915), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n912), .B1(new_n918), .B2(new_n920), .ZN(G397));
  INV_X1    g496(.A(G1384), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n842), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT114), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT45), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(G164), .A2(G1384), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT114), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(G40), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n464), .A2(new_n467), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(G1996), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(KEYINPUT46), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n806), .A2(G2067), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n801), .A2(new_n808), .A3(new_n805), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n938), .A2(new_n844), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n935), .B1(new_n931), .B2(new_n939), .ZN(new_n940));
  XOR2_X1   g515(.A(new_n940), .B(KEYINPUT47), .Z(new_n941));
  NAND3_X1  g516(.A1(new_n932), .A2(new_n933), .A3(new_n778), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT115), .ZN(new_n943));
  OR2_X1    g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n778), .A2(new_n933), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n932), .B1(new_n938), .B2(new_n946), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n944), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n948), .A2(new_n712), .A3(new_n714), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n931), .B1(new_n949), .B2(new_n937), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n711), .B(new_n714), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n948), .B1(new_n931), .B2(new_n951), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n931), .A2(G1986), .A3(G290), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT48), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n941), .A2(new_n950), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT116), .B1(G164), .B2(G1384), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT116), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n842), .A2(new_n958), .A3(new_n922), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT50), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n957), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT117), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n957), .A2(new_n959), .A3(KEYINPUT117), .A4(new_n960), .ZN(new_n964));
  NAND2_X1  g539(.A1(G160), .A2(G40), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n965), .B1(KEYINPUT50), .B2(new_n923), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n963), .A2(new_n763), .A3(new_n964), .A4(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT45), .B1(new_n957), .B2(new_n959), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n842), .A2(KEYINPUT45), .A3(new_n922), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n930), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n771), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n967), .A2(G168), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(G8), .ZN(new_n973));
  AOI21_X1  g548(.A(G168), .B1(new_n967), .B2(new_n971), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT51), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n972), .A2(new_n976), .A3(G8), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n979));
  AND3_X1   g554(.A1(G303), .A2(G8), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n979), .B1(G303), .B2(G8), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT120), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n960), .B1(new_n957), .B2(new_n959), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n983), .B1(new_n984), .B2(new_n965), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n958), .B1(new_n842), .B2(new_n922), .ZN(new_n986));
  AOI211_X1 g561(.A(KEYINPUT116), .B(G1384), .C1(new_n840), .C2(new_n841), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT50), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n988), .A2(KEYINPUT120), .A3(new_n930), .ZN(new_n989));
  INV_X1    g564(.A(G2090), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n926), .A2(new_n960), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n985), .A2(new_n989), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(G164), .B2(G1384), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n994), .A2(new_n969), .A3(new_n930), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n720), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n982), .B1(new_n997), .B2(G8), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n963), .A2(new_n990), .A3(new_n964), .A4(new_n966), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(new_n996), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n1000), .A2(G8), .A3(new_n982), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n730), .A2(G1976), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n957), .A2(new_n959), .A3(new_n930), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(G8), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT52), .ZN(new_n1005));
  INV_X1    g580(.A(G1976), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT52), .B1(G288), .B2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1002), .A2(new_n1007), .A3(G8), .A4(new_n1003), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT119), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(G305), .B2(G1981), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT49), .ZN(new_n1012));
  NAND3_X1  g587(.A1(G305), .A2(new_n1012), .A3(G1981), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1012), .B1(G305), .B2(G1981), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1011), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1015), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1017), .A2(new_n1010), .A3(new_n1013), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1016), .A2(new_n1018), .A3(G8), .A4(new_n1003), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n1005), .A2(new_n1008), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1001), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n998), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n930), .B1(new_n926), .B2(new_n960), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1024), .B1(new_n962), .B2(new_n961), .ZN(new_n1025));
  AOI21_X1  g600(.A(G1961), .B1(new_n1025), .B2(new_n964), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n994), .A2(new_n969), .A3(new_n930), .ZN(new_n1027));
  INV_X1    g602(.A(G2078), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT53), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n969), .A2(KEYINPUT53), .A3(new_n1028), .A4(new_n930), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1030), .B1(new_n927), .B2(new_n925), .ZN(new_n1031));
  NOR4_X1   g606(.A1(new_n1026), .A2(G171), .A3(new_n1029), .A4(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n963), .A2(new_n964), .A3(new_n966), .ZN(new_n1033));
  INV_X1    g608(.A(G1961), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1029), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OR2_X1    g610(.A1(new_n968), .A2(new_n1030), .ZN(new_n1036));
  AOI21_X1  g611(.A(G301), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1023), .B1(new_n1032), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1035), .A2(G301), .A3(new_n1036), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n1026), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1039), .B(KEYINPUT54), .C1(new_n1040), .C2(G301), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n978), .A2(new_n1022), .A3(new_n1038), .A4(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n794), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1043), .B1(new_n1025), .B2(new_n964), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1003), .A2(G2067), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n599), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g621(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n1047));
  XNOR2_X1  g622(.A(new_n1047), .B(G2072), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1027), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n985), .A2(new_n989), .A3(new_n991), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1050), .B1(new_n1051), .B2(new_n697), .ZN(new_n1052));
  NAND2_X1  g627(.A1(KEYINPUT121), .A2(KEYINPUT57), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT121), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(G299), .A2(new_n1053), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT123), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n562), .A2(new_n564), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1058), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1046), .B1(new_n1052), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT124), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1052), .A2(new_n1066), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1063), .A2(new_n1064), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1064), .B1(new_n1063), .B2(new_n1067), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1067), .B(KEYINPUT61), .C1(new_n1052), .C2(new_n1062), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT61), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1051), .A2(new_n697), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1066), .B1(new_n1073), .B2(new_n1049), .ZN(new_n1074));
  AOI211_X1 g649(.A(new_n1050), .B(new_n1065), .C1(new_n1051), .C2(new_n697), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1072), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NOR4_X1   g651(.A1(new_n1044), .A2(KEYINPUT60), .A3(new_n591), .A4(new_n1045), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT125), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT58), .B(G1341), .Z(new_n1080));
  NAND2_X1  g655(.A1(new_n1003), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(G1996), .B2(new_n995), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1079), .B1(new_n1082), .B2(new_n546), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1027), .A2(new_n933), .B1(new_n1003), .B2(new_n1080), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1084), .A2(KEYINPUT125), .A3(new_n545), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1078), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT125), .B1(new_n1084), .B2(new_n545), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1082), .A2(new_n1079), .A3(new_n546), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1087), .A2(new_n1088), .A3(KEYINPUT59), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1077), .B1(new_n1086), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1046), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n1044), .A2(new_n599), .A3(new_n1045), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT60), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1071), .A2(new_n1076), .A3(new_n1090), .A4(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1042), .B1(new_n1070), .B2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n978), .A2(KEYINPUT62), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1022), .A2(new_n1037), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT62), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1098), .B1(new_n975), .B2(new_n977), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1096), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT63), .ZN(new_n1101));
  INV_X1    g676(.A(G8), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1102), .B1(new_n992), .B2(new_n996), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1001), .B(new_n1020), .C1(new_n1103), .C2(new_n982), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n967), .A2(new_n971), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1105), .A2(G8), .A3(G168), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1101), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1106), .A2(new_n1101), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1000), .A2(G8), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n980), .B2(new_n981), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1108), .A2(new_n1110), .A3(new_n1001), .A4(new_n1020), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1001), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1019), .A2(new_n1006), .A3(new_n730), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(G1981), .B2(G305), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1003), .A2(G8), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1113), .A2(new_n1020), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1112), .A2(new_n1117), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1095), .A2(new_n1100), .A3(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(G290), .B(new_n674), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1120), .A2(new_n931), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n952), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n1119), .A2(KEYINPUT126), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT126), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1042), .ZN(new_n1126));
  AND4_X1   g701(.A1(new_n1071), .A2(new_n1076), .A3(new_n1090), .A4(new_n1093), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1063), .A2(new_n1067), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT124), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1063), .A2(new_n1064), .A3(new_n1067), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1126), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1132));
  OR3_X1    g707(.A1(new_n1096), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1112), .A2(new_n1117), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1125), .B1(new_n1135), .B2(new_n1122), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n956), .B1(new_n1124), .B2(new_n1136), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g712(.A1(new_n637), .A2(new_n457), .ZN(new_n1139));
  NOR2_X1   g713(.A1(G227), .A2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g714(.A(new_n862), .B(new_n1140), .C1(new_n685), .C2(new_n686), .ZN(new_n1141));
  INV_X1    g715(.A(new_n916), .ZN(new_n1142));
  NOR2_X1   g716(.A1(new_n1141), .A2(new_n1142), .ZN(G308));
  OR2_X1    g717(.A1(new_n1141), .A2(new_n1142), .ZN(G225));
endmodule


