//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n559, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n610, new_n611,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT64), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g025(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT66), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n453), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G125), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n464), .B1(new_n465), .B2(KEYINPUT67), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G137), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n465), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n470), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(G112), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G2105), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n483), .B1(new_n471), .B2(new_n473), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT68), .ZN(new_n486));
  AOI211_X1 g061(.A(new_n482), .B(new_n486), .C1(G136), .C2(new_n474), .ZN(G162));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n483), .A2(G114), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n492), .A2(new_n494), .A3(KEYINPUT69), .A4(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  AND3_X1   g071(.A1(new_n472), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n497));
  AOI21_X1  g072(.A(KEYINPUT3), .B1(new_n472), .B2(G2104), .ZN(new_n498));
  OAI211_X1 g073(.A(G126), .B(G2105), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n471), .A2(new_n473), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n483), .A2(G138), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n500), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n500), .A2(new_n483), .A3(G138), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n505), .B1(new_n466), .B2(new_n467), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n496), .B(new_n499), .C1(new_n504), .C2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  NAND2_X1  g083(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT70), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n517), .B1(new_n515), .B2(KEYINPUT71), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT70), .A2(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT6), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g096(.A(new_n517), .B(KEYINPUT6), .C1(new_n515), .C2(KEYINPUT71), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(G543), .A3(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G50), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n521), .A2(new_n513), .A3(G88), .A4(new_n522), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n516), .A2(new_n525), .A3(new_n526), .A4(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G50), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n527), .B1(new_n523), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n514), .A2(new_n515), .ZN(new_n531));
  OAI21_X1  g106(.A(KEYINPUT73), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n528), .A2(new_n532), .ZN(G166));
  NAND2_X1  g108(.A1(new_n524), .A2(G51), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n521), .A2(new_n513), .A3(new_n522), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G89), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n539));
  AND2_X1   g114(.A1(G63), .A2(G651), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n538), .A2(new_n539), .B1(new_n513), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n534), .A2(new_n536), .A3(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  AOI22_X1  g118(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n515), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n524), .A2(G52), .ZN(new_n546));
  XNOR2_X1  g121(.A(KEYINPUT74), .B(G90), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n535), .A2(new_n547), .ZN(new_n548));
  AND3_X1   g123(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(G171));
  NAND4_X1  g124(.A1(new_n521), .A2(new_n513), .A3(G81), .A4(new_n522), .ZN(new_n550));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n523), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n513), .A2(G56), .ZN(new_n553));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n515), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(new_n561));
  XOR2_X1   g136(.A(new_n561), .B(KEYINPUT75), .Z(G188));
  NAND2_X1  g137(.A1(new_n535), .A2(G91), .ZN(new_n563));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n523), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NOR3_X1   g142(.A1(new_n523), .A2(KEYINPUT9), .A3(new_n564), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n563), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n513), .A2(G65), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n515), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT76), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G299));
  NAND3_X1  g150(.A1(new_n545), .A2(new_n548), .A3(new_n546), .ZN(G301));
  AND2_X1   g151(.A1(new_n528), .A2(new_n532), .ZN(G303));
  NAND4_X1  g152(.A1(new_n521), .A2(new_n513), .A3(G87), .A4(new_n522), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n521), .A2(G49), .A3(G543), .A4(new_n522), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n582), .B1(new_n511), .B2(new_n512), .ZN(new_n583));
  AND2_X1   g158(.A1(G73), .A2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n521), .A2(new_n513), .A3(G86), .A4(new_n522), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n521), .A2(G48), .A3(G543), .A4(new_n522), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(G305));
  AOI22_X1  g163(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(new_n515), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n524), .A2(G47), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n535), .A2(G85), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n521), .A2(new_n513), .A3(G92), .A4(new_n522), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n595), .B(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(new_n515), .ZN(new_n599));
  INV_X1    g174(.A(G54), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n523), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT77), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n594), .B1(new_n604), .B2(G868), .ZN(G284));
  XOR2_X1   g180(.A(G284), .B(KEYINPUT78), .Z(G321));
  NAND2_X1  g181(.A1(G286), .A2(G868), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(new_n574), .B2(G868), .ZN(G297));
  OAI21_X1  g183(.A(new_n607), .B1(new_n574), .B2(G868), .ZN(G280));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n604), .B1(new_n610), .B2(G860), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(KEYINPUT79), .Z(G148));
  NAND2_X1  g187(.A1(new_n604), .A2(new_n610), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G868), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g191(.A1(new_n466), .A2(new_n467), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(new_n476), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2100), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n474), .A2(G135), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT80), .Z(new_n623));
  NAND2_X1  g198(.A1(new_n484), .A2(G123), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n483), .A2(G111), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n627), .A2(G2096), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(G2096), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n621), .A2(new_n628), .A3(new_n629), .ZN(G156));
  INV_X1    g205(.A(KEYINPUT14), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(new_n634), .B2(new_n633), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2451), .B(G2454), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n636), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(G14), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT81), .ZN(G401));
  XNOR2_X1  g221(.A(G2072), .B(G2078), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT17), .Z(new_n648));
  XNOR2_X1  g223(.A(G2067), .B(G2678), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n649), .B2(new_n647), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT82), .Z(new_n656));
  NAND3_X1  g231(.A1(new_n652), .A2(new_n649), .A3(new_n647), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT18), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n653), .A2(new_n649), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n658), .B1(new_n648), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2096), .B(G2100), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1971), .B(G1976), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  AND2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT20), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n666), .A2(new_n667), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n665), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n665), .B2(new_n671), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1991), .B(G1996), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1981), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G229));
  INV_X1    g255(.A(G16), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G22), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(G166), .B2(new_n681), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n683), .A2(G1971), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(G1971), .ZN(new_n685));
  NOR2_X1   g260(.A1(G6), .A2(G16), .ZN(new_n686));
  INV_X1    g261(.A(G305), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n686), .B1(new_n687), .B2(G16), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT32), .B(G1981), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n681), .A2(G23), .ZN(new_n691));
  INV_X1    g266(.A(G288), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(new_n681), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT33), .B(G1976), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT83), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n693), .B(new_n695), .ZN(new_n696));
  NAND4_X1  g271(.A1(new_n684), .A2(new_n685), .A3(new_n690), .A4(new_n696), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n697), .A2(KEYINPUT34), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(KEYINPUT34), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n474), .A2(G131), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n484), .A2(G119), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n483), .A2(G107), .ZN(new_n702));
  OAI21_X1  g277(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n700), .B(new_n701), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  MUX2_X1   g279(.A(G25), .B(new_n704), .S(G29), .Z(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT35), .B(G1991), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n705), .B(new_n706), .Z(new_n707));
  INV_X1    g282(.A(G1986), .ZN(new_n708));
  AND3_X1   g283(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n709), .A2(new_n681), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n681), .B2(G24), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n707), .B1(new_n708), .B2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n708), .B2(new_n711), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n698), .A2(new_n699), .A3(new_n713), .ZN(new_n714));
  OR2_X1    g289(.A1(KEYINPUT84), .A2(KEYINPUT36), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(KEYINPUT84), .A2(KEYINPUT36), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT85), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n716), .B(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(G29), .A2(G32), .ZN(new_n720));
  NAND3_X1  g295(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT26), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n723), .A2(new_n724), .B1(G105), .B2(new_n476), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n474), .A2(G141), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n484), .A2(G129), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT92), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n732), .A2(KEYINPUT93), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT93), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n730), .B2(new_n731), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n720), .B1(new_n736), .B2(G29), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT27), .B(G1996), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n737), .A2(new_n739), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n681), .A2(G20), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT97), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT23), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n574), .B2(new_n681), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G1956), .ZN(new_n746));
  NOR3_X1   g321(.A1(new_n740), .A2(new_n741), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n681), .A2(G4), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n604), .B2(new_n681), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT86), .B(G1348), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G29), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G35), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT96), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G162), .B2(new_n752), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT29), .ZN(new_n756));
  INV_X1    g331(.A(G2090), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT31), .B(G11), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT94), .B(G28), .Z(new_n760));
  NOR2_X1   g335(.A1(new_n760), .A2(KEYINPUT30), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(KEYINPUT30), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(new_n752), .ZN(new_n763));
  OAI221_X1 g338(.A(new_n759), .B1(new_n761), .B2(new_n763), .C1(new_n627), .C2(new_n752), .ZN(new_n764));
  INV_X1    g339(.A(G2084), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT24), .B(G34), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n766), .A2(G29), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n478), .B2(G29), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n764), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n681), .A2(G21), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G168), .B2(new_n681), .ZN(new_n771));
  INV_X1    g346(.A(G1966), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n681), .A2(G5), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G171), .B2(new_n681), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n769), .B(new_n773), .C1(G1961), .C2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n752), .A2(G26), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT28), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n474), .A2(G140), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n484), .A2(G128), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n483), .A2(G116), .ZN(new_n781));
  OAI21_X1  g356(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n779), .B(new_n780), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n778), .B1(new_n783), .B2(G29), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT90), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT89), .B(G2067), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n752), .A2(G33), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n483), .A2(G103), .A3(G2104), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT25), .Z(new_n790));
  NAND2_X1  g365(.A1(new_n474), .A2(G139), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n617), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n793), .A2(new_n483), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n788), .B1(new_n795), .B2(new_n752), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n796), .A2(G2072), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT91), .ZN(new_n798));
  INV_X1    g373(.A(G19), .ZN(new_n799));
  OR3_X1    g374(.A1(new_n799), .A2(KEYINPUT87), .A3(G16), .ZN(new_n800));
  OAI21_X1  g375(.A(KEYINPUT87), .B1(new_n799), .B2(G16), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n800), .B(new_n801), .C1(new_n556), .C2(new_n681), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT88), .B(G1341), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(G164), .A2(G29), .ZN(new_n805));
  OR2_X1    g380(.A1(G27), .A2(G29), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n808), .A2(G2078), .B1(new_n796), .B2(G2072), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n768), .A2(new_n765), .ZN(new_n810));
  INV_X1    g385(.A(G2078), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n810), .B1(new_n807), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n804), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  NOR4_X1   g388(.A1(new_n776), .A2(new_n787), .A3(new_n798), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n775), .A2(G1961), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT95), .Z(new_n816));
  AND4_X1   g391(.A1(new_n751), .A2(new_n758), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n719), .A2(new_n747), .A3(new_n817), .ZN(G150));
  INV_X1    g393(.A(G150), .ZN(G311));
  INV_X1    g394(.A(new_n555), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n524), .A2(G43), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT99), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n820), .A2(new_n821), .A3(new_n822), .A4(new_n550), .ZN(new_n823));
  OAI21_X1  g398(.A(KEYINPUT99), .B1(new_n552), .B2(new_n555), .ZN(new_n824));
  INV_X1    g399(.A(G67), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(new_n511), .B2(new_n512), .ZN(new_n826));
  AND2_X1   g401(.A1(G80), .A2(G543), .ZN(new_n827));
  OAI21_X1  g402(.A(G651), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  XOR2_X1   g403(.A(KEYINPUT98), .B(G93), .Z(new_n829));
  NAND4_X1  g404(.A1(new_n829), .A2(new_n521), .A3(new_n513), .A4(new_n522), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n521), .A2(G55), .A3(G543), .A4(new_n522), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n828), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n823), .A2(new_n824), .A3(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n832), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n556), .A2(new_n822), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT38), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n604), .A2(G559), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n839), .A2(KEYINPUT39), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n839), .A2(KEYINPUT39), .ZN(new_n841));
  NOR3_X1   g416(.A1(new_n840), .A2(new_n841), .A3(G860), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n832), .A2(G860), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT37), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n842), .A2(new_n844), .ZN(G145));
  NAND2_X1  g420(.A1(new_n474), .A2(G142), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n484), .A2(G130), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n483), .A2(G118), .ZN(new_n848));
  OAI21_X1  g423(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n846), .B(new_n847), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n619), .B(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n704), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n795), .B1(new_n733), .B2(new_n735), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n507), .B(new_n783), .Z(new_n855));
  OR2_X1    g430(.A1(new_n732), .A2(new_n795), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n855), .B1(new_n854), .B2(new_n856), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n853), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n854), .A2(new_n856), .ZN(new_n861));
  INV_X1    g436(.A(new_n855), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n863), .A2(new_n852), .A3(new_n857), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT100), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n860), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n627), .B(new_n478), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(G162), .Z(new_n868));
  AOI21_X1  g443(.A(G37), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n870), .A2(new_n865), .A3(new_n864), .A4(new_n860), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(KEYINPUT101), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT101), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n869), .A2(new_n874), .A3(new_n871), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n873), .A2(KEYINPUT40), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(KEYINPUT40), .B1(new_n873), .B2(new_n875), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(G395));
  INV_X1    g453(.A(G868), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n832), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n881));
  NAND2_X1  g456(.A1(G303), .A2(G305), .ZN(new_n882));
  NAND2_X1  g457(.A1(G166), .A2(new_n687), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n709), .A2(new_n692), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT103), .ZN(new_n886));
  NAND2_X1  g461(.A1(G290), .A2(G288), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n887), .ZN(new_n891));
  NOR2_X1   g466(.A1(G290), .A2(G288), .ZN(new_n892));
  OAI21_X1  g467(.A(KEYINPUT103), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n893), .A2(new_n882), .A3(new_n883), .A4(new_n888), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n881), .B1(new_n895), .B2(KEYINPUT104), .ZN(new_n896));
  AOI21_X1  g471(.A(KEYINPUT104), .B1(new_n895), .B2(KEYINPUT105), .ZN(new_n897));
  MUX2_X1   g472(.A(new_n896), .B(new_n881), .S(new_n897), .Z(new_n898));
  XNOR2_X1  g473(.A(new_n613), .B(new_n836), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n597), .A2(new_n602), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(new_n573), .B2(new_n569), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n565), .B(new_n566), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT76), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n572), .B(new_n903), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n603), .A2(new_n902), .A3(new_n904), .A4(new_n563), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n901), .A2(new_n905), .A3(KEYINPUT102), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n900), .B(new_n907), .C1(new_n573), .C2(new_n569), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n906), .A2(KEYINPUT41), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT41), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n901), .A2(new_n910), .A3(new_n905), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n899), .A2(new_n912), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n906), .A2(new_n908), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n913), .B1(new_n914), .B2(new_n899), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n898), .B(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n880), .B1(new_n916), .B2(new_n879), .ZN(G295));
  OAI21_X1  g492(.A(new_n880), .B1(new_n916), .B2(new_n879), .ZN(G331));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT110), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n921));
  NAND2_X1  g496(.A1(G171), .A2(G168), .ZN(new_n922));
  NAND2_X1  g497(.A1(G301), .A2(G286), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n836), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n922), .A2(new_n833), .A3(new_n923), .A4(new_n835), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n921), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n926), .A2(new_n921), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n911), .B(new_n909), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n924), .A2(new_n836), .ZN(new_n931));
  AOI22_X1  g506(.A1(new_n922), .A2(new_n923), .B1(new_n833), .B2(new_n835), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n914), .A2(new_n930), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n895), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n906), .A2(new_n925), .A3(new_n908), .A4(new_n926), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT107), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n929), .A2(new_n934), .A3(new_n935), .A4(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G37), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n890), .A2(new_n894), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n941), .B1(new_n890), .B2(new_n894), .ZN(new_n943));
  OR2_X1    g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n906), .A2(new_n908), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n910), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n910), .B1(new_n901), .B2(new_n905), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n947), .B1(new_n926), .B2(new_n925), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n927), .A2(new_n945), .A3(new_n928), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n949), .B1(new_n950), .B2(KEYINPUT109), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT106), .B1(new_n931), .B2(new_n932), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n926), .A2(new_n921), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(new_n914), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n944), .B1(new_n951), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n940), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n942), .A2(new_n943), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n936), .B(new_n930), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n960), .B1(new_n929), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n938), .A2(new_n939), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT43), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n920), .B1(new_n959), .B2(new_n964), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n954), .A2(new_n955), .B1(new_n946), .B2(new_n948), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n950), .A2(KEYINPUT109), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n960), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n968), .A2(new_n963), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT110), .B1(new_n969), .B2(new_n958), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n919), .B1(new_n965), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n962), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT43), .B1(new_n972), .B2(new_n940), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n968), .A2(new_n958), .A3(new_n963), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT44), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n971), .A2(new_n975), .ZN(G397));
  INV_X1    g551(.A(G1384), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n501), .A2(new_n503), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n506), .B1(new_n978), .B2(KEYINPUT4), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n496), .A2(new_n499), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n977), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n470), .A2(new_n475), .A3(G40), .A4(new_n477), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G1996), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT111), .ZN(new_n988));
  XOR2_X1   g563(.A(new_n988), .B(KEYINPUT46), .Z(new_n989));
  XNOR2_X1  g564(.A(new_n985), .B(KEYINPUT112), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n783), .B(G2067), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n990), .B1(new_n732), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT125), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n992), .B(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n989), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT47), .ZN(new_n996));
  INV_X1    g571(.A(new_n991), .ZN(new_n997));
  INV_X1    g572(.A(new_n732), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n997), .B1(new_n998), .B2(new_n986), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n988), .A2(new_n736), .B1(new_n999), .B2(new_n990), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n704), .A2(new_n706), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n783), .A2(G2067), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n990), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n985), .A2(new_n708), .A3(new_n709), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1005), .B(KEYINPUT127), .ZN(new_n1006));
  XNOR2_X1  g581(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n704), .A2(new_n706), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n990), .B1(new_n1009), .B2(new_n1001), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1008), .A2(new_n1000), .A3(new_n1010), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n996), .A2(new_n1004), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1971), .ZN(new_n1013));
  INV_X1    g588(.A(new_n984), .ZN(new_n1014));
  AOI22_X1  g589(.A1(G126), .A2(new_n484), .B1(new_n491), .B2(new_n495), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n617), .A2(new_n500), .A3(new_n503), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n502), .B1(new_n471), .B2(new_n473), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1016), .B1(new_n1017), .B2(new_n500), .ZN(new_n1018));
  AOI21_X1  g593(.A(G1384), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1014), .B1(new_n1019), .B2(KEYINPUT45), .ZN(new_n1020));
  AOI211_X1 g595(.A(new_n982), .B(G1384), .C1(new_n1015), .C2(new_n1018), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1013), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n981), .A2(KEYINPUT50), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1023), .A2(new_n1025), .A3(new_n757), .A4(new_n1014), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1022), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(G8), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n528), .A2(new_n532), .A3(G8), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n528), .A2(new_n532), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1028), .A2(KEYINPUT115), .A3(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n578), .A2(new_n579), .A3(new_n580), .A4(G1976), .ZN(new_n1035));
  OAI211_X1 g610(.A(G8), .B(new_n1035), .C1(new_n981), .C2(new_n984), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT52), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(new_n692), .B2(G1976), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1037), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1040));
  XOR2_X1   g615(.A(KEYINPUT113), .B(G1981), .Z(new_n1041));
  NAND4_X1  g616(.A1(new_n585), .A2(new_n586), .A3(new_n587), .A4(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G1981), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1042), .B1(new_n687), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT49), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT114), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1044), .A2(new_n1048), .A3(new_n1045), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1014), .A2(new_n1019), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(G8), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1040), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n1056));
  INV_X1    g631(.A(G8), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1057), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1056), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1034), .A2(new_n1055), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1014), .B1(new_n1019), .B2(new_n1024), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n981), .A2(KEYINPUT50), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT117), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G1961), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1023), .A2(new_n1025), .A3(new_n1067), .A4(new_n1014), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1065), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n984), .B1(new_n981), .B2(new_n982), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1019), .A2(KEYINPUT45), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n811), .A3(new_n1071), .ZN(new_n1072));
  XOR2_X1   g647(.A(KEYINPUT122), .B(KEYINPUT53), .Z(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT45), .B1(new_n507), .B2(new_n977), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1075), .B1(new_n1076), .B2(new_n984), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1014), .B(KEYINPUT116), .C1(new_n1019), .C2(KEYINPUT45), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n811), .A2(KEYINPUT53), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1077), .A2(new_n1071), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1069), .A2(new_n1074), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G171), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1062), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n1084));
  NAND3_X1  g659(.A1(G286), .A2(new_n1084), .A3(G8), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1084), .B1(G286), .B2(G8), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT51), .B1(new_n1088), .B2(KEYINPUT121), .ZN(new_n1089));
  NOR3_X1   g664(.A1(new_n1063), .A2(new_n1064), .A3(G2084), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1077), .A2(new_n1071), .A3(new_n1078), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1090), .B1(new_n1091), .B2(new_n772), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1089), .B(new_n1088), .C1(new_n1092), .C2(new_n1057), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT62), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1087), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n1085), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1078), .A2(new_n1071), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT116), .B1(new_n983), .B2(new_n1014), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n772), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1090), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1096), .B1(new_n1101), .B2(G8), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT51), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1103), .B1(new_n1096), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n1092), .B2(new_n1088), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1093), .B(new_n1094), .C1(new_n1102), .C2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1021), .B1(new_n1070), .B2(KEYINPUT116), .ZN(new_n1109));
  AOI21_X1  g684(.A(G1966), .B1(new_n1109), .B2(new_n1077), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1096), .B1(new_n1110), .B2(new_n1090), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1057), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1111), .B(new_n1105), .C1(new_n1112), .C2(new_n1096), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1094), .B1(new_n1113), .B2(new_n1093), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1083), .B1(new_n1108), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1055), .A2(new_n1059), .A3(new_n1058), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1050), .A2(new_n1054), .ZN(new_n1117));
  NOR2_X1   g692(.A1(G288), .A2(G1976), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1117), .A2(new_n1118), .B1(new_n687), .B2(new_n1041), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1116), .B1(new_n1119), .B2(new_n1053), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT63), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1112), .A2(G168), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1121), .B1(new_n1062), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1122), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1121), .B1(new_n1028), .B2(new_n1033), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1124), .A2(new_n1125), .A3(new_n1061), .A4(new_n1055), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1120), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(G1956), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT56), .B(G2072), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1070), .A2(new_n1071), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT57), .B1(new_n569), .B2(new_n573), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT57), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n902), .A2(new_n904), .A3(new_n1134), .A4(new_n563), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1132), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n900), .ZN(new_n1139));
  INV_X1    g714(.A(G1348), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1065), .A2(new_n1140), .A3(new_n1068), .ZN(new_n1141));
  OR2_X1    g716(.A1(new_n1052), .A2(G2067), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1136), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1132), .ZN(new_n1145));
  OAI22_X1  g720(.A1(new_n1139), .A2(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1129), .A2(new_n1131), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1147), .B1(new_n1137), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT59), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT118), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1070), .A2(new_n986), .A3(new_n1071), .ZN(new_n1152));
  XOR2_X1   g727(.A(KEYINPUT58), .B(G1341), .Z(new_n1153));
  NAND2_X1  g728(.A1(new_n1052), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1151), .B1(new_n1155), .B2(new_n556), .ZN(new_n1156));
  INV_X1    g731(.A(new_n556), .ZN(new_n1157));
  XOR2_X1   g732(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n1158));
  AOI211_X1 g733(.A(new_n1157), .B(new_n1158), .C1(new_n1152), .C2(new_n1154), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1141), .A2(KEYINPUT60), .A3(new_n603), .A4(new_n1142), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1149), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1141), .A2(KEYINPUT60), .A3(new_n1142), .ZN(new_n1163));
  AOI21_X1  g738(.A(KEYINPUT60), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1163), .A2(new_n1164), .A3(new_n603), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT119), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1138), .B1(new_n1167), .B2(new_n1148), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1145), .A2(KEYINPUT119), .A3(new_n1144), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1168), .A2(KEYINPUT61), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1146), .B1(new_n1166), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1093), .B1(new_n1102), .B2(new_n1106), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1070), .A2(new_n1071), .A3(new_n1079), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT123), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1070), .A2(KEYINPUT123), .A3(new_n1071), .A4(new_n1079), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1177), .A2(G301), .A3(new_n1069), .A4(new_n1074), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT54), .B1(new_n1082), .B2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1172), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1177), .A2(new_n1069), .A3(new_n1074), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(G171), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1069), .A2(new_n1074), .A3(G301), .A4(new_n1080), .ZN(new_n1183));
  AND2_X1   g758(.A1(new_n1183), .A2(KEYINPUT54), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1062), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1180), .A2(new_n1185), .ZN(new_n1186));
  OAI211_X1 g761(.A(new_n1115), .B(new_n1127), .C1(new_n1171), .C2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1000), .A2(new_n1010), .ZN(new_n1188));
  XNOR2_X1  g763(.A(G290), .B(G1986), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1188), .B1(new_n985), .B2(new_n1189), .ZN(new_n1190));
  AND3_X1   g765(.A1(new_n1187), .A2(KEYINPUT124), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g766(.A(KEYINPUT124), .B1(new_n1187), .B2(new_n1190), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1012), .B1(new_n1191), .B2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g768(.A1(new_n965), .A2(new_n970), .ZN(new_n1195));
  NOR2_X1   g769(.A1(G227), .A2(new_n461), .ZN(new_n1196));
  NAND2_X1  g770(.A1(new_n1196), .A2(new_n645), .ZN(new_n1197));
  NOR2_X1   g771(.A1(G229), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g772(.A(new_n875), .ZN(new_n1199));
  AOI21_X1  g773(.A(new_n874), .B1(new_n869), .B2(new_n871), .ZN(new_n1200));
  OAI21_X1  g774(.A(new_n1198), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g775(.A1(new_n1195), .A2(new_n1201), .ZN(G308));
  OAI221_X1 g776(.A(new_n1198), .B1(new_n1199), .B2(new_n1200), .C1(new_n965), .C2(new_n970), .ZN(G225));
endmodule


