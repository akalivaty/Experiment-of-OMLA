//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0 1 0 0 0 0 1 0 1 0 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967,
    new_n968, new_n969;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  INV_X1    g001(.A(G211gat), .ZN(new_n203));
  INV_X1    g002(.A(G218gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n202), .B1(KEYINPUT22), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G211gat), .B(G218gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G141gat), .B(G148gat), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n209), .B(new_n211), .C1(new_n212), .C2(KEYINPUT2), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(KEYINPUT73), .ZN(new_n214));
  INV_X1    g013(.A(G141gat), .ZN(new_n215));
  INV_X1    g014(.A(G148gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT73), .ZN(new_n218));
  NAND2_X1  g017(.A1(G141gat), .A2(G148gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT74), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n209), .B1(new_n211), .B2(KEYINPUT2), .ZN(new_n223));
  AND3_X1   g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n222), .B1(new_n221), .B2(new_n223), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n213), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  XOR2_X1   g025(.A(KEYINPUT75), .B(KEYINPUT3), .Z(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n208), .B1(new_n229), .B2(KEYINPUT29), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n227), .B1(new_n208), .B2(KEYINPUT29), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n232), .A2(new_n226), .ZN(new_n233));
  INV_X1    g032(.A(G228gat), .ZN(new_n234));
  INV_X1    g033(.A(G233gat), .ZN(new_n235));
  OAI22_X1  g034(.A1(new_n231), .A2(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n230), .A2(KEYINPUT80), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n234), .A2(new_n235), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n208), .A2(KEYINPUT29), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n239), .A2(KEYINPUT79), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(new_n239), .B2(KEYINPUT79), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n226), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n237), .A2(new_n238), .A3(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n230), .A2(KEYINPUT80), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n236), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G22gat), .ZN(new_n247));
  INV_X1    g046(.A(G22gat), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n236), .B(new_n248), .C1(new_n244), .C2(new_n245), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(G78gat), .ZN(new_n251));
  INV_X1    g050(.A(G78gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n247), .A2(new_n252), .A3(new_n249), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT31), .B(G50gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(KEYINPUT81), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(G106gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n251), .A2(new_n253), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n256), .ZN(new_n258));
  INV_X1    g057(.A(new_n253), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n252), .B1(new_n247), .B2(new_n249), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(G169gat), .A2(G176gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT23), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(G169gat), .ZN(new_n265));
  INV_X1    g064(.A(G176gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT24), .ZN(new_n268));
  INV_X1    g067(.A(G183gat), .ZN(new_n269));
  INV_X1    g068(.A(G190gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n267), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n269), .A2(new_n270), .ZN(new_n273));
  NAND2_X1  g072(.A1(G183gat), .A2(G190gat), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(KEYINPUT24), .A3(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n264), .A2(new_n272), .A3(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  AND2_X1   g077(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n279));
  OR2_X1    g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G127gat), .B(G134gat), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT66), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G113gat), .B(G120gat), .ZN(new_n284));
  OR2_X1    g083(.A1(new_n284), .A2(KEYINPUT1), .ZN(new_n285));
  AND2_X1   g084(.A1(new_n281), .A2(new_n282), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n283), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT1), .B1(new_n284), .B2(KEYINPUT67), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT67), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n281), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n288), .B1(new_n290), .B2(new_n284), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(KEYINPUT27), .B(G183gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(KEYINPUT65), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n295), .A2(KEYINPUT28), .A3(new_n270), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n294), .A2(new_n270), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n297), .A2(KEYINPUT28), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NOR3_X1   g098(.A1(new_n267), .A2(KEYINPUT26), .A3(new_n262), .ZN(new_n300));
  AOI211_X1 g099(.A(new_n271), .B(new_n300), .C1(KEYINPUT26), .C2(new_n262), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n280), .A2(new_n293), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n302), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n278), .A2(new_n279), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n292), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G227gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n307), .A2(new_n235), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n303), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  XOR2_X1   g108(.A(G71gat), .B(G99gat), .Z(new_n310));
  XNOR2_X1  g109(.A(G15gat), .B(G43gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n310), .B(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT33), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n309), .A2(KEYINPUT32), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT68), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n314), .B(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n309), .A2(KEYINPUT32), .ZN(new_n317));
  INV_X1    g116(.A(new_n309), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n317), .B(new_n312), .C1(new_n318), .C2(KEYINPUT33), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n306), .ZN(new_n320));
  INV_X1    g119(.A(new_n308), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n322), .A2(KEYINPUT34), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(KEYINPUT34), .ZN(new_n325));
  AND2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n316), .B(new_n319), .C1(KEYINPUT69), .C2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n316), .A2(new_n319), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n324), .A2(new_n325), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT69), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  AND4_X1   g130(.A1(new_n257), .A2(new_n261), .A3(new_n327), .A4(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G1gat), .B(G29gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n333), .B(KEYINPUT0), .ZN(new_n334));
  XNOR2_X1  g133(.A(G57gat), .B(G85gat), .ZN(new_n335));
  XOR2_X1   g134(.A(new_n334), .B(new_n335), .Z(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n226), .A2(new_n293), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT77), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n292), .B(new_n213), .C1(new_n225), .C2(new_n224), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(G225gat), .A2(G233gat), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n226), .A2(KEYINPUT77), .A3(new_n293), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT5), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT78), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT78), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n345), .A2(new_n348), .A3(KEYINPUT5), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n292), .B1(new_n226), .B2(KEYINPUT3), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n350), .B1(new_n226), .B2(new_n228), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n342), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT4), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n340), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(KEYINPUT76), .B(KEYINPUT4), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n355), .B1(new_n340), .B2(new_n356), .ZN(new_n357));
  AOI22_X1  g156(.A1(new_n347), .A2(new_n349), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n340), .A2(new_n354), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n359), .B1(new_n340), .B2(new_n356), .ZN(new_n360));
  NOR3_X1   g159(.A1(new_n352), .A2(new_n360), .A3(KEYINPUT5), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n337), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT6), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n353), .A2(new_n357), .ZN(new_n364));
  AND3_X1   g163(.A1(new_n345), .A2(new_n348), .A3(KEYINPUT5), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n348), .B1(new_n345), .B2(KEYINPUT5), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n361), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n367), .A2(new_n336), .A3(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n362), .A2(new_n363), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n336), .B1(new_n367), .B2(new_n368), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT6), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  AND2_X1   g172(.A1(G226gat), .A2(G233gat), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n280), .A2(new_n374), .A3(new_n302), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n280), .A2(KEYINPUT71), .A3(new_n302), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT71), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n377), .B1(new_n304), .B2(new_n305), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n374), .A2(KEYINPUT29), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n375), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n381), .A2(new_n208), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n376), .A2(new_n378), .A3(new_n374), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n380), .B1(new_n304), .B2(new_n305), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n208), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  XOR2_X1   g185(.A(G8gat), .B(G36gat), .Z(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(KEYINPUT72), .ZN(new_n388));
  XNOR2_X1  g187(.A(G64gat), .B(G92gat), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n388), .B(new_n389), .Z(new_n390));
  OR4_X1    g189(.A1(KEYINPUT30), .A2(new_n382), .A3(new_n386), .A4(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n208), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n379), .A2(new_n380), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n392), .B1(new_n393), .B2(new_n375), .ZN(new_n394));
  INV_X1    g193(.A(new_n390), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n394), .A2(new_n385), .A3(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n390), .B1(new_n382), .B2(new_n386), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(new_n397), .A3(KEYINPUT30), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n391), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n373), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n332), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT35), .ZN(new_n403));
  INV_X1    g202(.A(new_n399), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n328), .A2(new_n329), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n326), .A2(new_n316), .A3(new_n319), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NOR3_X1   g206(.A1(new_n404), .A2(new_n407), .A3(KEYINPUT35), .ZN(new_n408));
  OR2_X1    g207(.A1(new_n370), .A2(KEYINPUT82), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n370), .A2(KEYINPUT82), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n372), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n261), .A2(new_n257), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n408), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n403), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n351), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n343), .B1(new_n416), .B2(new_n360), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n341), .A2(new_n344), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n417), .B(KEYINPUT39), .C1(new_n343), .C2(new_n418), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n419), .B(new_n336), .C1(KEYINPUT39), .C2(new_n417), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT40), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n422), .A2(new_n371), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n404), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT37), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n425), .B1(new_n394), .B2(new_n385), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n385), .B(new_n425), .C1(new_n381), .C2(new_n208), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n390), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT38), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n396), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n208), .B1(new_n383), .B2(new_n384), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT83), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n431), .A2(new_n432), .B1(new_n381), .B2(new_n208), .ZN(new_n433));
  OR2_X1    g232(.A1(new_n431), .A2(new_n432), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n425), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n435), .A2(KEYINPUT38), .A3(new_n428), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n430), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n424), .B(new_n413), .C1(new_n411), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n412), .A2(new_n400), .ZN(new_n439));
  XNOR2_X1  g238(.A(KEYINPUT70), .B(KEYINPUT36), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n407), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n327), .A2(new_n331), .A3(KEYINPUT36), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n438), .A2(new_n439), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n415), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(G15gat), .B(G22gat), .ZN(new_n446));
  OR2_X1    g245(.A1(new_n446), .A2(G1gat), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT87), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT16), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n446), .B1(new_n449), .B2(G1gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n448), .A2(new_n451), .A3(G8gat), .ZN(new_n452));
  INV_X1    g251(.A(G8gat), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n447), .B(new_n450), .C1(KEYINPUT87), .C2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT86), .ZN(new_n457));
  XNOR2_X1  g256(.A(KEYINPUT14), .B(G29gat), .ZN(new_n458));
  INV_X1    g257(.A(G36gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(G29gat), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n462));
  INV_X1    g261(.A(G43gat), .ZN(new_n463));
  INV_X1    g262(.A(G50gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(G43gat), .A2(G50gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n460), .A2(KEYINPUT15), .A3(new_n462), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n460), .A2(new_n462), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(KEYINPUT15), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT15), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n465), .A2(new_n471), .A3(new_n466), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n469), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n468), .B1(new_n473), .B2(KEYINPUT85), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT85), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n470), .A2(new_n472), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n475), .B1(new_n476), .B2(new_n469), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n457), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n473), .A2(KEYINPUT85), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n476), .A2(new_n475), .A3(new_n469), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n479), .A2(KEYINPUT86), .A3(new_n480), .A4(new_n468), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT17), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT17), .ZN(new_n483));
  INV_X1    g282(.A(new_n474), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n483), .B1(new_n484), .B2(new_n479), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n456), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(G229gat), .A2(G233gat), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT88), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n455), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n452), .A2(KEYINPUT88), .A3(new_n454), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n478), .A2(new_n489), .A3(new_n481), .A4(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n486), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  XOR2_X1   g291(.A(KEYINPUT89), .B(KEYINPUT18), .Z(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT91), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n486), .A2(KEYINPUT18), .A3(new_n487), .A4(new_n491), .ZN(new_n496));
  XOR2_X1   g295(.A(new_n487), .B(KEYINPUT13), .Z(new_n497));
  NAND2_X1  g296(.A1(new_n478), .A2(new_n481), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n489), .A2(new_n490), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n491), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n497), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G113gat), .B(G141gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G169gat), .B(G197gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n509), .B(KEYINPUT12), .Z(new_n510));
  INV_X1    g309(.A(KEYINPUT91), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n492), .A2(new_n511), .A3(new_n493), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n495), .A2(new_n504), .A3(new_n510), .A4(new_n512), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n492), .A2(KEYINPUT90), .A3(new_n493), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT90), .B1(new_n492), .B2(new_n493), .ZN(new_n515));
  NOR3_X1   g314(.A1(new_n514), .A2(new_n515), .A3(new_n503), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n513), .B1(new_n516), .B2(new_n510), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n445), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G120gat), .B(G148gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(G176gat), .B(G204gat), .ZN(new_n520));
  XOR2_X1   g319(.A(new_n519), .B(new_n520), .Z(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(G57gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n523), .A2(G64gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(G64gat), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n524), .B1(KEYINPUT92), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n526), .B1(KEYINPUT92), .B2(new_n525), .ZN(new_n527));
  NAND2_X1  g326(.A1(G71gat), .A2(G78gat), .ZN(new_n528));
  INV_X1    g327(.A(G71gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(new_n252), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT9), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n525), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT9), .B1(new_n534), .B2(new_n524), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n535), .A2(new_n528), .A3(new_n530), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G99gat), .B(G106gat), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT97), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G99gat), .A2(G106gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT95), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT95), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n544), .A2(G99gat), .A3(G106gat), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n545), .A3(KEYINPUT8), .ZN(new_n546));
  NOR2_X1   g345(.A1(G85gat), .A2(G92gat), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT96), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT96), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n546), .A2(new_n551), .A3(new_n548), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G85gat), .A2(G92gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT7), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n541), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT8), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n557), .B1(new_n542), .B2(KEYINPUT95), .ZN(new_n558));
  AOI211_X1 g357(.A(KEYINPUT96), .B(new_n547), .C1(new_n558), .C2(new_n545), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n551), .B1(new_n546), .B2(new_n548), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n541), .B(new_n555), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n538), .B1(new_n556), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT98), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n555), .B1(new_n559), .B2(new_n560), .ZN(new_n565));
  INV_X1    g364(.A(new_n541), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n567), .A2(new_n537), .A3(new_n561), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n563), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n561), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n570), .A2(KEYINPUT98), .A3(new_n538), .ZN(new_n571));
  AOI21_X1  g370(.A(KEYINPUT10), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT99), .ZN(new_n573));
  AND4_X1   g372(.A1(new_n573), .A2(new_n570), .A3(KEYINPUT10), .A4(new_n538), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n537), .B1(new_n567), .B2(new_n561), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n573), .B1(new_n575), .B2(KEYINPUT10), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G230gat), .A2(G233gat), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n569), .A2(new_n571), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n582), .A2(new_n579), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n522), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT10), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n564), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n586), .A2(new_n575), .ZN(new_n587));
  INV_X1    g386(.A(new_n571), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n585), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n576), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n575), .A2(new_n573), .A3(KEYINPUT10), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n589), .A2(KEYINPUT100), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT100), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n594), .B1(new_n572), .B2(new_n577), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n593), .A2(new_n595), .A3(new_n579), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n583), .A2(new_n522), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n584), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT101), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT101), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n584), .A2(new_n598), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n498), .ZN(new_n605));
  AND2_X1   g404(.A1(G232gat), .A2(G233gat), .ZN(new_n606));
  AOI22_X1  g405(.A1(new_n605), .A2(new_n570), .B1(KEYINPUT41), .B2(new_n606), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n561), .B(new_n567), .C1(new_n482), .C2(new_n485), .ZN(new_n608));
  XOR2_X1   g407(.A(G190gat), .B(G218gat), .Z(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n607), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n606), .A2(KEYINPUT41), .ZN(new_n613));
  XNOR2_X1  g412(.A(G134gat), .B(G162gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n610), .B1(new_n607), .B2(new_n608), .ZN(new_n617));
  OR3_X1    g416(.A1(new_n612), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n616), .B1(new_n612), .B2(new_n617), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT21), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n499), .B1(new_n622), .B2(new_n537), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n537), .A2(new_n622), .ZN(new_n624));
  XOR2_X1   g423(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n623), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G127gat), .B(G155gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT20), .ZN(new_n629));
  NAND2_X1  g428(.A1(G231gat), .A2(G233gat), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n630), .B(KEYINPUT93), .Z(new_n631));
  XNOR2_X1  g430(.A(new_n629), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G183gat), .B(G211gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n627), .B(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n621), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n604), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n518), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT102), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n373), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n370), .A2(KEYINPUT102), .A3(new_n372), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(G1gat), .ZN(G1324gat));
  INV_X1    g444(.A(new_n517), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n646), .B1(new_n415), .B2(new_n444), .ZN(new_n647));
  INV_X1    g446(.A(new_n637), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(new_n404), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(G8gat), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(KEYINPUT103), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT103), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n649), .A2(new_n652), .A3(G8gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g453(.A(KEYINPUT16), .B(G8gat), .Z(new_n655));
  NAND4_X1  g454(.A1(new_n647), .A2(new_n404), .A3(new_n648), .A4(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(KEYINPUT104), .B1(new_n654), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n656), .B(KEYINPUT42), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n660), .A2(new_n661), .A3(new_n651), .A4(new_n653), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(new_n662), .ZN(G1325gat));
  INV_X1    g462(.A(KEYINPUT106), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n443), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n441), .A2(KEYINPUT106), .A3(new_n442), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n638), .A2(G15gat), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n407), .ZN(new_n670));
  AOI21_X1  g469(.A(G15gat), .B1(new_n638), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n669), .B1(new_n673), .B2(new_n674), .ZN(G1326gat));
  NOR2_X1   g474(.A1(new_n518), .A2(new_n413), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n648), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT43), .B(G22gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  INV_X1    g478(.A(new_n635), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n603), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n621), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n518), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n683), .A2(new_n461), .A3(new_n643), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT45), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n621), .A2(KEYINPUT44), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n445), .A2(new_n686), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n603), .A2(new_n646), .A3(new_n680), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n412), .A2(new_n400), .A3(KEYINPUT107), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT107), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n439), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n438), .A2(new_n443), .A3(new_n689), .A4(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n620), .B1(new_n692), .B2(new_n415), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n687), .B(new_n688), .C1(new_n693), .C2(KEYINPUT44), .ZN(new_n694));
  OAI21_X1  g493(.A(G29gat), .B1(new_n694), .B2(new_n642), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n685), .A2(new_n695), .ZN(G1328gat));
  NOR2_X1   g495(.A1(new_n399), .A2(G36gat), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n683), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(KEYINPUT108), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n683), .A2(new_n700), .A3(new_n697), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT46), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(G36gat), .B1(new_n694), .B2(new_n399), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n699), .A2(KEYINPUT46), .A3(new_n701), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(G1329gat));
  OAI21_X1  g506(.A(G43gat), .B1(new_n694), .B2(new_n443), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n683), .A2(new_n463), .A3(new_n670), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n708), .A2(KEYINPUT47), .A3(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n709), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n694), .A2(new_n667), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n711), .B1(new_n712), .B2(G43gat), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n710), .B1(new_n713), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g513(.A(G50gat), .B1(new_n694), .B2(new_n413), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n676), .A2(new_n464), .A3(new_n621), .A4(new_n681), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT48), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n715), .A2(KEYINPUT48), .A3(new_n716), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(G1331gat));
  NAND3_X1  g520(.A1(new_n636), .A2(new_n646), .A3(new_n603), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n722), .B1(new_n692), .B2(new_n415), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n370), .A2(KEYINPUT102), .A3(new_n372), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT102), .B1(new_n370), .B2(new_n372), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n640), .A2(KEYINPUT109), .A3(new_n641), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n723), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(G57gat), .ZN(G1332gat));
  INV_X1    g530(.A(KEYINPUT110), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n692), .A2(new_n415), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n733), .B2(new_n722), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n723), .A2(KEYINPUT110), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n404), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n738));
  XOR2_X1   g537(.A(KEYINPUT49), .B(G64gat), .Z(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n737), .B2(new_n739), .ZN(G1333gat));
  NAND3_X1  g539(.A1(new_n734), .A2(new_n735), .A3(new_n668), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G71gat), .ZN(new_n742));
  AND3_X1   g541(.A1(new_n723), .A2(KEYINPUT111), .A3(new_n670), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT111), .B1(new_n723), .B2(new_n670), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n529), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT50), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n742), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n746), .B1(new_n742), .B2(new_n745), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(G1334gat));
  NAND2_X1  g548(.A1(new_n736), .A2(new_n412), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g550(.A1(new_n517), .A2(new_n680), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n693), .A2(KEYINPUT51), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT51), .B1(new_n693), .B2(new_n752), .ZN(new_n754));
  OR2_X1    g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n642), .A2(G85gat), .A3(new_n604), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT112), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n752), .A2(new_n603), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n687), .B(new_n759), .C1(new_n693), .C2(KEYINPUT44), .ZN(new_n760));
  OAI21_X1  g559(.A(G85gat), .B1(new_n760), .B2(new_n642), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n758), .A2(new_n761), .ZN(G1336gat));
  OAI21_X1  g561(.A(G92gat), .B1(new_n760), .B2(new_n399), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n399), .A2(G92gat), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n603), .B(new_n764), .C1(new_n753), .C2(new_n754), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(KEYINPUT52), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n763), .A2(new_n765), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(G1337gat));
  NOR2_X1   g569(.A1(new_n407), .A2(G99gat), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n755), .A2(new_n603), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(G99gat), .B1(new_n760), .B2(new_n667), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(G1338gat));
  XNOR2_X1  g573(.A(KEYINPUT113), .B(G106gat), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n775), .B1(new_n760), .B2(new_n413), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n413), .A2(G106gat), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n603), .B(new_n777), .C1(new_n753), .C2(new_n754), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g578(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n776), .A2(new_n778), .A3(new_n780), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(G1339gat));
  NOR2_X1   g583(.A1(new_n646), .A2(G113gat), .ZN(new_n785));
  XOR2_X1   g584(.A(new_n785), .B(KEYINPUT118), .Z(new_n786));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n787), .B(new_n579), .C1(new_n572), .C2(new_n577), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n788), .A2(KEYINPUT55), .A3(new_n522), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n787), .B1(new_n578), .B2(new_n580), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n789), .B1(new_n596), .B2(new_n790), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n596), .A2(new_n597), .ZN(new_n792));
  OAI21_X1  g591(.A(KEYINPUT115), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n589), .A2(new_n580), .A3(new_n592), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT54), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n589), .A2(new_n592), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n580), .B1(new_n797), .B2(new_n594), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n796), .B1(new_n798), .B2(new_n593), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n794), .B(new_n598), .C1(new_n799), .C2(new_n789), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n596), .A2(new_n790), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n788), .A2(new_n522), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n793), .A2(new_n800), .A3(new_n517), .A4(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n509), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n487), .B1(new_n486), .B2(new_n491), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n500), .A2(new_n501), .A3(new_n497), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n513), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n602), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n601), .B1(new_n584), .B2(new_n598), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n621), .B1(new_n806), .B2(new_n814), .ZN(new_n815));
  AND4_X1   g614(.A1(new_n513), .A2(new_n618), .A3(new_n619), .A4(new_n810), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n816), .A2(new_n800), .A3(new_n793), .A4(new_n805), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n635), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n648), .A2(new_n646), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n821), .A2(new_n729), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n822), .A2(KEYINPUT116), .A3(new_n332), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(new_n332), .A3(new_n729), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n404), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n827), .A2(KEYINPUT117), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n827), .A2(KEYINPUT117), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n786), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n412), .B1(new_n819), .B2(new_n820), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n831), .A2(new_n399), .A3(new_n670), .A4(new_n643), .ZN(new_n832));
  OAI21_X1  g631(.A(G113gat), .B1(new_n832), .B2(new_n646), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n830), .A2(new_n833), .ZN(G1340gat));
  NOR2_X1   g633(.A1(new_n604), .A2(G120gat), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n835), .B1(new_n828), .B2(new_n829), .ZN(new_n836));
  OAI21_X1  g635(.A(G120gat), .B1(new_n832), .B2(new_n604), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(G1341gat));
  INV_X1    g637(.A(G127gat), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n827), .A2(new_n839), .A3(new_n680), .ZN(new_n840));
  OAI21_X1  g639(.A(G127gat), .B1(new_n832), .B2(new_n635), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1342gat));
  NAND2_X1  g641(.A1(new_n823), .A2(new_n826), .ZN(new_n843));
  INV_X1    g642(.A(G134gat), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n399), .A2(new_n621), .ZN(new_n845));
  XOR2_X1   g644(.A(new_n845), .B(KEYINPUT119), .Z(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n843), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n848), .A2(KEYINPUT56), .ZN(new_n849));
  OAI21_X1  g648(.A(G134gat), .B1(new_n832), .B2(new_n620), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(KEYINPUT56), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(G1343gat));
  AOI21_X1  g651(.A(KEYINPUT122), .B1(new_n667), .B2(new_n412), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n441), .A2(KEYINPUT106), .A3(new_n442), .ZN(new_n854));
  AOI21_X1  g653(.A(KEYINPUT106), .B1(new_n441), .B2(new_n442), .ZN(new_n855));
  OAI211_X1 g654(.A(KEYINPUT122), .B(new_n412), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n646), .A2(G141gat), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n858), .A2(new_n822), .A3(new_n399), .A4(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n791), .A2(new_n792), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n517), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n803), .A2(KEYINPUT120), .ZN(new_n863));
  AOI21_X1  g662(.A(KEYINPUT55), .B1(new_n803), .B2(KEYINPUT120), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n814), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n620), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n680), .B1(new_n867), .B2(new_n817), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n637), .A2(new_n517), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n412), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(KEYINPUT57), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n413), .B1(new_n819), .B2(new_n820), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n643), .A2(new_n399), .A3(new_n443), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n871), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(new_n646), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n860), .B1(new_n877), .B2(new_n215), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n860), .A2(KEYINPUT121), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(KEYINPUT58), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n880), .B(new_n860), .C1(new_n877), .C2(new_n215), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1344gat));
  NOR2_X1   g683(.A1(new_n876), .A2(new_n604), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n885), .A2(KEYINPUT59), .A3(new_n216), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n872), .A2(new_n873), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n873), .B(new_n412), .C1(new_n868), .C2(new_n869), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n888), .A2(new_n603), .A3(new_n875), .A4(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n887), .B1(new_n890), .B2(G148gat), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n858), .A2(new_n822), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n399), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n603), .A2(new_n216), .ZN(new_n894));
  OAI22_X1  g693(.A1(new_n886), .A2(new_n891), .B1(new_n893), .B2(new_n894), .ZN(G1345gat));
  NAND4_X1  g694(.A1(new_n858), .A2(new_n822), .A3(new_n399), .A4(new_n680), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(G155gat), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n899), .B1(new_n896), .B2(new_n897), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n635), .A2(new_n899), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  OAI22_X1  g701(.A1(new_n898), .A2(new_n900), .B1(new_n876), .B2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT124), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI221_X1 g704(.A(KEYINPUT124), .B1(new_n876), .B2(new_n902), .C1(new_n898), .C2(new_n900), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(G1346gat));
  OAI21_X1  g706(.A(G162gat), .B1(new_n876), .B2(new_n620), .ZN(new_n908));
  INV_X1    g707(.A(G162gat), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n892), .A2(new_n909), .A3(new_n847), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(G1347gat));
  AOI21_X1  g710(.A(new_n643), .B1(new_n819), .B2(new_n820), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n332), .A2(new_n404), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(G169gat), .B1(new_n915), .B2(new_n517), .ZN(new_n916));
  AND4_X1   g715(.A1(new_n404), .A2(new_n727), .A3(new_n728), .A4(new_n670), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n806), .A2(new_n814), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n620), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n680), .B1(new_n919), .B2(new_n817), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n413), .B(new_n917), .C1(new_n920), .C2(new_n869), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT125), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT125), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n831), .A2(new_n924), .A3(new_n917), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n646), .A2(new_n265), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n916), .B1(new_n927), .B2(new_n928), .ZN(G1348gat));
  NAND3_X1  g728(.A1(new_n915), .A2(new_n266), .A3(new_n603), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n923), .A2(new_n926), .A3(new_n604), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n930), .B1(new_n931), .B2(new_n266), .ZN(G1349gat));
  NAND3_X1  g731(.A1(new_n915), .A2(new_n295), .A3(new_n680), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n923), .A2(new_n926), .A3(new_n635), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n933), .B1(new_n934), .B2(new_n269), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g735(.A1(new_n915), .A2(new_n270), .A3(new_n621), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n922), .A2(new_n621), .A3(new_n925), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n938), .A2(new_n939), .A3(G190gat), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n939), .B1(new_n938), .B2(G190gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI211_X1 g743(.A(KEYINPUT126), .B(new_n937), .C1(new_n940), .C2(new_n941), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1351gat));
  AND4_X1   g745(.A1(new_n404), .A2(new_n912), .A3(new_n412), .A4(new_n667), .ZN(new_n947));
  AOI21_X1  g746(.A(G197gat), .B1(new_n947), .B2(new_n517), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n668), .A2(new_n399), .A3(new_n729), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n888), .A2(new_n889), .A3(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n517), .A2(G197gat), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n948), .B1(new_n951), .B2(new_n952), .ZN(G1352gat));
  INV_X1    g752(.A(G204gat), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n947), .A2(new_n954), .A3(new_n603), .ZN(new_n955));
  XOR2_X1   g754(.A(new_n955), .B(KEYINPUT62), .Z(new_n956));
  OAI21_X1  g755(.A(G204gat), .B1(new_n950), .B2(new_n604), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(G1353gat));
  NAND3_X1  g757(.A1(new_n947), .A2(new_n203), .A3(new_n680), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n951), .A2(new_n680), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n960), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g761(.A(KEYINPUT63), .B1(new_n960), .B2(G211gat), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(G1354gat));
  OAI21_X1  g763(.A(new_n621), .B1(new_n951), .B2(KEYINPUT127), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT127), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n950), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g766(.A(G218gat), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n947), .A2(new_n204), .A3(new_n621), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(G1355gat));
endmodule


