//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 0 1 0 1 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(G143), .B(G146), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT67), .B(G128), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT1), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n188), .B1(new_n189), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT1), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  AND4_X1   g010(.A1(new_n194), .A2(new_n191), .A3(new_n196), .A4(G128), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n193), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(G125), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n191), .A2(new_n196), .A3(KEYINPUT0), .A4(G128), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n188), .A2(KEYINPUT64), .A3(KEYINPUT0), .A4(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n188), .ZN(new_n206));
  XOR2_X1   g020(.A(KEYINPUT0), .B(G128), .Z(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n200), .B1(G125), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G953), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G224), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT7), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n210), .B(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(G116), .B(G119), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT2), .B(G113), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n215), .B(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G101), .ZN(new_n218));
  INV_X1    g032(.A(G104), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(KEYINPUT3), .ZN(new_n220));
  OR2_X1    g034(.A1(KEYINPUT85), .A2(G107), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT85), .A2(G107), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT86), .A4(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G104), .ZN(new_n225));
  AND2_X1   g039(.A1(KEYINPUT85), .A2(G107), .ZN(new_n226));
  NOR2_X1   g040(.A1(KEYINPUT85), .A2(G107), .ZN(new_n227));
  NOR3_X1   g041(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT3), .B1(new_n219), .B2(G107), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT86), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n223), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n219), .A2(G107), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n218), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT4), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n217), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT87), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n233), .A2(new_n218), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n239));
  INV_X1    g053(.A(G107), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G104), .ZN(new_n241));
  AOI21_X1  g055(.A(KEYINPUT86), .B1(new_n241), .B2(KEYINPUT3), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  AOI211_X1 g057(.A(new_n237), .B(new_n238), .C1(new_n243), .C2(new_n223), .ZN(new_n244));
  INV_X1    g058(.A(new_n238), .ZN(new_n245));
  AOI21_X1  g059(.A(KEYINPUT87), .B1(new_n232), .B2(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  AOI22_X1  g061(.A1(new_n243), .A2(new_n223), .B1(new_n219), .B2(G107), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT4), .B1(new_n248), .B2(new_n218), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n236), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n221), .A2(new_n222), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n219), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n218), .B1(new_n252), .B2(new_n241), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n215), .A2(KEYINPUT5), .ZN(new_n255));
  INV_X1    g069(.A(G116), .ZN(new_n256));
  NOR3_X1   g070(.A1(new_n256), .A2(KEYINPUT5), .A3(G119), .ZN(new_n257));
  INV_X1    g071(.A(G113), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n216), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n255), .A2(new_n259), .B1(new_n260), .B2(new_n215), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n254), .B(new_n261), .C1(new_n244), .C2(new_n246), .ZN(new_n262));
  XNOR2_X1  g076(.A(G110), .B(G122), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n250), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n214), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n254), .B1(new_n244), .B2(new_n246), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n266), .B(new_n261), .ZN(new_n267));
  XOR2_X1   g081(.A(new_n263), .B(KEYINPUT8), .Z(new_n268));
  OR2_X1    g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(G902), .B1(new_n265), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n250), .A2(new_n262), .ZN(new_n271));
  INV_X1    g085(.A(new_n263), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  XOR2_X1   g087(.A(KEYINPUT96), .B(KEYINPUT6), .Z(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n264), .A2(KEYINPUT6), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n263), .B1(new_n250), .B2(new_n262), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT95), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT95), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n273), .A2(new_n279), .A3(KEYINPUT6), .A4(new_n264), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n275), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT97), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n210), .B(new_n212), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n282), .B1(new_n281), .B2(new_n283), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n187), .B(new_n270), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT99), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n270), .B1(new_n284), .B2(new_n285), .ZN(new_n288));
  XOR2_X1   g102(.A(new_n187), .B(KEYINPUT98), .Z(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n278), .A2(new_n280), .ZN(new_n291));
  INV_X1    g105(.A(new_n275), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n292), .A3(new_n283), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT97), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT99), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n296), .A2(new_n297), .A3(new_n187), .A4(new_n270), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n287), .A2(new_n290), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G214), .B1(G237), .B2(G902), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G952), .ZN(new_n302));
  AOI211_X1 g116(.A(G953), .B(new_n302), .C1(G234), .C2(G237), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT75), .B(G902), .ZN(new_n304));
  AOI211_X1 g118(.A(new_n211), .B(new_n304), .C1(G234), .C2(G237), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT21), .B(G898), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n256), .A2(G122), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n240), .B1(new_n308), .B2(KEYINPUT14), .ZN(new_n309));
  XNOR2_X1  g123(.A(G116), .B(G122), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n309), .B1(KEYINPUT14), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G128), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n313), .A2(G143), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n314), .B(KEYINPUT104), .ZN(new_n315));
  XOR2_X1   g129(.A(KEYINPUT67), .B(G128), .Z(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G143), .ZN(new_n317));
  INV_X1    g131(.A(G134), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n315), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n318), .B1(new_n315), .B2(new_n317), .ZN(new_n320));
  OAI221_X1 g134(.A(new_n312), .B1(new_n251), .B2(new_n311), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT13), .ZN(new_n322));
  OR2_X1    g136(.A1(new_n315), .A2(new_n322), .ZN(new_n323));
  AOI22_X1  g137(.A1(new_n315), .A2(new_n322), .B1(G143), .B2(new_n316), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n318), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n251), .B(new_n310), .ZN(new_n326));
  OR2_X1    g140(.A1(new_n319), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n321), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT9), .B(G234), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(G217), .A3(new_n211), .ZN(new_n331));
  OR2_X1    g145(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT105), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n328), .A2(new_n331), .ZN(new_n335));
  OR3_X1    g149(.A1(new_n328), .A2(new_n333), .A3(new_n331), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n304), .ZN(new_n338));
  INV_X1    g152(.A(G478), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT106), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n340), .A2(KEYINPUT15), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(KEYINPUT15), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n339), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n338), .B(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G902), .ZN(new_n346));
  INV_X1    g160(.A(G237), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(new_n211), .A3(G214), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n348), .B(new_n195), .ZN(new_n349));
  OR2_X1    g163(.A1(new_n349), .A2(G131), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(G131), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  MUX2_X1   g166(.A(new_n352), .B(new_n351), .S(KEYINPUT17), .Z(new_n353));
  INV_X1    g167(.A(G140), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G125), .ZN(new_n355));
  INV_X1    g169(.A(G125), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G140), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n355), .A2(new_n357), .A3(KEYINPUT16), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT77), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT77), .B1(new_n355), .B2(KEYINPUT16), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n360), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n362), .B(new_n190), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT103), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n362), .B(G146), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT103), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n353), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(G113), .B(G122), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n369), .B(new_n219), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n349), .B1(KEYINPUT18), .B2(G131), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n355), .A2(new_n357), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT101), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n372), .B(new_n373), .ZN(new_n374));
  OR2_X1    g188(.A1(new_n374), .A2(new_n190), .ZN(new_n375));
  INV_X1    g189(.A(new_n372), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n190), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n371), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n349), .A2(KEYINPUT18), .A3(G131), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(KEYINPUT100), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n368), .A2(new_n370), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n370), .B1(new_n368), .B2(new_n381), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n346), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G475), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n362), .A2(G146), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n376), .A2(KEYINPUT19), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n388), .B1(new_n374), .B2(KEYINPUT19), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n352), .B(new_n387), .C1(G146), .C2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n381), .A2(new_n390), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n391), .A2(KEYINPUT102), .ZN(new_n392));
  INV_X1    g206(.A(new_n370), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n393), .B1(new_n391), .B2(KEYINPUT102), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n382), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT20), .ZN(new_n396));
  NOR2_X1   g210(.A1(G475), .A2(G902), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n396), .B1(new_n395), .B2(new_n397), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n386), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OR2_X1    g214(.A1(new_n345), .A2(new_n400), .ZN(new_n401));
  NOR3_X1   g215(.A1(new_n301), .A2(new_n307), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n304), .ZN(new_n403));
  INV_X1    g217(.A(G234), .ZN(new_n404));
  OAI21_X1  g218(.A(G217), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n313), .A2(G119), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT23), .ZN(new_n408));
  INV_X1    g222(.A(G119), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n408), .B1(new_n409), .B2(G128), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n316), .A2(G119), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n407), .B(new_n410), .C1(new_n411), .C2(new_n408), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G110), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT76), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n411), .A2(new_n414), .A3(new_n407), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n189), .A2(new_n409), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT76), .B1(new_n416), .B2(new_n406), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(KEYINPUT24), .B(G110), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n413), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n363), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n211), .A2(G221), .A3(G234), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n423), .B(KEYINPUT79), .ZN(new_n424));
  XNOR2_X1  g238(.A(KEYINPUT22), .B(G137), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n424), .B(new_n425), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n412), .A2(G110), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n418), .A2(new_n419), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT78), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n412), .A2(G110), .ZN(new_n431));
  INV_X1    g245(.A(new_n419), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n432), .B1(new_n415), .B2(new_n417), .ZN(new_n433));
  OAI21_X1  g247(.A(KEYINPUT78), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n387), .A2(new_n377), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n422), .B(new_n426), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n426), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n436), .B1(new_n430), .B2(new_n434), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n438), .B1(new_n439), .B2(new_n421), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n437), .A2(new_n440), .A3(new_n304), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT80), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT25), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n405), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n441), .A2(new_n442), .A3(KEYINPUT25), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT81), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT81), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n445), .A2(new_n449), .A3(new_n446), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n437), .A2(new_n440), .ZN(new_n451));
  XOR2_X1   g265(.A(new_n451), .B(KEYINPUT82), .Z(new_n452));
  NAND2_X1  g266(.A1(new_n405), .A2(new_n346), .ZN(new_n453));
  XOR2_X1   g267(.A(new_n453), .B(KEYINPUT83), .Z(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n448), .A2(new_n450), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(G472), .A2(G902), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT11), .B1(new_n318), .B2(G137), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT11), .ZN(new_n461));
  INV_X1    g275(.A(G137), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n461), .A2(new_n462), .A3(G134), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(G131), .ZN(new_n465));
  OAI21_X1  g279(.A(KEYINPUT65), .B1(new_n462), .B2(G134), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT65), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(new_n318), .A3(G137), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n464), .A2(new_n465), .A3(new_n466), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT66), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n466), .A2(new_n468), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT66), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n471), .A2(new_n472), .A3(new_n465), .A4(new_n464), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n189), .A2(new_n192), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n206), .ZN(new_n476));
  INV_X1    g290(.A(new_n197), .ZN(new_n477));
  XOR2_X1   g291(.A(G134), .B(G137), .Z(new_n478));
  AOI22_X1  g292(.A1(new_n476), .A2(new_n477), .B1(G131), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT68), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n474), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n471), .A2(new_n464), .ZN(new_n482));
  AOI22_X1  g296(.A1(new_n470), .A2(new_n473), .B1(G131), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n481), .B1(new_n483), .B2(new_n209), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n478), .A2(G131), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n485), .B1(new_n193), .B2(new_n197), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n486), .B1(new_n473), .B2(new_n470), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n487), .A2(new_n480), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT30), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n482), .A2(G131), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n474), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n209), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT30), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n474), .A2(new_n479), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n489), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n217), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n495), .A2(KEYINPUT68), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n500), .A2(new_n493), .A3(new_n217), .A4(new_n481), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n347), .A2(new_n211), .A3(G210), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(KEYINPUT27), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT26), .B(G101), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n503), .B(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT69), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT69), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n501), .A2(new_n508), .A3(new_n505), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n499), .A2(KEYINPUT70), .A3(new_n507), .A4(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT31), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n217), .B1(new_n489), .B2(new_n496), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n501), .A2(new_n508), .A3(new_n505), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n515), .A2(KEYINPUT70), .A3(KEYINPUT31), .A4(new_n507), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT72), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n483), .A2(new_n209), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n498), .B1(new_n519), .B2(new_n487), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n501), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT28), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT71), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT71), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n521), .A2(new_n524), .A3(KEYINPUT28), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n519), .A2(new_n498), .A3(new_n487), .ZN(new_n526));
  OR2_X1    g340(.A1(new_n526), .A2(KEYINPUT28), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n523), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n505), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n517), .A2(new_n518), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n518), .B1(new_n517), .B2(new_n530), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n459), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT32), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT32), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n535), .B(new_n459), .C1(new_n531), .C2(new_n532), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n526), .A2(KEYINPUT28), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n498), .B1(new_n484), .B2(new_n488), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n501), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n538), .B1(new_n540), .B2(KEYINPUT28), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT29), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n529), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  OR2_X1    g358(.A1(new_n544), .A2(KEYINPUT74), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(KEYINPUT74), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n403), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n501), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n513), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n549), .A2(new_n505), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(KEYINPUT73), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n542), .B1(new_n528), .B2(new_n529), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n547), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(G472), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n458), .B1(new_n537), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(G221), .B1(new_n329), .B2(G902), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n313), .B1(new_n191), .B2(KEYINPUT1), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n477), .B1(new_n188), .B2(new_n559), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n254), .B(new_n560), .C1(new_n244), .C2(new_n246), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT10), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n209), .B1(new_n234), .B2(new_n235), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n564), .B1(new_n247), .B2(new_n249), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n198), .A2(new_n562), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n566), .B(new_n254), .C1(new_n244), .C2(new_n246), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n563), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(new_n491), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n232), .A2(new_n245), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n237), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n232), .A2(KEYINPUT87), .A3(new_n245), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n253), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OAI211_X1 g388(.A(KEYINPUT89), .B(new_n561), .C1(new_n574), .C2(new_n199), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT89), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n266), .A2(new_n576), .A3(new_n198), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n575), .A2(KEYINPUT88), .A3(new_n491), .A4(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT90), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n579), .A3(KEYINPUT12), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n578), .A2(new_n579), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n575), .A2(KEYINPUT90), .A3(new_n491), .A4(new_n577), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT12), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n570), .B(new_n580), .C1(new_n581), .C2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT91), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(G110), .B(G140), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(KEYINPUT84), .ZN(new_n589));
  INV_X1    g403(.A(G227), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(G953), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n589), .B(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n578), .A2(new_n579), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(new_n583), .A3(new_n582), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n594), .A2(KEYINPUT91), .A3(new_n570), .A4(new_n580), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n587), .A2(new_n592), .A3(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n569), .A2(new_n592), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  OR2_X1    g412(.A1(new_n598), .A2(KEYINPUT92), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT93), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n568), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n563), .A2(new_n565), .A3(KEYINPUT93), .A4(new_n567), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n491), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n598), .A2(KEYINPUT92), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n599), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n596), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT94), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n596), .A2(KEYINPUT94), .A3(new_n605), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(G469), .A3(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(G469), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(new_n346), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n603), .A2(new_n570), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n592), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n597), .B(new_n580), .C1(new_n581), .C2(new_n584), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n403), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n612), .B1(new_n616), .B2(new_n611), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n558), .B1(new_n610), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n402), .A2(new_n556), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G101), .ZN(G3));
  OAI21_X1  g434(.A(new_n304), .B1(new_n531), .B2(new_n532), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(G472), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n622), .A2(new_n533), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n457), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n337), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n332), .A2(KEYINPUT33), .A3(new_n335), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n403), .A2(new_n339), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n338), .A2(new_n339), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n307), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n632), .A2(new_n400), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n187), .B1(new_n296), .B2(new_n270), .ZN(new_n635));
  INV_X1    g449(.A(new_n187), .ZN(new_n636));
  INV_X1    g450(.A(new_n270), .ZN(new_n637));
  AOI211_X1 g451(.A(new_n636), .B(new_n637), .C1(new_n294), .C2(new_n295), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n634), .B(new_n300), .C1(new_n635), .C2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(KEYINPUT107), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n288), .A2(new_n636), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n286), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT107), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n642), .A2(new_n643), .A3(new_n300), .A4(new_n634), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n625), .A2(new_n618), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT34), .B(G104), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  INV_X1    g462(.A(new_n300), .ZN(new_n649));
  INV_X1    g463(.A(new_n400), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n650), .A2(new_n633), .A3(new_n345), .ZN(new_n651));
  AOI211_X1 g465(.A(new_n649), .B(new_n651), .C1(new_n286), .C2(new_n641), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n625), .A2(new_n618), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT35), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  AND2_X1   g469(.A1(new_n448), .A2(new_n450), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n439), .A2(new_n421), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n438), .A2(KEYINPUT36), .ZN(new_n658));
  XOR2_X1   g472(.A(new_n657), .B(new_n658), .Z(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n455), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n402), .A2(new_n618), .A3(new_n623), .A4(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT37), .B(G110), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G12));
  AND2_X1   g478(.A1(new_n656), .A2(new_n660), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n665), .B1(new_n537), .B2(new_n555), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n649), .B1(new_n641), .B2(new_n286), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n650), .A2(new_n345), .ZN(new_n668));
  INV_X1    g482(.A(G900), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n305), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n670), .A2(KEYINPUT108), .ZN(new_n671));
  INV_X1    g485(.A(new_n303), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n670), .A2(KEYINPUT108), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n668), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n666), .A2(new_n618), .A3(new_n667), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G128), .ZN(G30));
  AND2_X1   g491(.A1(new_n515), .A2(new_n507), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n678), .B1(new_n529), .B2(new_n540), .ZN(new_n679));
  OAI21_X1  g493(.A(G472), .B1(new_n679), .B2(G902), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n537), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n345), .A2(new_n400), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n681), .A2(new_n300), .A3(new_n665), .A4(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT109), .B(KEYINPUT38), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n299), .B(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(new_n674), .B(KEYINPUT39), .Z(new_n687));
  NAND2_X1  g501(.A1(new_n618), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n686), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G143), .ZN(G45));
  INV_X1    g506(.A(new_n632), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n693), .A2(new_n650), .A3(new_n674), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n666), .A2(new_n618), .A3(new_n667), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G146), .ZN(G48));
  NAND2_X1  g510(.A1(new_n616), .A2(new_n611), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n557), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT111), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT110), .ZN(new_n700));
  OAI21_X1  g514(.A(G469), .B1(new_n616), .B2(new_n700), .ZN(new_n701));
  AOI211_X1 g515(.A(KEYINPUT110), .B(new_n403), .C1(new_n614), .C2(new_n615), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n699), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n614), .A2(new_n615), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n304), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(KEYINPUT110), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n616), .A2(new_n700), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n706), .A2(KEYINPUT111), .A3(G469), .A4(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n698), .B1(new_n703), .B2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n556), .A2(new_n645), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT41), .B(G113), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G15));
  NAND2_X1  g526(.A1(new_n517), .A2(new_n530), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT72), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n517), .A2(new_n518), .A3(new_n530), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n535), .B1(new_n716), .B2(new_n459), .ZN(new_n717));
  INV_X1    g531(.A(new_n536), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n555), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n719), .A2(new_n652), .A3(new_n457), .A4(new_n709), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G116), .ZN(G18));
  NAND2_X1  g535(.A1(new_n703), .A2(new_n708), .ZN(new_n722));
  INV_X1    g536(.A(new_n698), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n722), .A2(new_n667), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n401), .A2(new_n307), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n724), .A2(new_n719), .A3(new_n725), .A4(new_n661), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G119), .ZN(G21));
  OAI21_X1  g541(.A(new_n517), .B1(new_n505), .B2(new_n541), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n459), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n403), .B1(new_n714), .B2(new_n715), .ZN(new_n730));
  INV_X1    g544(.A(G472), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n457), .B(new_n729), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n667), .A2(new_n682), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n733), .A2(new_n734), .A3(new_n633), .A4(new_n709), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  NAND2_X1  g550(.A1(new_n709), .A2(new_n667), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n661), .A2(new_n622), .A3(new_n694), .A4(new_n729), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n356), .ZN(G27));
  OAI21_X1  g554(.A(new_n617), .B1(new_n606), .B2(new_n611), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n558), .A2(new_n649), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n299), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n719), .A2(new_n744), .A3(new_n457), .A4(new_n694), .ZN(new_n745));
  XNOR2_X1  g559(.A(KEYINPUT112), .B(KEYINPUT42), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(KEYINPUT42), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n556), .A2(new_n694), .A3(new_n744), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(KEYINPUT113), .B(G131), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G33));
  NAND3_X1  g569(.A1(new_n556), .A2(new_n675), .A3(new_n744), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G134), .ZN(G36));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n596), .A2(KEYINPUT94), .A3(new_n605), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT94), .B1(new_n596), .B2(new_n605), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n606), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n611), .B1(new_n762), .B2(KEYINPUT45), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n612), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n697), .B1(new_n764), .B2(KEYINPUT46), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT46), .ZN(new_n766));
  AOI211_X1 g580(.A(new_n766), .B(new_n612), .C1(new_n761), .C2(new_n763), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n557), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n687), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n693), .A2(new_n400), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT43), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n661), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT44), .ZN(new_n774));
  OR3_X1    g588(.A1(new_n773), .A2(new_n623), .A3(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n774), .B1(new_n773), .B2(new_n623), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n299), .A2(new_n649), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n770), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(new_n462), .ZN(G39));
  INV_X1    g594(.A(KEYINPUT47), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n768), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(KEYINPUT47), .B(new_n557), .C1(new_n765), .C2(new_n767), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AOI22_X1  g598(.A1(new_n534), .A2(new_n536), .B1(new_n554), .B2(G472), .ZN(new_n785));
  AND4_X1   g599(.A1(new_n458), .A2(new_n785), .A3(new_n694), .A4(new_n777), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G140), .ZN(G42));
  NAND3_X1  g602(.A1(new_n733), .A2(new_n303), .A3(new_n772), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n789), .A2(new_n649), .A3(new_n299), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n782), .A2(KEYINPUT118), .A3(new_n783), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n722), .A2(new_n558), .A3(new_n697), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT118), .B1(new_n782), .B2(new_n783), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n790), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n722), .A2(new_n723), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n672), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n777), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n537), .A2(new_n457), .A3(new_n680), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n632), .A2(new_n400), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n797), .A2(new_n772), .A3(new_n777), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n661), .A2(new_n622), .A3(new_n729), .ZN(new_n803));
  AOI22_X1  g617(.A1(new_n800), .A2(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n789), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n796), .A2(new_n300), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n805), .A2(KEYINPUT50), .A3(new_n685), .A4(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT50), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n685), .A2(new_n806), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n808), .B1(new_n809), .B2(new_n789), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n804), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT51), .B1(new_n795), .B2(new_n813), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n804), .A2(new_n811), .A3(KEYINPUT51), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n782), .A2(new_n792), .A3(new_n783), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n790), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n797), .A2(new_n772), .A3(new_n777), .ZN(new_n819));
  INV_X1    g633(.A(new_n556), .ZN(new_n820));
  OR3_X1    g634(.A1(new_n819), .A2(KEYINPUT48), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(KEYINPUT48), .B1(new_n819), .B2(new_n820), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI211_X1 g637(.A(new_n302), .B(G953), .C1(new_n805), .C2(new_n724), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n693), .A2(new_n650), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n800), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n818), .A2(new_n823), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT119), .B1(new_n814), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n827), .A2(new_n823), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n830), .B1(new_n815), .B2(new_n817), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT119), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n784), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n834), .A2(new_n791), .A3(new_n792), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n812), .B1(new_n835), .B2(new_n790), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n831), .B(new_n832), .C1(new_n836), .C2(KEYINPUT51), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n829), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n739), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n674), .A2(new_n558), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n741), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n681), .A2(new_n665), .A3(new_n734), .A4(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n676), .A2(new_n695), .A3(new_n839), .A4(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT52), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n846));
  INV_X1    g660(.A(new_n675), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n785), .A2(new_n847), .A3(new_n665), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n618), .A2(new_n667), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n739), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n850), .A2(KEYINPUT52), .A3(new_n695), .A4(new_n842), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n845), .A2(new_n846), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n843), .A2(KEYINPUT116), .A3(new_n844), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n642), .A2(new_n633), .A3(new_n300), .A4(new_n682), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n796), .A2(new_n855), .A3(new_n732), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n785), .A2(new_n796), .A3(new_n458), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n856), .B1(new_n857), .B2(new_n645), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT114), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n858), .A2(new_n859), .A3(new_n720), .A4(new_n726), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n710), .A2(new_n726), .A3(new_n720), .A4(new_n735), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT114), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n825), .B1(new_n345), .B2(new_n650), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n301), .A2(new_n864), .A3(new_n307), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n625), .A2(new_n865), .A3(new_n618), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n866), .A2(new_n619), .A3(new_n662), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n738), .A2(new_n299), .A3(new_n743), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n401), .A2(new_n674), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n618), .A2(new_n777), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n869), .B1(new_n871), .B2(new_n666), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n753), .A2(new_n872), .A3(new_n756), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n863), .A2(new_n868), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n854), .B1(KEYINPUT115), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n867), .B1(new_n860), .B2(new_n862), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT115), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n876), .A2(new_n877), .A3(new_n873), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT53), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n845), .A2(new_n851), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n876), .A2(new_n873), .A3(new_n880), .ZN(new_n881));
  XOR2_X1   g695(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n882));
  NOR2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT54), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n881), .A2(new_n882), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n867), .A2(new_n886), .A3(new_n861), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n852), .A2(new_n873), .A3(new_n887), .A4(new_n853), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT54), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n885), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n838), .A2(KEYINPUT120), .A3(new_n884), .A4(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT120), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n874), .A2(KEYINPUT115), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n852), .A2(new_n853), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n893), .A2(new_n894), .A3(new_n878), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n883), .B1(new_n895), .B2(new_n886), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n890), .B1(new_n896), .B2(new_n889), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n829), .A2(new_n837), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n892), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n302), .A2(new_n211), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n891), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n685), .A2(new_n742), .A3(new_n771), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n722), .A2(new_n697), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n799), .B1(KEYINPUT49), .B2(new_n903), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n902), .B(new_n904), .C1(KEYINPUT49), .C2(new_n903), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n901), .A2(new_n905), .ZN(G75));
  NOR2_X1   g720(.A1(new_n211), .A2(G952), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n304), .B1(new_n885), .B2(new_n888), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT56), .B1(new_n909), .B2(new_n636), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n281), .B(new_n283), .Z(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT55), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n908), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n909), .A2(new_n289), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT121), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n909), .A2(KEYINPUT121), .A3(new_n289), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT56), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n912), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n916), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT122), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n916), .A2(KEYINPUT122), .A3(new_n917), .A4(new_n919), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n913), .B1(new_n922), .B2(new_n923), .ZN(G51));
  NAND2_X1  g738(.A1(new_n885), .A2(new_n888), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(KEYINPUT54), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n890), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n612), .B(KEYINPUT57), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n704), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n909), .A2(new_n761), .A3(new_n763), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n907), .B1(new_n930), .B2(new_n931), .ZN(G54));
  AND3_X1   g746(.A1(new_n909), .A2(KEYINPUT58), .A3(G475), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n908), .B1(new_n933), .B2(new_n395), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n934), .B1(new_n395), .B2(new_n933), .ZN(G60));
  AND2_X1   g749(.A1(new_n627), .A2(new_n628), .ZN(new_n936));
  NAND2_X1  g750(.A1(G478), .A2(G902), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT59), .Z(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n936), .B1(new_n897), .B2(new_n939), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n927), .A2(new_n936), .A3(new_n939), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n940), .A2(new_n941), .A3(new_n907), .ZN(G63));
  NAND2_X1  g756(.A1(G217), .A2(G902), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT60), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n885), .B2(new_n888), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n659), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n946), .B(new_n908), .C1(new_n452), .C2(new_n945), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT61), .Z(G66));
  OR2_X1    g762(.A1(new_n876), .A2(G953), .ZN(new_n949));
  INV_X1    g763(.A(G224), .ZN(new_n950));
  OAI21_X1  g764(.A(G953), .B1(new_n306), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n949), .A2(KEYINPUT123), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n952), .B1(KEYINPUT123), .B2(new_n949), .ZN(new_n953));
  INV_X1    g767(.A(G898), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n281), .B1(new_n954), .B2(G953), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n953), .B(new_n955), .ZN(G69));
  XOR2_X1   g770(.A(new_n497), .B(new_n389), .Z(new_n957));
  AND2_X1   g771(.A1(new_n850), .A2(new_n695), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n691), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n864), .A2(new_n649), .A3(new_n299), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n961), .A2(new_n556), .A3(new_n618), .A4(new_n687), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n787), .B1(new_n770), .B2(new_n778), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n963), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n957), .B1(new_n967), .B2(new_n211), .ZN(new_n968));
  OR2_X1    g782(.A1(new_n968), .A2(KEYINPUT124), .ZN(new_n969));
  OAI21_X1  g783(.A(G953), .B1(new_n590), .B2(new_n669), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT125), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n957), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n958), .A2(new_n753), .A3(new_n756), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n769), .A2(new_n556), .A3(new_n687), .A4(new_n734), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n211), .B1(new_n976), .B2(new_n964), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n211), .A2(G900), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n973), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(KEYINPUT124), .B1(new_n968), .B2(new_n980), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n969), .A2(new_n972), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n972), .B1(new_n969), .B2(new_n981), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n982), .A2(new_n983), .ZN(G72));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT63), .Z(new_n986));
  OAI21_X1  g800(.A(new_n986), .B1(new_n552), .B2(new_n678), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n965), .A2(new_n876), .A3(new_n975), .A4(new_n974), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n988), .A2(new_n986), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n549), .A2(new_n529), .ZN(new_n990));
  OAI221_X1 g804(.A(new_n908), .B1(new_n896), .B2(new_n987), .C1(new_n989), .C2(new_n990), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n549), .A2(new_n529), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n963), .A2(new_n965), .A3(new_n876), .A4(new_n966), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n993), .A2(KEYINPUT126), .A3(new_n986), .ZN(new_n994));
  AOI21_X1  g808(.A(KEYINPUT126), .B1(new_n993), .B2(new_n986), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT127), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI211_X1 g812(.A(KEYINPUT127), .B(new_n992), .C1(new_n994), .C2(new_n995), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n991), .B1(new_n998), .B2(new_n999), .ZN(G57));
endmodule


