//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 1 0 1 0 0 1 0 0 0 0 0 1 1 0 1 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 1 1 1 0 1 0 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1228, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G50), .A2(G226), .ZN(new_n207));
  INV_X1    g0007(.A(G116), .ZN(new_n208));
  INV_X1    g0008(.A(G270), .ZN(new_n209));
  OAI21_X1  g0009(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AOI21_X1  g0010(.A(new_n210), .B1(G58), .B2(G232), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G87), .A2(G250), .ZN(new_n213));
  AND2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G68), .A2(G238), .ZN(new_n215));
  XOR2_X1   g0015(.A(KEYINPUT66), .B(G244), .Z(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G77), .ZN(new_n217));
  NAND4_X1  g0017(.A1(new_n211), .A2(new_n214), .A3(new_n215), .A4(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G20), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT1), .Z(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(KEYINPUT65), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT65), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G20), .ZN(new_n225));
  AND2_X1   g0025(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(G50), .B1(G58), .B2(G68), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n226), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n219), .A2(G13), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n232), .B(G250), .C1(G257), .C2(G264), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT0), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n221), .A2(new_n231), .A3(new_n234), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G226), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G264), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n209), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G358));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G97), .B(G107), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(G87), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(new_n208), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  XNOR2_X1  g0052(.A(KEYINPUT69), .B(G58), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT8), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(KEYINPUT8), .B2(G58), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n227), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(G1), .B2(new_n222), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G13), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n261), .A2(new_n222), .A3(G1), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n260), .B1(new_n262), .B2(new_n255), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT3), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G33), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT68), .ZN(new_n269));
  AND3_X1   g0069(.A1(new_n266), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n269), .B1(new_n266), .B2(new_n268), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(KEYINPUT7), .B1(new_n272), .B2(new_n222), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n267), .A2(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n275));
  OAI21_X1  g0075(.A(KEYINPUT7), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(KEYINPUT76), .B1(new_n276), .B2(new_n226), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT7), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n278), .B1(new_n266), .B2(new_n268), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT76), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n223), .A2(new_n225), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(G68), .B1(new_n273), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n201), .B1(new_n253), .B2(G68), .ZN(new_n285));
  INV_X1    g0085(.A(G159), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI22_X1  g0088(.A1(new_n285), .A2(new_n222), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n264), .B1(new_n284), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT74), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n266), .A2(new_n268), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n274), .A2(KEYINPUT74), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(new_n294), .A3(new_n222), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT7), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n265), .A2(KEYINPUT74), .A3(KEYINPUT3), .ZN(new_n297));
  XNOR2_X1  g0097(.A(KEYINPUT3), .B(G33), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n297), .B1(new_n298), .B2(new_n292), .ZN(new_n299));
  AOI21_X1  g0099(.A(KEYINPUT7), .B1(new_n223), .B2(new_n225), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n296), .A2(new_n301), .A3(G68), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(new_n290), .A3(KEYINPUT16), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n257), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n263), .B1(new_n291), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n293), .A2(new_n294), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n306), .A2(G226), .A3(G1698), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT77), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(G1698), .B1(new_n293), .B2(new_n294), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n310), .A2(G223), .B1(G33), .B2(G87), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n306), .A2(KEYINPUT77), .A3(G226), .A4(G1698), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n309), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n314), .ZN(new_n316));
  INV_X1    g0116(.A(G1), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(G41), .B2(G45), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G232), .ZN(new_n320));
  INV_X1    g0120(.A(G274), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  AND4_X1   g0123(.A1(G179), .A2(new_n315), .A3(new_n320), .A4(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G169), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n322), .B1(new_n313), .B2(new_n314), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n325), .B1(new_n326), .B2(new_n320), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n305), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n328), .B(KEYINPUT18), .ZN(new_n329));
  INV_X1    g0129(.A(new_n264), .ZN(new_n330));
  INV_X1    g0130(.A(G68), .ZN(new_n331));
  AND3_X1   g0131(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n280), .B1(new_n279), .B2(new_n281), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n298), .A2(new_n269), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT68), .B1(new_n274), .B2(new_n275), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(new_n336), .A3(new_n222), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n278), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n331), .B1(new_n334), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n330), .B1(new_n339), .B2(new_n289), .ZN(new_n340));
  AOI22_X1  g0140(.A1(KEYINPUT7), .A2(new_n295), .B1(new_n299), .B2(new_n300), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n289), .B1(new_n341), .B2(G68), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n258), .B1(new_n342), .B2(KEYINPUT16), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n315), .A2(G190), .A3(new_n320), .A4(new_n323), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n344), .A2(new_n263), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n320), .ZN(new_n347));
  AOI211_X1 g0147(.A(new_n347), .B(new_n322), .C1(new_n313), .C2(new_n314), .ZN(new_n348));
  INV_X1    g0148(.A(G200), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT17), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n263), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(new_n340), .B2(new_n343), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n315), .A2(new_n320), .A3(new_n323), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G200), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT17), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n353), .A2(new_n355), .A3(new_n356), .A4(new_n345), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n351), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT78), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n351), .A2(KEYINPUT78), .A3(new_n357), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n329), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n319), .A2(new_n216), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n335), .A2(new_n336), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n364), .A2(G238), .A3(G1698), .ZN(new_n365));
  INV_X1    g0165(.A(G1698), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(G232), .A3(new_n366), .ZN(new_n367));
  XOR2_X1   g0167(.A(KEYINPUT70), .B(G107), .Z(new_n368));
  OAI211_X1 g0168(.A(new_n365), .B(new_n367), .C1(new_n364), .C2(new_n368), .ZN(new_n369));
  AOI211_X1 g0169(.A(new_n322), .B(new_n363), .C1(new_n369), .C2(new_n314), .ZN(new_n370));
  OR2_X1    g0170(.A1(new_n370), .A2(G169), .ZN(new_n371));
  INV_X1    g0171(.A(G179), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  XOR2_X1   g0173(.A(KEYINPUT8), .B(G58), .Z(new_n374));
  OR2_X1    g0174(.A1(new_n287), .A2(KEYINPUT71), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n287), .A2(KEYINPUT71), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G77), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n281), .A2(G33), .ZN(new_n379));
  XOR2_X1   g0179(.A(KEYINPUT15), .B(G87), .Z(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  OAI221_X1 g0181(.A(new_n377), .B1(new_n378), .B2(new_n281), .C1(new_n379), .C2(new_n381), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n382), .A2(new_n257), .B1(new_n378), .B2(new_n262), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n378), .B2(new_n259), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n371), .A2(new_n373), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n370), .A2(G190), .ZN(new_n386));
  INV_X1    g0186(.A(new_n384), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n386), .B(new_n387), .C1(new_n349), .C2(new_n370), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n362), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n203), .A2(G20), .ZN(new_n390));
  INV_X1    g0190(.A(G150), .ZN(new_n391));
  OAI221_X1 g0191(.A(new_n390), .B1(new_n391), .B2(new_n288), .C1(new_n255), .C2(new_n379), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n392), .A2(new_n257), .B1(new_n202), .B2(new_n262), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(new_n202), .B2(new_n259), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT9), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n364), .A2(G223), .A3(G1698), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n364), .A2(G222), .A3(new_n366), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n396), .B(new_n397), .C1(new_n378), .C2(new_n364), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n314), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n319), .A2(G226), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(new_n323), .A3(new_n400), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n394), .A2(new_n395), .B1(new_n401), .B2(G200), .ZN(new_n402));
  INV_X1    g0202(.A(new_n401), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G190), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n402), .B(new_n404), .C1(new_n395), .C2(new_n394), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n405), .B(KEYINPUT10), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT13), .ZN(new_n407));
  OAI211_X1 g0207(.A(G226), .B(new_n366), .C1(new_n270), .C2(new_n271), .ZN(new_n408));
  OAI211_X1 g0208(.A(G232), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G33), .A2(G97), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n314), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n319), .A2(G238), .ZN(new_n413));
  AND4_X1   g0213(.A1(new_n407), .A2(new_n412), .A3(new_n323), .A4(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n411), .A2(new_n314), .B1(G238), .B2(new_n319), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n407), .B1(new_n416), .B2(new_n323), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n415), .A2(new_n418), .A3(G190), .ZN(new_n419));
  OAI21_X1  g0219(.A(G200), .B1(new_n414), .B2(new_n417), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n331), .A2(G20), .ZN(new_n421));
  OAI221_X1 g0221(.A(new_n421), .B1(new_n202), .B2(new_n288), .C1(new_n379), .C2(new_n378), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n422), .A2(KEYINPUT11), .A3(new_n257), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(new_n331), .B2(new_n259), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n262), .A2(new_n331), .ZN(new_n425));
  XOR2_X1   g0225(.A(new_n425), .B(KEYINPUT12), .Z(new_n426));
  AOI21_X1  g0226(.A(KEYINPUT11), .B1(new_n422), .B2(new_n257), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n424), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n419), .A2(new_n420), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT72), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT72), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n419), .A2(new_n420), .A3(new_n431), .A4(new_n428), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n394), .B1(new_n401), .B2(G179), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(new_n325), .B2(new_n401), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n406), .A2(new_n430), .A3(new_n432), .A4(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(G169), .B1(new_n414), .B2(new_n417), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT14), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n415), .A2(new_n418), .A3(G179), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT14), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n440), .B(G169), .C1(new_n414), .C2(new_n417), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n438), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT73), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT73), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n438), .A2(new_n444), .A3(new_n439), .A4(new_n441), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n428), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n389), .A2(new_n436), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n262), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n448), .B(new_n258), .C1(G1), .C2(new_n265), .ZN(new_n449));
  INV_X1    g0249(.A(G107), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g0251(.A(KEYINPUT70), .B(G107), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(new_n222), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT23), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT22), .B1(KEYINPUT23), .B2(G107), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  OAI22_X1  g0256(.A1(new_n453), .A2(new_n454), .B1(new_n281), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT22), .ZN(new_n458));
  OAI21_X1  g0258(.A(G87), .B1(new_n270), .B2(new_n271), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  XNOR2_X1  g0260(.A(KEYINPUT84), .B(KEYINPUT24), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n222), .A2(G33), .A3(G116), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n306), .A2(KEYINPUT22), .A3(G87), .A4(new_n281), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n460), .A2(new_n461), .A3(new_n462), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n459), .A2(new_n458), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n368), .A2(G20), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n466), .A2(KEYINPUT23), .B1(new_n226), .B2(new_n455), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n465), .A2(new_n467), .A3(new_n462), .A4(new_n463), .ZN(new_n468));
  INV_X1    g0268(.A(new_n461), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n464), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n451), .B1(new_n471), .B2(new_n257), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n262), .A2(new_n450), .B1(KEYINPUT85), .B2(KEYINPUT25), .ZN(new_n473));
  NOR2_X1   g0273(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n474));
  XNOR2_X1  g0274(.A(new_n473), .B(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n306), .B1(G250), .B2(G1698), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n366), .A2(G257), .ZN(new_n478));
  INV_X1    g0278(.A(G294), .ZN(new_n479));
  OAI22_X1  g0279(.A1(new_n477), .A2(new_n478), .B1(new_n265), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n317), .A2(G45), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT80), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT5), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G41), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G41), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n317), .B(G45), .C1(new_n486), .C2(KEYINPUT5), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT80), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n486), .A2(KEYINPUT5), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT81), .ZN(new_n491));
  XNOR2_X1  g0291(.A(new_n490), .B(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n314), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n480), .A2(new_n314), .B1(G264), .B2(new_n493), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n489), .A2(new_n492), .A3(G274), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n316), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n325), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n494), .A2(new_n372), .A3(new_n496), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n476), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n272), .A2(G303), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G264), .A2(G1698), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT83), .B1(new_n299), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n310), .A2(G257), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT83), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n306), .A2(new_n505), .A3(G264), .A4(G1698), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n501), .A2(new_n503), .A3(new_n504), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n314), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n495), .A2(new_n316), .B1(new_n493), .B2(G270), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n325), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n262), .A2(new_n208), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n258), .B1(G20), .B2(new_n208), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G283), .ZN(new_n513));
  INV_X1    g0313(.A(G97), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n281), .B(new_n513), .C1(G33), .C2(new_n514), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n512), .A2(KEYINPUT20), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(KEYINPUT20), .B1(new_n512), .B2(new_n515), .ZN(new_n517));
  OAI221_X1 g0317(.A(new_n511), .B1(new_n208), .B2(new_n449), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n510), .A2(KEYINPUT21), .A3(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n518), .A2(G179), .A3(new_n509), .A4(new_n508), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT21), .B1(new_n510), .B2(new_n518), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n448), .A2(new_n380), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n306), .A2(G68), .A3(new_n281), .ZN(new_n525));
  XNOR2_X1  g0325(.A(KEYINPUT82), .B(KEYINPUT19), .ZN(new_n526));
  XNOR2_X1  g0326(.A(new_n526), .B(new_n410), .ZN(new_n527));
  NOR3_X1   g0327(.A1(new_n452), .A2(G87), .A3(G97), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n525), .B(new_n527), .C1(new_n281), .C2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n524), .B1(new_n529), .B2(new_n257), .ZN(new_n530));
  INV_X1    g0330(.A(new_n449), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n380), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n306), .A2(G238), .A3(new_n366), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n306), .A2(G244), .A3(G1698), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G33), .A2(G116), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n314), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n314), .A2(new_n481), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G250), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n481), .A2(G274), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n325), .B1(new_n538), .B2(new_n543), .ZN(new_n544));
  AOI211_X1 g0344(.A(new_n372), .B(new_n542), .C1(new_n537), .C2(new_n314), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n533), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(G87), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n449), .A2(new_n547), .ZN(new_n548));
  AOI211_X1 g0348(.A(new_n524), .B(new_n548), .C1(new_n529), .C2(new_n257), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n542), .B1(new_n537), .B2(new_n314), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G190), .ZN(new_n551));
  INV_X1    g0351(.A(G244), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n552), .B1(new_n293), .B2(new_n294), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n553), .A2(G1698), .B1(G33), .B2(G116), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n316), .B1(new_n554), .B2(new_n534), .ZN(new_n555));
  OAI21_X1  g0355(.A(G200), .B1(new_n555), .B2(new_n542), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n549), .A2(new_n551), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n546), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n500), .A2(new_n523), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n368), .B1(new_n334), .B2(new_n338), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n450), .A2(G97), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n514), .A2(G107), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT6), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n450), .A2(KEYINPUT6), .A3(G97), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n281), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n288), .A2(new_n378), .ZN(new_n568));
  OAI21_X1  g0368(.A(KEYINPUT79), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT79), .ZN(new_n570));
  INV_X1    g0370(.A(new_n568), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n450), .A2(KEYINPUT6), .A3(G97), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n249), .B2(new_n564), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n570), .B(new_n571), .C1(new_n573), .C2(new_n281), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n257), .B1(new_n561), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n448), .A2(G97), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n531), .A2(G97), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n576), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(G250), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n581));
  AND2_X1   g0381(.A1(KEYINPUT4), .A2(G244), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n366), .B(new_n582), .C1(new_n270), .C2(new_n271), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n581), .A2(new_n583), .A3(new_n513), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT4), .B1(new_n553), .B2(new_n366), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n314), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n495), .A2(new_n316), .B1(new_n493), .B2(G257), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n325), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n586), .A2(new_n587), .A3(new_n372), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n580), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n494), .A2(G190), .A3(new_n496), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n497), .A2(G200), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n472), .A2(new_n475), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n580), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n586), .A2(new_n587), .A3(G190), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n588), .A2(G200), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n508), .A2(new_n509), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n518), .B1(new_n599), .B2(G200), .ZN(new_n600));
  INV_X1    g0400(.A(G190), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n600), .B1(new_n601), .B2(new_n599), .ZN(new_n602));
  AND4_X1   g0402(.A1(new_n591), .A2(new_n594), .A3(new_n598), .A4(new_n602), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n447), .A2(new_n560), .A3(new_n603), .ZN(G372));
  AND3_X1   g0404(.A1(new_n580), .A2(new_n589), .A3(new_n590), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT26), .ZN(new_n606));
  OAI21_X1  g0406(.A(KEYINPUT86), .B1(new_n544), .B2(new_n545), .ZN(new_n607));
  OAI21_X1  g0407(.A(G169), .B1(new_n555), .B2(new_n542), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n538), .A2(G179), .A3(new_n543), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT86), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n607), .A2(new_n533), .A3(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n605), .A2(new_n606), .A3(new_n612), .A4(new_n557), .ZN(new_n613));
  OAI21_X1  g0413(.A(KEYINPUT26), .B1(new_n591), .B2(new_n558), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n614), .A3(new_n612), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT87), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n500), .A2(new_n523), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n598), .A2(new_n591), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n612), .A2(new_n557), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n618), .A2(new_n619), .A3(new_n594), .A4(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n613), .A2(new_n614), .A3(KEYINPUT87), .A4(new_n612), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n617), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n447), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n385), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n625), .A2(new_n429), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n351), .A2(KEYINPUT78), .A3(new_n357), .ZN(new_n627));
  AOI21_X1  g0427(.A(KEYINPUT78), .B1(new_n351), .B2(new_n357), .ZN(new_n628));
  OAI22_X1  g0428(.A1(new_n446), .A2(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT18), .ZN(new_n630));
  XNOR2_X1  g0430(.A(new_n328), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n434), .B1(new_n632), .B2(new_n406), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n624), .A2(new_n633), .ZN(G369));
  NOR2_X1   g0434(.A1(new_n226), .A2(new_n261), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  OR3_X1    g0436(.A1(new_n636), .A2(KEYINPUT27), .A3(G1), .ZN(new_n637));
  OAI21_X1  g0437(.A(KEYINPUT27), .B1(new_n636), .B2(G1), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(G213), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(G343), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n518), .ZN(new_n642));
  XNOR2_X1  g0442(.A(new_n523), .B(new_n642), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n643), .A2(new_n602), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(G330), .ZN(new_n645));
  INV_X1    g0445(.A(new_n500), .ZN(new_n646));
  INV_X1    g0446(.A(new_n641), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n594), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n647), .B1(new_n472), .B2(new_n475), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n500), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n645), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n523), .A2(new_n641), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n651), .A2(new_n655), .B1(new_n646), .B2(new_n647), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n654), .A2(new_n656), .ZN(G399));
  INV_X1    g0457(.A(new_n232), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n658), .A2(G41), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(G1), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n528), .A2(new_n208), .ZN(new_n662));
  OAI22_X1  g0462(.A1(new_n661), .A2(new_n662), .B1(new_n229), .B2(new_n660), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT28), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT29), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n586), .A2(new_n372), .A3(new_n587), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n452), .B1(new_n273), .B2(new_n283), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n569), .A2(new_n574), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n577), .B1(new_n669), .B2(new_n257), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n666), .B1(new_n670), .B2(new_n579), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n612), .A2(new_n671), .A3(new_n557), .A4(new_n589), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(KEYINPUT26), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n559), .A2(new_n605), .A3(new_n606), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(new_n612), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT90), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n673), .A2(KEYINPUT90), .A3(new_n612), .A4(new_n674), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(new_n621), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n665), .B1(new_n679), .B2(new_n647), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n623), .A2(new_n647), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(KEYINPUT29), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n508), .A2(G179), .A3(new_n509), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT88), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n508), .A2(KEYINPUT88), .A3(new_n509), .A4(G179), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n494), .A2(new_n586), .A3(new_n550), .A4(new_n587), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT30), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT30), .ZN(new_n691));
  AOI211_X1 g0491(.A(new_n691), .B(new_n688), .C1(new_n685), .C2(new_n686), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n550), .A2(G179), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n497), .A2(new_n693), .A3(new_n599), .A4(new_n588), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n690), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT31), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n696), .A2(new_n697), .A3(new_n647), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n687), .A2(new_n689), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n691), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n687), .A2(KEYINPUT30), .A3(new_n689), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(new_n694), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(KEYINPUT31), .B1(new_n702), .B2(new_n641), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT89), .B1(new_n698), .B2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n560), .A2(new_n603), .A3(new_n647), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n697), .B1(new_n696), .B2(new_n647), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n702), .A2(KEYINPUT31), .A3(new_n641), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT89), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n704), .A2(new_n705), .A3(new_n709), .ZN(new_n710));
  AOI211_X1 g0510(.A(new_n680), .B(new_n682), .C1(G330), .C2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n664), .B1(new_n711), .B2(G1), .ZN(G364));
  AOI21_X1  g0512(.A(new_n317), .B1(new_n635), .B2(G45), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(new_n659), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n645), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n644), .A2(G330), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n248), .A2(G45), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n306), .A2(new_n658), .ZN(new_n721));
  OAI211_X1 g0521(.A(new_n720), .B(new_n721), .C1(G45), .C2(new_n229), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n272), .A2(new_n658), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G355), .ZN(new_n724));
  OAI211_X1 g0524(.A(new_n722), .B(new_n724), .C1(G116), .C2(new_n232), .ZN(new_n725));
  NOR2_X1   g0525(.A1(G13), .A2(G33), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G20), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n227), .B1(G20), .B2(new_n325), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n725), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n281), .A2(new_n372), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G200), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(new_n601), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n601), .A2(G200), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n372), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n226), .A2(new_n736), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n734), .A2(G326), .B1(G294), .B2(new_n737), .ZN(new_n738));
  XOR2_X1   g0538(.A(new_n738), .B(KEYINPUT92), .Z(new_n739));
  NOR2_X1   g0539(.A1(new_n733), .A2(G190), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(G317), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n741), .B1(KEYINPUT33), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(KEYINPUT33), .B2(new_n742), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n349), .A2(G179), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n226), .A2(new_n601), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT91), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G283), .ZN(new_n749));
  NOR4_X1   g0549(.A1(new_n281), .A2(new_n372), .A3(G190), .A4(G200), .ZN(new_n750));
  NOR4_X1   g0550(.A1(new_n281), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n751));
  AOI22_X1  g0551(.A1(G311), .A2(new_n750), .B1(new_n751), .B2(G329), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n732), .A2(new_n735), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n364), .B1(new_n754), .B2(G322), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n744), .A2(new_n749), .A3(new_n752), .A4(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n745), .A2(G20), .A3(G190), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI211_X1 g0558(.A(new_n739), .B(new_n756), .C1(G303), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n740), .A2(G68), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n751), .A2(G159), .ZN(new_n761));
  INV_X1    g0561(.A(new_n734), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n760), .B1(KEYINPUT32), .B2(new_n761), .C1(new_n762), .C2(new_n202), .ZN(new_n763));
  INV_X1    g0563(.A(new_n750), .ZN(new_n764));
  INV_X1    g0564(.A(new_n253), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n764), .A2(new_n378), .B1(new_n765), .B2(new_n753), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(G87), .B2(new_n758), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n272), .B1(G97), .B2(new_n737), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n767), .B(new_n768), .C1(new_n450), .C2(new_n747), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n763), .B(new_n769), .C1(KEYINPUT32), .C2(new_n761), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n729), .B1(new_n759), .B2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n728), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n731), .B(new_n771), .C1(new_n644), .C2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n719), .B1(new_n716), .B2(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT93), .Z(G396));
  NAND3_X1  g0576(.A1(new_n625), .A2(KEYINPUT95), .A3(new_n641), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n385), .B(new_n388), .C1(new_n387), .C2(new_n647), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT95), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(new_n385), .B2(new_n647), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n777), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n681), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n710), .A2(G330), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n716), .ZN(new_n785));
  INV_X1    g0585(.A(G303), .ZN(new_n786));
  INV_X1    g0586(.A(new_n737), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n762), .A2(new_n786), .B1(new_n514), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n751), .ZN(new_n789));
  INV_X1    g0589(.A(G311), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n789), .A2(new_n790), .B1(new_n479), .B2(new_n753), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n272), .B1(new_n450), .B2(new_n757), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n788), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n748), .A2(G87), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G283), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n740), .A2(KEYINPUT94), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n740), .A2(KEYINPUT94), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n795), .B1(new_n208), .B2(new_n764), .C1(new_n796), .C2(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n306), .B1(new_n787), .B2(new_n765), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(G132), .B2(new_n751), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n331), .B2(new_n747), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT34), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n734), .A2(G137), .B1(G159), .B2(new_n750), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n754), .A2(G143), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n805), .B(new_n806), .C1(new_n391), .C2(new_n741), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n803), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n808), .B1(new_n804), .B2(new_n807), .C1(new_n202), .C2(new_n757), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n800), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n729), .A2(new_n726), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n810), .A2(new_n729), .B1(new_n378), .B2(new_n811), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n812), .B(new_n715), .C1(new_n727), .C2(new_n781), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n785), .A2(new_n813), .ZN(G384));
  NAND3_X1  g0614(.A1(new_n706), .A2(new_n705), .A3(new_n707), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n443), .A2(new_n445), .A3(new_n430), .A4(new_n432), .ZN(new_n816));
  INV_X1    g0616(.A(new_n428), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n641), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n429), .A2(new_n818), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n446), .A2(new_n821), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n815), .B(new_n781), .C1(new_n820), .C2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(KEYINPUT98), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT37), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n353), .A2(new_n355), .A3(new_n345), .ZN(new_n826));
  INV_X1    g0626(.A(new_n639), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n305), .A2(new_n827), .ZN(new_n828));
  AND4_X1   g0628(.A1(new_n825), .A2(new_n328), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n303), .B(new_n257), .C1(new_n342), .C2(new_n264), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n639), .B1(new_n830), .B2(new_n263), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n315), .A2(G179), .A3(new_n320), .A4(new_n323), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n348), .B2(new_n325), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n830), .A2(new_n263), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n831), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n825), .B1(new_n835), .B2(new_n826), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n829), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n831), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n838), .B1(new_n362), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT38), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI211_X1 g0642(.A(KEYINPUT38), .B(new_n838), .C1(new_n362), .C2(new_n839), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n816), .A2(new_n819), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n446), .B2(new_n821), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT98), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n847), .A2(KEYINPUT40), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n846), .A2(new_n781), .A3(new_n815), .A4(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n824), .A2(new_n844), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n828), .B1(new_n631), .B2(new_n358), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n328), .A2(new_n826), .A3(new_n828), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(new_n825), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n841), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n843), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(KEYINPUT40), .B1(new_n856), .B2(new_n823), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n851), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(G330), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n815), .A2(G330), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n447), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT99), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n858), .A2(new_n447), .A3(new_n815), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n443), .A2(new_n445), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n817), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n868), .A2(new_n641), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n631), .B1(new_n627), .B2(new_n628), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n831), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT38), .B1(new_n872), .B2(new_n838), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n841), .B(new_n837), .C1(new_n871), .C2(new_n831), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT39), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT39), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n843), .A2(new_n876), .A3(new_n855), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n870), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n821), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n868), .A2(new_n879), .B1(new_n816), .B2(new_n819), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n623), .A2(new_n647), .A3(new_n781), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n385), .A2(new_n641), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n880), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n884), .A2(new_n844), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n631), .A2(new_n827), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n878), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n447), .B1(new_n682), .B2(new_n680), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n633), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n887), .B(new_n889), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n866), .B(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n317), .B2(new_n635), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n573), .B(KEYINPUT96), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT35), .ZN(new_n894));
  AOI211_X1 g0694(.A(new_n227), .B(new_n281), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n895), .B(G116), .C1(new_n894), .C2(new_n893), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n896), .B(KEYINPUT36), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n378), .B(new_n229), .C1(new_n253), .C2(G68), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(KEYINPUT97), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n331), .A2(G50), .ZN(new_n900));
  OAI211_X1 g0700(.A(G1), .B(new_n261), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n892), .A2(new_n897), .A3(new_n901), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(KEYINPUT100), .ZN(G367));
  OAI22_X1  g0703(.A1(new_n764), .A2(new_n796), .B1(new_n746), .B2(new_n514), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n758), .A2(G116), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT46), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n299), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n790), .B2(new_n762), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n789), .A2(new_n742), .B1(new_n786), .B2(new_n753), .ZN(new_n910));
  NAND2_X1  g0710(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n911));
  OR2_X1    g0711(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n905), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT106), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n909), .A2(new_n910), .A3(new_n914), .ZN(new_n915));
  OAI221_X1 g0715(.A(new_n915), .B1(new_n479), .B2(new_n799), .C1(new_n368), .C2(new_n787), .ZN(new_n916));
  INV_X1    g0716(.A(new_n799), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(G159), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n764), .A2(new_n202), .B1(new_n746), .B2(new_n378), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(G68), .B2(new_n737), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n751), .A2(G137), .B1(new_n253), .B2(new_n758), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT107), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n364), .B1(new_n753), .B2(new_n391), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(G143), .B2(new_n734), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n918), .A2(new_n920), .A3(new_n922), .A4(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n916), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT47), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n716), .B1(new_n927), .B2(new_n729), .ZN(new_n928));
  INV_X1    g0728(.A(new_n721), .ZN(new_n929));
  OAI221_X1 g0729(.A(new_n730), .B1(new_n232), .B2(new_n381), .C1(new_n244), .C2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n620), .B1(new_n549), .B2(new_n647), .ZN(new_n931));
  OR3_X1    g0731(.A1(new_n612), .A2(new_n549), .A3(new_n647), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n928), .B(new_n930), .C1(new_n772), .C2(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n659), .B(KEYINPUT41), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n619), .B1(new_n595), .B2(new_n647), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n605), .A2(new_n641), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n656), .A2(new_n939), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n940), .A2(KEYINPUT104), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(KEYINPUT104), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT45), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n656), .A2(new_n939), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT44), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n941), .A2(KEYINPUT45), .A3(new_n942), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n945), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n653), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n945), .A2(new_n947), .A3(new_n654), .A4(new_n948), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n652), .B(new_n655), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(new_n645), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n950), .A2(new_n711), .A3(new_n951), .A4(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n936), .B1(new_n954), .B2(new_n711), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n937), .A2(new_n938), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n654), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n648), .A2(new_n651), .A3(new_n655), .ZN(new_n959));
  OR3_X1    g0759(.A1(new_n956), .A2(KEYINPUT42), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(KEYINPUT42), .B1(new_n956), .B2(new_n959), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n591), .B1(new_n937), .B2(new_n500), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n647), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT101), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(KEYINPUT101), .B1(new_n961), .B2(new_n963), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n958), .B(new_n960), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT102), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n964), .B(new_n965), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n971), .A2(KEYINPUT102), .A3(new_n958), .A4(new_n960), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n958), .B1(new_n971), .B2(new_n960), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n970), .A2(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n955), .A2(new_n714), .B1(new_n957), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n972), .A2(new_n970), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n973), .A2(new_n974), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n977), .A2(new_n978), .A3(new_n957), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT103), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n975), .A2(KEYINPUT103), .A3(new_n957), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n934), .B1(new_n976), .B2(new_n983), .ZN(G387));
  NAND2_X1  g0784(.A1(new_n953), .A2(new_n714), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n734), .A2(G322), .B1(G303), .B2(new_n750), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n742), .B2(new_n753), .C1(new_n799), .C2(new_n790), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT48), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n796), .B2(new_n787), .C1(new_n479), .C2(new_n757), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT49), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n306), .B1(new_n751), .B2(G326), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n208), .B2(new_n746), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT110), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n989), .A2(new_n990), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n993), .A2(new_n994), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n991), .A2(new_n995), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n754), .A2(G50), .B1(G150), .B2(new_n751), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n999), .B1(new_n331), .B2(new_n764), .C1(new_n378), .C2(new_n757), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n737), .A2(new_n380), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n741), .B2(new_n255), .ZN(new_n1002));
  NOR3_X1   g0802(.A1(new_n1000), .A2(new_n299), .A3(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n514), .B2(new_n747), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n734), .A2(G159), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT109), .Z(new_n1006));
  OAI21_X1  g0806(.A(new_n998), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n1007), .A2(new_n729), .B1(new_n652), .B2(new_n728), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n929), .B1(new_n241), .B2(G45), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(new_n662), .B2(new_n723), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n374), .A2(new_n202), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT50), .Z(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n331), .B2(new_n378), .ZN(new_n1013));
  NOR3_X1   g0813(.A1(new_n1013), .A2(G45), .A3(new_n662), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n1010), .A2(new_n1014), .B1(G107), .B2(new_n232), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n716), .B1(new_n1015), .B2(new_n730), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT108), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1008), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n711), .A2(new_n953), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(KEYINPUT111), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n659), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n711), .A2(new_n953), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n1019), .B2(KEYINPUT111), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n985), .B(new_n1018), .C1(new_n1021), .C2(new_n1023), .ZN(G393));
  NAND2_X1  g0824(.A1(new_n950), .A2(new_n951), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n1022), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1026), .A2(new_n659), .A3(new_n954), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n950), .A2(new_n714), .A3(new_n951), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n917), .A2(G303), .B1(G116), .B2(new_n737), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n479), .B2(new_n764), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT112), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n748), .A2(G107), .B1(G322), .B2(new_n751), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n734), .A2(G317), .B1(new_n754), .B2(G311), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT52), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n364), .B(new_n1036), .C1(G283), .C2(new_n758), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .A4(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G143), .A2(new_n751), .B1(new_n750), .B2(new_n374), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n331), .B2(new_n757), .C1(new_n378), .C2(new_n787), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n734), .A2(G150), .B1(new_n754), .B2(G159), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n299), .B(new_n1040), .C1(KEYINPUT51), .C2(new_n1041), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1041), .A2(KEYINPUT51), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n917), .A2(G50), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1042), .A2(new_n794), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1038), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n716), .B1(new_n1046), .B2(new_n729), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n730), .B1(new_n514), .B2(new_n232), .C1(new_n251), .C2(new_n929), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(new_n772), .C2(new_n939), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1027), .A2(new_n1028), .A3(new_n1049), .ZN(G390));
  NAND3_X1  g0850(.A1(new_n679), .A2(new_n647), .A3(new_n781), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n883), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n846), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n843), .A2(new_n855), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n870), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n875), .B(new_n877), .C1(new_n884), .C2(new_n869), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n710), .A2(G330), .A3(new_n781), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1059), .A2(new_n880), .ZN(new_n1060));
  AND3_X1   g0860(.A1(new_n1057), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n781), .ZN(new_n1062));
  NOR3_X1   g0862(.A1(new_n860), .A2(new_n880), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n1051), .A2(new_n883), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n880), .B1(new_n860), .B2(new_n1062), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1066), .B(new_n1067), .C1(new_n1059), .C2(new_n880), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1063), .B1(new_n1059), .B2(new_n880), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n881), .A2(new_n883), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1068), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT113), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n888), .A2(new_n633), .A3(new_n862), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  AND3_X1   g0875(.A1(new_n1072), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1073), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1065), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1065), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1078), .A2(new_n1080), .A3(new_n659), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT114), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n875), .A2(new_n877), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n869), .B1(new_n1070), .B2(new_n846), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n880), .B1(new_n1051), .B2(new_n883), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n1083), .A2(new_n1084), .B1(new_n1085), .B2(new_n1055), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1063), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1057), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n713), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n875), .A2(new_n726), .A3(new_n877), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n754), .A2(G116), .B1(G294), .B2(new_n751), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1092), .B1(new_n378), .B2(new_n787), .C1(new_n514), .C2(new_n764), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(G87), .B2(new_n758), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n272), .B1(new_n762), .B2(new_n796), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(G68), .B2(new_n748), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1094), .B(new_n1096), .C1(new_n368), .C2(new_n799), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n917), .A2(G137), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n758), .A2(G150), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(KEYINPUT53), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n746), .ZN(new_n1101));
  XOR2_X1   g0901(.A(KEYINPUT54), .B(G143), .Z(new_n1102));
  AOI22_X1  g0902(.A1(new_n1101), .A2(G50), .B1(new_n750), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(G125), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1103), .B1(new_n1104), .B2(new_n789), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(G132), .B2(new_n754), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n787), .A2(new_n286), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n364), .B1(new_n1099), .B2(KEYINPUT53), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1107), .B(new_n1108), .C1(G128), .C2(new_n734), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1098), .A2(new_n1100), .A3(new_n1106), .A4(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1097), .A2(new_n1110), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1111), .A2(new_n729), .B1(new_n255), .B2(new_n811), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1091), .A2(new_n715), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1082), .B1(new_n1090), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n714), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1116), .A2(KEYINPUT114), .A3(new_n1113), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1115), .A2(KEYINPUT115), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(KEYINPUT115), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1081), .B1(new_n1118), .B2(new_n1119), .ZN(G378));
  OAI21_X1  g0920(.A(new_n1075), .B1(new_n1065), .B2(new_n1079), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n859), .A2(new_n887), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1083), .A2(new_n869), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n886), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n884), .A2(new_n844), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(G330), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(new_n851), .B2(new_n857), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT55), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n406), .A2(new_n435), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1131), .A2(new_n394), .A3(new_n827), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n394), .A2(new_n827), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n406), .A2(new_n435), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1130), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1132), .A2(new_n1130), .A3(new_n1134), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1136), .A2(KEYINPUT56), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(KEYINPUT56), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1122), .A2(new_n1129), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1140), .B1(new_n1122), .B2(new_n1129), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1121), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT57), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1140), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n859), .A2(new_n887), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1122), .A2(new_n1129), .A3(new_n1140), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1151), .A2(KEYINPUT57), .A3(new_n1121), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1145), .A2(new_n659), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1140), .A2(new_n726), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n716), .B1(new_n202), .B2(new_n811), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n1155), .A2(KEYINPUT119), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(KEYINPUT119), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n754), .A2(G107), .B1(new_n380), .B2(new_n750), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1101), .A2(new_n253), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1158), .B(new_n1159), .C1(new_n796), .C2(new_n789), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(G68), .B2(new_n737), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n762), .A2(new_n208), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n741), .A2(new_n514), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n299), .B1(new_n378), .B2(new_n757), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1161), .A2(new_n486), .A3(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT116), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT58), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G125), .A2(new_n734), .B1(new_n740), .B2(G132), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n758), .A2(new_n1102), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT117), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n737), .A2(G150), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n754), .A2(G128), .B1(G137), .B2(new_n750), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1171), .A2(new_n1173), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  XOR2_X1   g0976(.A(new_n1176), .B(KEYINPUT59), .Z(new_n1177));
  AOI21_X1  g0977(.A(G41), .B1(new_n751), .B2(G124), .ZN(new_n1178));
  AOI21_X1  g0978(.A(G33), .B1(new_n1101), .B2(G159), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n486), .B1(new_n299), .B2(new_n265), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n202), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1169), .A2(new_n1170), .A3(new_n1180), .A4(new_n1182), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1183), .A2(new_n729), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1157), .B1(new_n1184), .B2(KEYINPUT118), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(KEYINPUT118), .B2(new_n1184), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1154), .A2(new_n1156), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n1151), .B2(new_n714), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1153), .A2(new_n1189), .ZN(G375));
  NAND2_X1  g0990(.A1(new_n811), .A2(new_n331), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n880), .A2(new_n726), .ZN(new_n1192));
  OR2_X1    g0992(.A1(new_n1192), .A2(KEYINPUT120), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(KEYINPUT120), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n799), .A2(new_n208), .B1(new_n368), .B2(new_n764), .ZN(new_n1195));
  OR2_X1    g0995(.A1(new_n1195), .A2(KEYINPUT121), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(KEYINPUT121), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n272), .B1(new_n514), .B2(new_n757), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(G294), .B2(new_n734), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1001), .B1(new_n753), .B2(new_n796), .C1(new_n789), .C2(new_n786), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(G77), .B2(new_n748), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1196), .A2(new_n1197), .A3(new_n1199), .A4(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n757), .A2(new_n286), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n917), .A2(new_n1102), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n754), .A2(G137), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1205), .B(new_n1159), .C1(new_n391), .C2(new_n764), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(G128), .B2(new_n751), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n306), .B1(new_n787), .B2(new_n202), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n734), .B2(G132), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1204), .A2(new_n1207), .A3(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1202), .B1(new_n1203), .B2(new_n1210), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT122), .Z(new_n1212));
  AOI21_X1  g1012(.A(new_n716), .B1(new_n1212), .B2(new_n729), .ZN(new_n1213));
  AND4_X1   g1013(.A1(new_n1191), .A2(new_n1193), .A3(new_n1194), .A4(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n1072), .B2(new_n714), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT123), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1068), .B(new_n1074), .C1(new_n1069), .C2(new_n1071), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1216), .B1(new_n936), .B2(new_n1218), .ZN(G381));
  OAI21_X1  g1019(.A(new_n714), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n1187), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n660), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1221), .B1(new_n1222), .B2(new_n1152), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(G387), .A2(G381), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1081), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1225));
  NOR4_X1   g1025(.A1(G390), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .A4(new_n1226), .ZN(G407));
  NAND3_X1  g1027(.A1(new_n1223), .A2(new_n640), .A3(new_n1225), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(G407), .A2(G213), .A3(new_n1228), .ZN(G409));
  INV_X1    g1029(.A(G390), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(G387), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT126), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  OAI211_X1 g1033(.A(G390), .B(new_n934), .C1(new_n976), .C2(new_n983), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1231), .A2(new_n1234), .ZN(new_n1235));
  XOR2_X1   g1035(.A(G393), .B(G396), .Z(new_n1236));
  AOI21_X1  g1036(.A(new_n1233), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1236), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1238), .A2(new_n1232), .A3(new_n1234), .A4(new_n1231), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT61), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(G213), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1241), .A2(G343), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1153), .A2(G378), .A3(new_n1189), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1121), .B(new_n935), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT124), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1151), .A2(KEYINPUT124), .A3(new_n935), .A4(new_n1121), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1246), .A2(new_n1189), .A3(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1225), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1242), .B1(new_n1243), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT60), .ZN(new_n1251));
  OR2_X1    g1051(.A1(new_n1217), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n660), .B1(new_n1217), .B2(new_n1251), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1252), .A2(new_n1079), .A3(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT125), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1252), .A2(new_n1253), .A3(KEYINPUT125), .A4(new_n1079), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1256), .A2(new_n1216), .A3(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(new_n785), .A3(new_n813), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1256), .A2(new_n1216), .A3(G384), .A4(new_n1257), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1250), .A2(KEYINPUT63), .A3(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT63), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1243), .A2(new_n1249), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1242), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1242), .A2(G2897), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1259), .A2(new_n1260), .A3(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1268), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1264), .B1(new_n1267), .B2(new_n1271), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1267), .A2(new_n1261), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1240), .B(new_n1263), .C1(new_n1272), .C2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT61), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1268), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1261), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1259), .A2(new_n1260), .A3(new_n1268), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1275), .B1(new_n1279), .B2(new_n1250), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n1223), .A2(G378), .B1(new_n1248), .B2(new_n1225), .ZN(new_n1281));
  NOR4_X1   g1081(.A1(new_n1281), .A2(KEYINPUT62), .A3(new_n1242), .A4(new_n1261), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT62), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1283), .B1(new_n1250), .B2(new_n1262), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1280), .A2(new_n1282), .A3(new_n1284), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1274), .B1(new_n1285), .B2(new_n1287), .ZN(G405));
  NAND2_X1  g1088(.A1(new_n1262), .A2(KEYINPUT127), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(G375), .A2(new_n1225), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1289), .A2(new_n1243), .A3(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1243), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(KEYINPUT127), .A3(new_n1262), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1291), .A2(new_n1293), .ZN(new_n1294));
  XNOR2_X1  g1094(.A(new_n1294), .B(new_n1286), .ZN(G402));
endmodule


