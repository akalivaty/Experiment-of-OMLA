//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 1 0 1 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1280, new_n1281, new_n1282, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1288, new_n1289, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(KEYINPUT64), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  OAI21_X1  g0009(.A(new_n208), .B1(new_n209), .B2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G13), .ZN(new_n211));
  NAND4_X1  g0011(.A1(new_n211), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT0), .Z(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G116), .ZN(new_n218));
  INV_X1    g0018(.A(G270), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n202), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  INV_X1    g0023(.A(G97), .ZN(new_n224));
  INV_X1    g0024(.A(G257), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n220), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT1), .ZN(new_n228));
  AND3_X1   g0028(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n229));
  AOI21_X1  g0029(.A(KEYINPUT65), .B1(G1), .B2(G13), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(G20), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(G68), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n222), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n235), .A2(G50), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  AOI211_X1 g0037(.A(new_n215), .B(new_n228), .C1(new_n233), .C2(new_n237), .ZN(G361));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT66), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G232), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT2), .B(G226), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n242), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n248), .B(new_n249), .Z(new_n250));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XOR2_X1   g0051(.A(G107), .B(G116), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n250), .B(new_n253), .Z(G351));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n255), .B1(new_n229), .B2(new_n230), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT3), .B(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G222), .A2(G1698), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G223), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n258), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n257), .B(new_n262), .C1(G77), .C2(new_n258), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT67), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT67), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n267), .B(new_n264), .C1(G41), .C2(G45), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G274), .ZN(new_n270));
  AND2_X1   g0070(.A1(G1), .A2(G13), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n270), .B1(new_n271), .B2(new_n255), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  INV_X1    g0074(.A(G45), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n264), .A2(new_n276), .B1(new_n271), .B2(new_n255), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n263), .B(new_n273), .C1(new_n217), .C2(new_n278), .ZN(new_n279));
  OR2_X1    g0079(.A1(new_n279), .A2(G179), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G1), .A2(G13), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT65), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n264), .A2(G13), .A3(G20), .ZN(new_n284));
  NAND3_X1  g0084(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n283), .A2(new_n284), .A3(new_n285), .A4(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n264), .A2(G20), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(G50), .A3(new_n289), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT8), .B(G58), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n232), .A2(G33), .ZN(new_n292));
  INV_X1    g0092(.A(G150), .ZN(new_n293));
  INV_X1    g0093(.A(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n232), .A2(new_n294), .ZN(new_n295));
  OAI22_X1  g0095(.A1(new_n291), .A2(new_n292), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(G20), .B2(new_n203), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n283), .A2(new_n285), .A3(new_n286), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI221_X1 g0099(.A(new_n290), .B1(G50), .B2(new_n284), .C1(new_n297), .C2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n279), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n280), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n300), .B(KEYINPUT9), .ZN(new_n304));
  INV_X1    g0104(.A(G190), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n279), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(G200), .B2(new_n279), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(KEYINPUT10), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT10), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n310), .B1(new_n304), .B2(new_n307), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n303), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  XOR2_X1   g0112(.A(KEYINPUT15), .B(G87), .Z(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT68), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT15), .B(G87), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT68), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n318), .A2(new_n292), .ZN(new_n319));
  XOR2_X1   g0119(.A(KEYINPUT8), .B(G58), .Z(new_n320));
  NOR2_X1   g0120(.A1(G20), .A2(G33), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n320), .A2(new_n321), .B1(G20), .B2(G77), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n299), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n289), .A2(G77), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n287), .A2(new_n324), .B1(G77), .B2(new_n284), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(G232), .A2(G1698), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n260), .A2(G238), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n258), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n257), .B(new_n329), .C1(G107), .C2(new_n258), .ZN(new_n330));
  INV_X1    g0130(.A(G244), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n330), .B(new_n273), .C1(new_n331), .C2(new_n278), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G200), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n326), .B(new_n333), .C1(new_n305), .C2(new_n332), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(new_n301), .ZN(new_n335));
  OAI221_X1 g0135(.A(new_n335), .B1(G179), .B2(new_n332), .C1(new_n323), .C2(new_n325), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n312), .A2(new_n337), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n321), .A2(G50), .B1(G20), .B2(new_n234), .ZN(new_n339));
  INV_X1    g0139(.A(G77), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n339), .B1(new_n340), .B2(new_n292), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n298), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n342), .B(KEYINPUT11), .ZN(new_n343));
  INV_X1    g0143(.A(new_n284), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n234), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT12), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n288), .A2(G68), .A3(new_n289), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(new_n347), .A3(KEYINPUT70), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(KEYINPUT70), .B1(new_n346), .B2(new_n347), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n277), .A2(G238), .ZN(new_n352));
  NOR2_X1   g0152(.A1(G226), .A2(G1698), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(new_n223), .B2(G1698), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n354), .A2(new_n258), .B1(G33), .B2(G97), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n273), .B(new_n352), .C1(new_n355), .C2(new_n256), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT69), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n223), .A2(G1698), .ZN(new_n358));
  AND2_X1   g0158(.A1(KEYINPUT3), .A2(G33), .ZN(new_n359));
  NOR2_X1   g0159(.A1(KEYINPUT3), .A2(G33), .ZN(new_n360));
  OAI221_X1 g0160(.A(new_n358), .B1(G226), .B2(G1698), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G33), .A2(G97), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n257), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT69), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n364), .A2(new_n365), .A3(new_n273), .A4(new_n352), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n357), .A2(KEYINPUT13), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G179), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n256), .B1(new_n361), .B2(new_n362), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n277), .A2(G238), .ZN(new_n370));
  AND2_X1   g0170(.A1(G33), .A2(G41), .ZN(new_n371));
  OAI21_X1  g0171(.A(G274), .B1(new_n371), .B2(new_n281), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n372), .B1(new_n266), .B2(new_n268), .ZN(new_n373));
  NOR3_X1   g0173(.A1(new_n369), .A2(new_n370), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT13), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n368), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n367), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT71), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT71), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n367), .A2(new_n379), .A3(new_n376), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n356), .A2(KEYINPUT13), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n364), .A2(new_n375), .A3(new_n273), .A4(new_n352), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n301), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  XNOR2_X1  g0184(.A(new_n384), .B(KEYINPUT14), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n351), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n367), .A2(G190), .A3(new_n383), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n382), .A2(new_n383), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(G200), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n387), .A2(new_n351), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n320), .A2(new_n289), .ZN(new_n393));
  OAI22_X1  g0193(.A1(new_n393), .A2(new_n287), .B1(new_n284), .B2(new_n320), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT74), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n394), .B(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n359), .A2(new_n360), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT7), .B1(new_n397), .B2(new_n232), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT3), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n294), .ZN(new_n400));
  NAND2_X1  g0200(.A1(KEYINPUT3), .A2(G33), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n400), .A2(KEYINPUT7), .A3(new_n232), .A4(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(G68), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT73), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G58), .A2(G68), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n232), .B1(new_n235), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(G159), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n295), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n405), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  AND2_X1   g0210(.A1(G58), .A2(G68), .ZN(new_n411));
  OAI21_X1  g0211(.A(G20), .B1(new_n411), .B2(new_n201), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n412), .B(KEYINPUT73), .C1(new_n408), .C2(new_n295), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n404), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT16), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n299), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT72), .B1(new_n359), .B2(new_n360), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT72), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n400), .A2(new_n418), .A3(new_n401), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(new_n419), .A3(new_n232), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT7), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n402), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(G68), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n410), .A2(new_n413), .A3(KEYINPUT16), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n396), .B1(new_n416), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n217), .A2(G1698), .ZN(new_n429));
  OAI221_X1 g0229(.A(new_n429), .B1(G223), .B2(G1698), .C1(new_n359), .C2(new_n360), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G33), .A2(G87), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n257), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n269), .A2(new_n272), .B1(new_n277), .B2(G232), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n301), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n277), .A2(G232), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n273), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n256), .B1(new_n430), .B2(new_n431), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n435), .B1(G179), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT18), .B1(new_n428), .B2(new_n440), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n394), .B(KEYINPUT74), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n410), .A2(new_n413), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n400), .A2(new_n232), .A3(new_n401), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n421), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n234), .B1(new_n445), .B2(new_n402), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n415), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n298), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n425), .B1(new_n423), .B2(G68), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n442), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT18), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n439), .A2(G179), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n439), .B2(new_n301), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n450), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G200), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(new_n437), .B2(new_n438), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n433), .A2(new_n305), .A3(new_n434), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n458), .B(new_n442), .C1(new_n448), .C2(new_n449), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT17), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n234), .B1(new_n422), .B2(new_n402), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n447), .B(new_n298), .C1(new_n462), .C2(new_n425), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n463), .A2(KEYINPUT17), .A3(new_n442), .A4(new_n458), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n441), .A2(new_n454), .A3(new_n461), .A4(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n338), .A2(new_n392), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n275), .A2(G1), .ZN(new_n469));
  AND2_X1   g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  NOR2_X1   g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n271), .A2(new_n255), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(G264), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT83), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT83), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n472), .A2(new_n476), .A3(G264), .A4(new_n473), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g0278(.A(KEYINPUT5), .B(G41), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n272), .A2(new_n469), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G294), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n294), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G250), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n260), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n225), .A2(G1698), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n485), .B(new_n486), .C1(new_n359), .C2(new_n360), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n256), .B1(new_n483), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n478), .A2(G179), .A3(new_n480), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT84), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n488), .B1(new_n475), .B2(new_n477), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT84), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n492), .A2(new_n493), .A3(G179), .A4(new_n480), .ZN(new_n494));
  NOR2_X1   g0294(.A1(G250), .A2(G1698), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n495), .B1(new_n225), .B2(G1698), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n482), .B1(new_n496), .B2(new_n258), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n474), .B(new_n480), .C1(new_n497), .C2(new_n256), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G169), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT82), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT82), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n498), .A2(new_n501), .A3(G169), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n491), .A2(new_n494), .A3(new_n500), .A4(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n232), .B(G87), .C1(new_n359), .C2(new_n360), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT22), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT22), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n258), .A2(new_n506), .A3(new_n232), .A4(G87), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT23), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n232), .B2(G107), .ZN(new_n510));
  INV_X1    g0310(.A(G107), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n511), .A2(KEYINPUT23), .A3(G20), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n294), .A2(new_n218), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n232), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n508), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT24), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(KEYINPUT80), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n516), .B1(new_n505), .B2(new_n507), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT80), .ZN(new_n522));
  OAI21_X1  g0322(.A(KEYINPUT24), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n508), .A2(new_n522), .A3(new_n517), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n520), .B(new_n298), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n264), .A2(G33), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n288), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G107), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT81), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n344), .B(new_n511), .C1(new_n530), .C2(KEYINPUT25), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(KEYINPUT25), .ZN(new_n532));
  XNOR2_X1  g0332(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n525), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n503), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n492), .A2(new_n480), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n455), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(G190), .B2(new_n498), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n518), .A2(KEYINPUT80), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n521), .A2(new_n522), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(KEYINPUT24), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n522), .B1(new_n508), .B2(new_n517), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n299), .B1(new_n544), .B2(new_n519), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n534), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n540), .A2(new_n546), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n537), .A2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT6), .ZN(new_n549));
  AND2_X1   g0349(.A1(G97), .A2(G107), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n549), .B1(new_n550), .B2(new_n205), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n511), .A2(KEYINPUT6), .A3(G97), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n553), .A2(G20), .B1(G77), .B2(new_n321), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n511), .B1(new_n445), .B2(new_n402), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT75), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AOI211_X1 g0357(.A(KEYINPUT75), .B(new_n511), .C1(new_n445), .C2(new_n402), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n298), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT76), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT76), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n561), .B(new_n298), .C1(new_n557), .C2(new_n558), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n284), .A2(G97), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n564), .B1(new_n528), .B2(G97), .ZN(new_n565));
  AND2_X1   g0365(.A1(KEYINPUT4), .A2(G244), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n260), .B(new_n566), .C1(new_n359), .C2(new_n360), .ZN(new_n567));
  NAND2_X1  g0367(.A1(G33), .A2(G283), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n331), .B1(new_n400), .B2(new_n401), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n567), .B(new_n568), .C1(new_n569), .C2(KEYINPUT4), .ZN(new_n570));
  OAI21_X1  g0370(.A(G250), .B1(new_n359), .B2(new_n360), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n260), .B1(new_n571), .B2(KEYINPUT4), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n257), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n472), .A2(new_n372), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n472), .A2(new_n473), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n574), .B1(new_n575), .B2(G257), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT77), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT77), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n573), .A2(new_n579), .A3(new_n576), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(G190), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n577), .A2(G200), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n563), .A2(new_n565), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n562), .ZN(new_n584));
  OAI21_X1  g0384(.A(G107), .B1(new_n398), .B2(new_n403), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT75), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n555), .A2(new_n556), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(new_n587), .A3(new_n554), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n561), .B1(new_n588), .B2(new_n298), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n565), .B1(new_n584), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n577), .A2(G179), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n578), .A2(new_n580), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n591), .B1(new_n592), .B2(new_n301), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n473), .B(G250), .C1(G1), .C2(new_n275), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n272), .A2(new_n469), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(G238), .B(new_n260), .C1(new_n359), .C2(new_n360), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(KEYINPUT78), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT78), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n258), .A2(new_n600), .A3(G238), .A4(new_n260), .ZN(new_n601));
  INV_X1    g0401(.A(new_n514), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n258), .A2(G244), .A3(G1698), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n599), .A2(new_n601), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n597), .B1(new_n604), .B2(new_n257), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(G179), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n301), .B2(new_n605), .ZN(new_n607));
  INV_X1    g0407(.A(new_n318), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n528), .A2(new_n608), .A3(KEYINPUT79), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT79), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n527), .B2(new_n318), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n258), .A2(new_n232), .A3(G68), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT19), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n232), .B1(new_n362), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(G87), .B2(new_n206), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n613), .B1(new_n292), .B2(new_n224), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n612), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n298), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n318), .A2(new_n344), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n609), .A2(new_n611), .A3(new_n618), .A4(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n288), .A2(G87), .A3(new_n526), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n618), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n604), .A2(new_n257), .ZN(new_n623));
  INV_X1    g0423(.A(new_n597), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n622), .B1(new_n625), .B2(G200), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n605), .A2(G190), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n607), .A2(new_n620), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n548), .A2(new_n583), .A3(new_n594), .A4(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n258), .A2(G257), .A3(new_n260), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n258), .A2(G264), .A3(G1698), .ZN(new_n631));
  INV_X1    g0431(.A(G303), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n630), .B(new_n631), .C1(new_n632), .C2(new_n258), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n257), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n472), .A2(new_n473), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n480), .B1(new_n635), .B2(new_n219), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n288), .A2(G116), .A3(new_n526), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n344), .A2(new_n218), .ZN(new_n640));
  AOI21_X1  g0440(.A(G20), .B1(G33), .B2(G283), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n294), .A2(G97), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n641), .A2(new_n642), .B1(G20), .B2(new_n218), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n643), .A2(new_n298), .A3(KEYINPUT20), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT20), .B1(new_n643), .B2(new_n298), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n639), .B(new_n640), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n638), .A2(new_n646), .A3(KEYINPUT21), .A4(G169), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n636), .B1(new_n257), .B2(new_n633), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n648), .A2(new_n646), .A3(G179), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n301), .B1(new_n634), .B2(new_n637), .ZN(new_n651));
  AOI21_X1  g0451(.A(KEYINPUT21), .B1(new_n651), .B2(new_n646), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n648), .A2(G190), .ZN(new_n654));
  INV_X1    g0454(.A(new_n646), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n654), .B(new_n655), .C1(new_n455), .C2(new_n648), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n468), .A2(new_n629), .A3(new_n657), .ZN(G372));
  NAND3_X1  g0458(.A1(new_n628), .A2(new_n590), .A3(new_n593), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n659), .A2(KEYINPUT26), .B1(new_n607), .B2(new_n620), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n594), .A2(new_n583), .A3(new_n628), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n494), .A2(new_n500), .A3(new_n502), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n546), .B1(new_n662), .B2(new_n491), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n651), .A2(new_n646), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT21), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n666), .A2(new_n649), .A3(new_n647), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n547), .B1(new_n663), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT85), .ZN(new_n669));
  INV_X1    g0469(.A(new_n565), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n670), .B1(new_n560), .B2(new_n562), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n573), .A2(new_n579), .A3(new_n576), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n579), .B1(new_n573), .B2(new_n576), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n301), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n591), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n669), .B1(new_n671), .B2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n590), .A2(KEYINPUT85), .A3(new_n593), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(new_n678), .A3(new_n628), .ZN(new_n679));
  OAI221_X1 g0479(.A(new_n660), .B1(new_n661), .B2(new_n668), .C1(KEYINPUT26), .C2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n467), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g0481(.A(new_n681), .B(KEYINPUT86), .Z(new_n682));
  INV_X1    g0482(.A(new_n303), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT14), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n384), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n384), .A2(new_n684), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n367), .A2(new_n379), .A3(new_n376), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n379), .B1(new_n367), .B2(new_n376), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n685), .B(new_n686), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n351), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n391), .B2(new_n336), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n692), .A2(new_n461), .A3(new_n464), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n441), .A2(new_n454), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n309), .A2(new_n311), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n683), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n682), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g0498(.A(new_n698), .B(KEYINPUT87), .Z(G369));
  NAND3_X1  g0499(.A1(new_n264), .A2(new_n232), .A3(G13), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G213), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(G343), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n655), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n667), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n657), .B2(new_n707), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(G330), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n537), .B(new_n547), .C1(new_n546), .C2(new_n706), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n663), .A2(new_n705), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n537), .A2(new_n667), .A3(new_n547), .A4(new_n706), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n663), .A2(new_n706), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n714), .A2(new_n717), .ZN(G399));
  INV_X1    g0518(.A(new_n213), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G41), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n721), .A2(G1), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n723), .B1(new_n237), .B2(new_n720), .ZN(new_n724));
  XNOR2_X1  g0524(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n724), .B(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n648), .A2(new_n605), .A3(G179), .A4(new_n492), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n727), .B1(new_n592), .B2(new_n728), .ZN(new_n729));
  AND4_X1   g0529(.A1(G179), .A2(new_n648), .A3(new_n605), .A4(new_n492), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n672), .A2(new_n673), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(new_n731), .A3(KEYINPUT30), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n648), .A2(G179), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n733), .A2(new_n538), .A3(new_n577), .A4(new_n625), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n729), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n705), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT31), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n705), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n653), .A2(new_n656), .A3(new_n706), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n738), .B(new_n739), .C1(new_n629), .C2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G330), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n680), .A2(new_n706), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT29), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n581), .A2(new_n582), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n590), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n671), .A2(new_n676), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT89), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n537), .A2(new_n653), .B1(new_n540), .B2(new_n546), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n750), .A2(new_n751), .A3(new_n628), .A4(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(KEYINPUT89), .B1(new_n661), .B2(new_n668), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n679), .A2(KEYINPUT26), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT26), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n628), .A2(new_n590), .A3(new_n757), .A4(new_n593), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n607), .A2(new_n620), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  OAI211_X1 g0561(.A(KEYINPUT29), .B(new_n706), .C1(new_n755), .C2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n743), .B1(new_n746), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n726), .B1(new_n763), .B2(G1), .ZN(G364));
  NOR2_X1   g0564(.A1(new_n211), .A2(G20), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n264), .B1(new_n765), .B2(G45), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n720), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n231), .B1(G20), .B2(new_n301), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n770), .A2(KEYINPUT91), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(KEYINPUT91), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n211), .A2(new_n294), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT90), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n213), .A2(new_n258), .ZN(new_n780));
  INV_X1    g0580(.A(G355), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n780), .A2(new_n781), .B1(G116), .B2(new_n213), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n417), .A2(new_n419), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n719), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n785), .B1(new_n275), .B2(new_n237), .ZN(new_n786));
  OR2_X1    g0586(.A1(new_n250), .A2(new_n275), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n782), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n768), .B1(new_n779), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n232), .A2(G179), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G190), .A2(G200), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G159), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT32), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n232), .A2(new_n368), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G200), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n305), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n790), .A2(new_n305), .A3(G200), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n799), .A2(new_n202), .B1(new_n800), .B2(new_n511), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n795), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n796), .A2(G190), .A3(new_n455), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n258), .B1(new_n803), .B2(new_n222), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n305), .A2(G179), .A3(G200), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n232), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n790), .A2(G190), .A3(G200), .ZN(new_n807));
  INV_X1    g0607(.A(G87), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n806), .A2(new_n224), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n796), .A2(new_n791), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n804), .B(new_n809), .C1(G77), .C2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n797), .A2(G190), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n813), .A2(KEYINPUT92), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n813), .A2(KEYINPUT92), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n802), .B(new_n812), .C1(new_n234), .C2(new_n816), .ZN(new_n817));
  XOR2_X1   g0617(.A(KEYINPUT33), .B(G317), .Z(new_n818));
  INV_X1    g0618(.A(G322), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n816), .A2(new_n818), .B1(new_n819), .B2(new_n803), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT93), .ZN(new_n821));
  INV_X1    g0621(.A(G311), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n810), .A2(new_n822), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n258), .B(new_n823), .C1(G329), .C2(new_n793), .ZN(new_n824));
  INV_X1    g0624(.A(new_n806), .ZN(new_n825));
  INV_X1    g0625(.A(new_n800), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n825), .A2(G294), .B1(new_n826), .B2(G283), .ZN(new_n827));
  INV_X1    g0627(.A(new_n807), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n798), .A2(G326), .B1(new_n828), .B2(G303), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n824), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n817), .B1(new_n821), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n789), .B1(new_n831), .B2(new_n773), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n709), .B2(new_n776), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT94), .Z(new_n834));
  INV_X1    g0634(.A(new_n710), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n768), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(G330), .B2(new_n709), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n834), .A2(new_n837), .ZN(G396));
  OAI21_X1  g0638(.A(new_n334), .B1(new_n326), .B2(new_n706), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n336), .ZN(new_n840));
  OR2_X1    g0640(.A1(new_n336), .A2(new_n705), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n744), .A2(new_n842), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n840), .A2(new_n841), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n659), .A2(KEYINPUT26), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n845), .B(new_n759), .C1(new_n661), .C2(new_n668), .ZN(new_n846));
  AND4_X1   g0646(.A1(new_n757), .A2(new_n677), .A3(new_n678), .A4(new_n628), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n706), .B(new_n844), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n768), .B1(new_n849), .B2(new_n742), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n742), .B2(new_n849), .ZN(new_n851));
  INV_X1    g0651(.A(new_n773), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n774), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n768), .B1(new_n853), .B2(G77), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n799), .A2(new_n632), .B1(new_n807), .B2(new_n511), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n806), .A2(new_n224), .B1(new_n800), .B2(new_n808), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n810), .A2(new_n218), .B1(new_n792), .B2(new_n822), .ZN(new_n858));
  INV_X1    g0658(.A(new_n803), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n258), .B(new_n858), .C1(G294), .C2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(G283), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n857), .B(new_n860), .C1(new_n861), .C2(new_n816), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT95), .Z(new_n863));
  AOI22_X1  g0663(.A1(new_n859), .A2(G143), .B1(new_n811), .B2(G159), .ZN(new_n864));
  INV_X1    g0664(.A(G137), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n864), .B1(new_n865), .B2(new_n799), .C1(new_n816), .C2(new_n293), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT34), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n202), .A2(new_n807), .B1(new_n800), .B2(new_n234), .ZN(new_n869));
  INV_X1    g0669(.A(G132), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n783), .B1(new_n870), .B2(new_n792), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n869), .B(new_n871), .C1(G58), .C2(new_n825), .ZN(new_n872));
  INV_X1    g0672(.A(new_n866), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n872), .B1(new_n873), .B2(KEYINPUT34), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n863), .B1(new_n868), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n854), .B1(new_n875), .B2(new_n773), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n844), .B2(new_n774), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n851), .A2(new_n877), .ZN(G384));
  NOR2_X1   g0678(.A1(new_n765), .A2(new_n264), .ZN(new_n879));
  XOR2_X1   g0679(.A(KEYINPUT99), .B(KEYINPUT40), .Z(new_n880));
  OAI21_X1  g0680(.A(new_n705), .B1(new_n349), .B2(new_n350), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT96), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n386), .B2(new_n391), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT96), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n881), .B(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n691), .A2(new_n390), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n741), .A2(new_n844), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n415), .B1(new_n462), .B2(new_n443), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n427), .A2(new_n889), .A3(new_n298), .ZN(new_n890));
  INV_X1    g0690(.A(new_n394), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n703), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n459), .A2(KEYINPUT37), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n890), .A2(new_n891), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n453), .ZN(new_n896));
  INV_X1    g0696(.A(new_n703), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n450), .B1(new_n453), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n459), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT37), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n894), .A2(new_n896), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n465), .A2(new_n892), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT38), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT38), .B1(new_n901), .B2(new_n902), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n880), .B1(new_n888), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n428), .A2(new_n703), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n465), .A2(new_n907), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n440), .A2(new_n703), .B1(new_n463), .B2(new_n442), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT37), .B1(new_n909), .B2(KEYINPUT97), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n899), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n898), .A2(new_n459), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT97), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n900), .B1(new_n898), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n908), .A2(new_n911), .A3(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT38), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT38), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n705), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT31), .B1(new_n735), .B2(new_n705), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n740), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n750), .A2(new_n924), .A3(new_n548), .A4(new_n628), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n842), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n920), .A2(KEYINPUT40), .A3(new_n926), .A4(new_n887), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n906), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n467), .A2(new_n741), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n930), .A2(G330), .A3(new_n931), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n932), .B(KEYINPUT100), .Z(new_n933));
  NAND3_X1  g0733(.A1(new_n746), .A2(new_n467), .A3(new_n762), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n697), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT98), .ZN(new_n936));
  INV_X1    g0736(.A(new_n887), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n848), .B2(new_n841), .ZN(new_n938));
  INV_X1    g0738(.A(new_n905), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT39), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n465), .A2(new_n907), .B1(new_n912), .B2(new_n914), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT38), .B1(new_n942), .B2(new_n911), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n941), .B1(new_n943), .B2(new_n903), .ZN(new_n944));
  INV_X1    g0744(.A(new_n904), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n945), .A2(KEYINPUT39), .A3(new_n919), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n691), .A2(new_n705), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n944), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n694), .A2(new_n897), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n940), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n936), .B(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n879), .B1(new_n933), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n933), .B2(new_n951), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n553), .A2(KEYINPUT35), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n553), .A2(KEYINPUT35), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n954), .A2(G116), .A3(new_n233), .A4(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT36), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n237), .A2(G77), .A3(new_n406), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(G50), .B2(new_n234), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n959), .A2(G1), .A3(new_n211), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n953), .A2(new_n957), .A3(new_n960), .ZN(G367));
  OAI211_X1 g0761(.A(new_n594), .B(new_n583), .C1(new_n671), .C2(new_n706), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n749), .A2(new_n705), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n717), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT45), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(KEYINPUT45), .B1(new_n964), .B2(new_n717), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n715), .A2(new_n716), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n969), .A2(new_n962), .A3(new_n963), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT44), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n970), .A2(new_n971), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n967), .A2(new_n968), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n713), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n714), .B1(new_n972), .B2(new_n973), .C1(new_n967), .C2(new_n968), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n667), .A2(new_n706), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n711), .A2(new_n712), .A3(new_n978), .ZN(new_n979));
  AND3_X1   g0779(.A1(new_n710), .A2(new_n715), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n710), .B1(new_n979), .B2(new_n715), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n763), .B1(new_n977), .B2(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n720), .B(KEYINPUT41), .Z(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n767), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n622), .A2(new_n705), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n759), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n628), .A2(new_n987), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT43), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n990), .A2(KEYINPUT43), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n964), .A2(new_n548), .A3(new_n667), .A4(new_n706), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT42), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n962), .A2(KEYINPUT101), .A3(new_n963), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(KEYINPUT101), .B1(new_n962), .B2(new_n963), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n663), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n705), .B1(new_n1000), .B2(new_n594), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n993), .B(new_n994), .C1(new_n996), .C2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n999), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n537), .B1(new_n1003), .B2(new_n997), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n706), .B1(new_n1004), .B2(new_n749), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT42), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n995), .B(new_n1006), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1005), .A2(new_n1007), .A3(new_n992), .A4(new_n991), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n998), .A2(new_n999), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n714), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1002), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(KEYINPUT103), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT103), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1002), .A2(new_n1008), .A3(new_n1013), .A4(new_n1010), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1010), .B1(new_n1002), .B2(new_n1008), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1016), .A2(KEYINPUT102), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1012), .B(new_n1014), .C1(KEYINPUT102), .C2(new_n1016), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n986), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n768), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n778), .B1(new_n213), .B2(new_n318), .C1(new_n242), .C2(new_n785), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1021), .B1(new_n1022), .B2(KEYINPUT104), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(KEYINPUT104), .B2(new_n1022), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n783), .B1(new_n798), .B2(G311), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n825), .A2(G107), .B1(new_n826), .B2(G97), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(new_n816), .C2(new_n481), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n859), .A2(G303), .B1(new_n793), .B2(G317), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n828), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT46), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n807), .B2(new_n218), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n811), .A2(G283), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1028), .A2(new_n1029), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n816), .A2(new_n408), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(G68), .A2(new_n825), .B1(new_n798), .B2(G143), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n397), .B1(new_n811), .B2(G50), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n859), .A2(G150), .B1(new_n793), .B2(G137), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n828), .A2(G58), .B1(new_n826), .B2(G77), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n1027), .A2(new_n1033), .B1(new_n1034), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT47), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n1042), .A2(new_n773), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1024), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n991), .A2(new_n777), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1020), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(G387));
  INV_X1    g0850(.A(new_n982), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n784), .B1(new_n246), .B2(new_n275), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n722), .B2(new_n780), .ZN(new_n1053));
  OR3_X1    g0853(.A1(new_n291), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1054));
  OAI21_X1  g0854(.A(KEYINPUT50), .B1(new_n291), .B2(G50), .ZN(new_n1055));
  AOI21_X1  g0855(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1054), .A2(new_n722), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n1053), .A2(new_n1057), .B1(new_n511), .B2(new_n719), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n768), .B1(new_n1058), .B2(new_n779), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n783), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n340), .A2(new_n807), .B1(new_n800), .B2(new_n224), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(G150), .C2(new_n793), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT105), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n816), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n320), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n608), .A2(new_n825), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n803), .A2(new_n202), .B1(new_n810), .B2(new_n234), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(G159), .B2(new_n798), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1063), .A2(new_n1065), .A3(new_n1066), .A4(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n859), .A2(G317), .B1(new_n811), .B2(G303), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT106), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1071), .B1(new_n819), .B2(new_n799), .C1(new_n822), .C2(new_n816), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT48), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n806), .A2(new_n861), .B1(new_n807), .B2(new_n481), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1074), .A2(KEYINPUT49), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n783), .B1(G326), .B2(new_n793), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1077), .B(new_n1078), .C1(new_n218), .C2(new_n800), .ZN(new_n1079));
  AOI21_X1  g0879(.A(KEYINPUT49), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1069), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1059), .B1(new_n1081), .B2(new_n773), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n711), .A2(new_n712), .A3(new_n777), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n1051), .A2(new_n767), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n763), .A2(new_n1051), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n720), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n763), .A2(new_n1051), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1084), .B1(new_n1086), .B2(new_n1087), .ZN(G393));
  INV_X1    g0888(.A(KEYINPUT109), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n720), .B1(new_n1085), .B2(new_n977), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n975), .A2(new_n976), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n743), .B(new_n982), .C1(new_n746), .C2(new_n762), .ZN(new_n1092));
  OAI21_X1  g0892(.A(KEYINPUT108), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT108), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1085), .A2(new_n977), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1090), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n253), .A2(new_n784), .B1(G97), .B2(new_n719), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1021), .B1(new_n778), .B2(new_n1097), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n806), .A2(new_n218), .B1(new_n810), .B2(new_n481), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(G317), .A2(new_n798), .B1(new_n859), .B2(G311), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT52), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1099), .B(new_n1101), .C1(G303), .C2(new_n1064), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n397), .B1(new_n792), .B2(new_n819), .C1(new_n511), .C2(new_n800), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(G283), .B2(new_n828), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT107), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n799), .A2(new_n293), .B1(new_n408), .B2(new_n803), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT51), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n793), .A2(G143), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1108), .B(new_n783), .C1(new_n291), .C2(new_n810), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n825), .A2(G77), .B1(new_n826), .B2(G87), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n234), .B2(new_n807), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1109), .B(new_n1111), .C1(new_n1064), .C2(G50), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1102), .A2(new_n1105), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1098), .B1(new_n1113), .B2(new_n852), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n1009), .B2(new_n777), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(new_n1091), .B2(new_n767), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1089), .B1(new_n1096), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n721), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1095), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1094), .B1(new_n1085), .B2(new_n977), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1119), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1122), .A2(KEYINPUT109), .A3(new_n1116), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1118), .A2(new_n1123), .ZN(G390));
  NAND4_X1  g0924(.A1(new_n741), .A2(G330), .A3(new_n887), .A4(new_n844), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n848), .A2(new_n841), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n887), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n947), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n1128), .A2(new_n1129), .B1(new_n944), .B2(new_n946), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT110), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n947), .B(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n920), .A2(new_n1132), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n706), .B(new_n840), .C1(new_n755), .C2(new_n761), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n841), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1133), .B1(new_n1135), .B2(new_n887), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1126), .B1(new_n1130), .B2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1125), .B(KEYINPUT111), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n944), .A2(new_n946), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n938), .B2(new_n947), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n937), .B1(new_n1134), .B2(new_n841), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1138), .B(new_n1140), .C1(new_n1141), .C2(new_n1133), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1137), .A2(new_n767), .A3(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n768), .B1(new_n853), .B2(new_n320), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1064), .A2(G137), .ZN(new_n1145));
  INV_X1    g0945(.A(G125), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n803), .A2(new_n870), .B1(new_n792), .B2(new_n1146), .ZN(new_n1147));
  XOR2_X1   g0947(.A(KEYINPUT54), .B(G143), .Z(new_n1148));
  AOI211_X1 g0948(.A(new_n397), .B(new_n1147), .C1(new_n811), .C2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(G128), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n799), .A2(new_n1150), .B1(new_n800), .B2(new_n202), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G159), .B2(new_n825), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n807), .A2(new_n293), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1145), .A2(new_n1149), .A3(new_n1152), .A4(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n816), .A2(new_n511), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(G77), .A2(new_n825), .B1(new_n798), .B2(G283), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n258), .B1(new_n793), .B2(G294), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n859), .A2(G116), .B1(new_n811), .B2(G97), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n828), .A2(G87), .B1(new_n826), .B2(G68), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1156), .B1(new_n1157), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1144), .B1(new_n1163), .B2(new_n773), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1139), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1164), .B1(new_n1165), .B2(new_n774), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1143), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n741), .A2(G330), .A3(new_n844), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n937), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n1125), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n1127), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT111), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1125), .B(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1169), .A2(new_n841), .A3(new_n1134), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1171), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT112), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n743), .A2(new_n467), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n934), .A2(new_n697), .A3(new_n1177), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n1175), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1176), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT113), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1137), .A2(new_n1142), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1175), .A2(new_n1178), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(KEYINPUT112), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1175), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1186), .A2(new_n1183), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT113), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1184), .A2(new_n1189), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1137), .A2(new_n1142), .A3(new_n1175), .A4(new_n1178), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n720), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1167), .B1(new_n1190), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(G378));
  INV_X1    g0995(.A(KEYINPUT57), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n1191), .A2(new_n1178), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n940), .A2(new_n948), .A3(new_n949), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n300), .A2(new_n897), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n312), .A2(new_n1200), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n303), .B(new_n1199), .C1(new_n309), .C2(new_n311), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1203));
  AND3_X1   g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1203), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  AND4_X1   g1006(.A1(G330), .A2(new_n906), .A3(new_n927), .A4(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(G330), .ZN(new_n1208));
  AND3_X1   g1008(.A1(new_n741), .A2(new_n844), .A3(new_n887), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT40), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n918), .B2(new_n919), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1208), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1206), .B1(new_n1212), .B2(new_n906), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1198), .B1(new_n1207), .B2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n906), .A2(new_n927), .A3(G330), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1206), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1212), .A2(new_n906), .A3(new_n1206), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1217), .A2(new_n950), .A3(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1214), .A2(KEYINPUT117), .A3(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT117), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1198), .B(new_n1221), .C1(new_n1207), .C2(new_n1213), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1196), .B1(new_n1197), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1191), .A2(new_n1178), .ZN(new_n1225));
  OR4_X1    g1025(.A1(KEYINPUT118), .A2(new_n1198), .A3(new_n1207), .A4(new_n1213), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1214), .A2(KEYINPUT118), .A3(new_n1219), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1225), .A2(new_n1226), .A3(KEYINPUT57), .A4(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1224), .A2(new_n720), .A3(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1220), .A2(new_n767), .A3(new_n1222), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n768), .B1(new_n853), .B2(G50), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n826), .A2(G58), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1232), .B1(new_n340), .B2(new_n807), .C1(new_n799), .C2(new_n218), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n803), .A2(new_n511), .B1(new_n792), .B2(new_n861), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1060), .A2(new_n274), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1234), .B(new_n1235), .C1(G68), .C2(new_n825), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n318), .B2(new_n810), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n1233), .B(new_n1237), .C1(G97), .C2(new_n1064), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1238), .A2(KEYINPUT58), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n803), .A2(new_n1150), .B1(new_n810), .B2(new_n865), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(G150), .B2(new_n825), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n798), .A2(G125), .B1(new_n828), .B2(new_n1148), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(new_n816), .C2(new_n870), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1243), .A2(KEYINPUT59), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(KEYINPUT59), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(KEYINPUT115), .B(G124), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n294), .B(new_n274), .C1(new_n792), .C2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G159), .B2(new_n826), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1244), .A2(new_n1245), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1238), .A2(KEYINPUT58), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1235), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1239), .A2(new_n1249), .A3(new_n1250), .A4(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1231), .B1(new_n1252), .B2(new_n773), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n1216), .B2(new_n774), .ZN(new_n1254));
  XOR2_X1   g1054(.A(new_n1254), .B(KEYINPUT116), .Z(new_n1255));
  AND2_X1   g1055(.A1(new_n1230), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1229), .A2(new_n1256), .ZN(G375));
  OAI211_X1 g1057(.A(new_n1181), .B(new_n985), .C1(new_n1175), .C2(new_n1178), .ZN(new_n1258));
  OR2_X1    g1058(.A1(new_n887), .A2(new_n774), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n816), .A2(new_n218), .B1(new_n511), .B2(new_n810), .ZN(new_n1260));
  XOR2_X1   g1060(.A(new_n1260), .B(KEYINPUT120), .Z(new_n1261));
  OAI22_X1  g1061(.A1(new_n340), .A2(new_n800), .B1(new_n807), .B2(new_n224), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(G294), .B2(new_n798), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n397), .B1(new_n792), .B2(new_n632), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(G283), .B2(new_n859), .ZN(new_n1265));
  AND4_X1   g1065(.A1(new_n1066), .A2(new_n1261), .A3(new_n1263), .A4(new_n1265), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(G150), .A2(new_n811), .B1(new_n793), .B2(G128), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n859), .A2(G137), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1267), .A2(new_n783), .A3(new_n1232), .A4(new_n1268), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(G50), .A2(new_n825), .B1(new_n798), .B2(G132), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1270), .B1(new_n408), .B2(new_n807), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n1269), .B(new_n1271), .C1(new_n1064), .C2(new_n1148), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n773), .B1(new_n1266), .B2(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n768), .B1(new_n853), .B2(G68), .ZN(new_n1274));
  XOR2_X1   g1074(.A(new_n1274), .B(KEYINPUT119), .Z(new_n1275));
  NAND2_X1  g1075(.A1(new_n1273), .A2(new_n1275), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1276), .B(KEYINPUT121), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n1175), .A2(new_n767), .B1(new_n1259), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1258), .A2(new_n1278), .ZN(G381));
  NOR4_X1   g1079(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1118), .A2(new_n1123), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1280), .A2(new_n1049), .A3(new_n1281), .A4(new_n1194), .ZN(new_n1282));
  OR2_X1    g1082(.A1(new_n1282), .A2(G375), .ZN(G407));
  INV_X1    g1083(.A(G213), .ZN(new_n1284));
  OR3_X1    g1084(.A1(new_n1284), .A2(KEYINPUT122), .A3(G343), .ZN(new_n1285));
  OAI21_X1  g1085(.A(KEYINPUT122), .B1(new_n1284), .B2(G343), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(new_n1287), .B(KEYINPUT123), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1194), .A2(new_n1288), .ZN(new_n1289));
  OAI211_X1 g1089(.A(G407), .B(G213), .C1(G375), .C2(new_n1289), .ZN(G409));
  OAI21_X1  g1090(.A(new_n1281), .B1(new_n1020), .B2(new_n1048), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n986), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1019), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1292), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1295), .A2(new_n1047), .A3(G390), .ZN(new_n1296));
  XOR2_X1   g1096(.A(G393), .B(G396), .Z(new_n1297));
  AND3_X1   g1097(.A1(new_n1291), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1297), .B1(new_n1291), .B2(new_n1296), .ZN(new_n1299));
  NOR3_X1   g1099(.A1(new_n1298), .A2(new_n1299), .A3(KEYINPUT126), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT126), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1297), .ZN(new_n1302));
  NOR3_X1   g1102(.A1(new_n1281), .A2(new_n1020), .A3(new_n1048), .ZN(new_n1303));
  AOI21_X1  g1103(.A(G390), .B1(new_n1295), .B2(new_n1047), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1302), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1291), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1301), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1300), .A2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1182), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1309));
  AND4_X1   g1109(.A1(new_n1182), .A2(new_n1186), .A3(new_n1183), .A4(new_n1187), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1193), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1226), .A2(new_n767), .A3(new_n1227), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1225), .A2(new_n1222), .A3(new_n1220), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1255), .B(new_n1312), .C1(new_n1313), .C2(new_n984), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1167), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1311), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1316), .B1(G375), .B2(new_n1194), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1175), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1178), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1318), .A2(KEYINPUT60), .A3(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n720), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT60), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1322), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1175), .A2(new_n1178), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1278), .B1(new_n1321), .B2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT124), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n851), .A2(new_n1327), .A3(new_n877), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1327), .B1(new_n851), .B2(new_n877), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1326), .A2(new_n1332), .ZN(new_n1333));
  OAI211_X1 g1133(.A(new_n1278), .B(new_n1328), .C1(new_n1321), .C2(new_n1325), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1317), .A2(new_n1287), .A3(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT62), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1192), .B1(new_n1184), .B2(new_n1189), .ZN(new_n1339));
  OAI211_X1 g1139(.A(new_n1229), .B(new_n1256), .C1(new_n1339), .C2(new_n1167), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1288), .B1(new_n1340), .B2(new_n1316), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1336), .A2(KEYINPUT62), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1342), .ZN(new_n1343));
  AOI22_X1  g1143(.A1(new_n1337), .A2(new_n1338), .B1(new_n1341), .B2(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT61), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT125), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1288), .A2(G2897), .ZN(new_n1347));
  AOI211_X1 g1147(.A(new_n1346), .B(new_n1347), .C1(new_n1333), .C2(new_n1334), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1285), .A2(G2897), .A3(new_n1286), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1278), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1325), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n721), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1350), .B1(new_n1351), .B2(new_n1352), .ZN(new_n1353));
  OAI211_X1 g1153(.A(new_n1334), .B(new_n1349), .C1(new_n1353), .C2(new_n1331), .ZN(new_n1354));
  AND2_X1   g1154(.A1(new_n1354), .A2(new_n1346), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1335), .A2(G2897), .A3(new_n1288), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1348), .B1(new_n1355), .B2(new_n1356), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1345), .B1(new_n1357), .B2(new_n1341), .ZN(new_n1358));
  OAI21_X1  g1158(.A(new_n1308), .B1(new_n1344), .B2(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1317), .A2(new_n1287), .ZN(new_n1360));
  AND2_X1   g1160(.A1(new_n1355), .A2(new_n1356), .ZN(new_n1361));
  OAI21_X1  g1161(.A(new_n1360), .B1(new_n1361), .B2(new_n1348), .ZN(new_n1362));
  INV_X1    g1162(.A(KEYINPUT63), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1337), .A2(new_n1363), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1341), .A2(KEYINPUT63), .A3(new_n1336), .ZN(new_n1365));
  NOR3_X1   g1165(.A1(new_n1298), .A2(new_n1299), .A3(KEYINPUT61), .ZN(new_n1366));
  NAND4_X1  g1166(.A1(new_n1362), .A2(new_n1364), .A3(new_n1365), .A4(new_n1366), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1359), .A2(new_n1367), .ZN(G405));
  NAND3_X1  g1168(.A1(G375), .A2(new_n1194), .A3(new_n1335), .ZN(new_n1369));
  INV_X1    g1169(.A(new_n1369), .ZN(new_n1370));
  AOI21_X1  g1170(.A(new_n1335), .B1(G375), .B2(new_n1194), .ZN(new_n1371));
  OAI211_X1 g1171(.A(KEYINPUT127), .B(new_n1340), .C1(new_n1370), .C2(new_n1371), .ZN(new_n1372));
  NOR2_X1   g1172(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1373));
  INV_X1    g1173(.A(new_n1371), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1340), .A2(KEYINPUT127), .ZN(new_n1375));
  NAND3_X1  g1175(.A1(new_n1374), .A2(new_n1375), .A3(new_n1369), .ZN(new_n1376));
  AND3_X1   g1176(.A1(new_n1372), .A2(new_n1373), .A3(new_n1376), .ZN(new_n1377));
  AOI21_X1  g1177(.A(new_n1373), .B1(new_n1372), .B2(new_n1376), .ZN(new_n1378));
  NOR2_X1   g1178(.A1(new_n1377), .A2(new_n1378), .ZN(G402));
endmodule


