

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760;

  AND2_X1 U367 ( .A1(n348), .A2(n347), .ZN(n641) );
  INV_X1 U368 ( .A(n728), .ZN(n347) );
  INV_X1 U369 ( .A(n638), .ZN(n349) );
  NOR2_X1 U370 ( .A1(n528), .A2(n392), .ZN(n350) );
  OR2_X1 U371 ( .A1(n699), .A2(n698), .ZN(n422) );
  NOR2_X1 U372 ( .A1(n561), .A2(n559), .ZN(n700) );
  XNOR2_X1 U373 ( .A(n609), .B(n586), .ZN(n699) );
  XNOR2_X1 U374 ( .A(n406), .B(G478), .ZN(n560) );
  AND2_X1 U375 ( .A1(n439), .A2(n434), .ZN(n433) );
  XOR2_X1 U376 ( .A(n549), .B(n548), .Z(n638) );
  XNOR2_X1 U377 ( .A(n544), .B(n490), .ZN(n743) );
  XNOR2_X1 U378 ( .A(n451), .B(n450), .ZN(n520) );
  XNOR2_X1 U379 ( .A(n430), .B(G119), .ZN(n451) );
  XOR2_X1 U380 ( .A(G101), .B(KEYINPUT68), .Z(n491) );
  INV_X1 U381 ( .A(KEYINPUT3), .ZN(n430) );
  BUF_X2 U382 ( .A(n479), .Z(n733) );
  XNOR2_X2 U383 ( .A(n395), .B(n603), .ZN(n615) );
  XNOR2_X1 U384 ( .A(n346), .B(n367), .ZN(n423) );
  NAND2_X1 U385 ( .A1(n425), .A2(n396), .ZN(n346) );
  XNOR2_X1 U386 ( .A(n637), .B(n349), .ZN(n348) );
  INV_X1 U387 ( .A(n619), .ZN(n455) );
  XNOR2_X2 U388 ( .A(n449), .B(n448), .ZN(n619) );
  NAND2_X1 U389 ( .A1(n350), .A2(n387), .ZN(n383) );
  XNOR2_X2 U390 ( .A(n351), .B(n618), .ZN(n623) );
  NAND2_X1 U391 ( .A1(n453), .A2(n454), .ZN(n351) );
  OR2_X1 U392 ( .A1(n609), .A2(n599), .ZN(n600) );
  AND2_X2 U393 ( .A1(n371), .A2(n370), .ZN(n369) );
  NAND2_X2 U394 ( .A1(n433), .A2(n382), .ZN(n485) );
  XNOR2_X2 U395 ( .A(n489), .B(n488), .ZN(n544) );
  NOR2_X1 U396 ( .A1(n553), .A2(n685), .ZN(n403) );
  NOR2_X1 U397 ( .A1(n376), .A2(n759), .ZN(n374) );
  XNOR2_X1 U398 ( .A(n403), .B(n402), .ZN(n564) );
  INV_X1 U399 ( .A(KEYINPUT45), .ZN(n448) );
  INV_X1 U400 ( .A(KEYINPUT4), .ZN(n404) );
  XOR2_X1 U401 ( .A(G902), .B(KEYINPUT15), .Z(n617) );
  NOR2_X1 U402 ( .A1(n635), .A2(n728), .ZN(n636) );
  NOR2_X1 U403 ( .A1(n722), .A2(n728), .ZN(n723) );
  NAND2_X1 U404 ( .A1(n378), .A2(n374), .ZN(n449) );
  XNOR2_X1 U405 ( .A(n375), .B(KEYINPUT99), .ZN(n759) );
  NOR2_X1 U406 ( .A1(n557), .A2(n554), .ZN(n569) );
  NOR2_X1 U407 ( .A1(n564), .A2(n572), .ZN(n527) );
  XNOR2_X1 U408 ( .A(n582), .B(KEYINPUT1), .ZN(n553) );
  NOR2_X1 U409 ( .A1(n726), .A2(G902), .ZN(n514) );
  XOR2_X1 U410 ( .A(n719), .B(KEYINPUT59), .Z(n721) );
  XNOR2_X1 U411 ( .A(n409), .B(n461), .ZN(n463) );
  XNOR2_X1 U412 ( .A(n404), .B(KEYINPUT65), .ZN(n487) );
  NAND2_X1 U413 ( .A1(n479), .A2(G224), .ZN(n409) );
  XNOR2_X1 U414 ( .A(G113), .B(KEYINPUT69), .ZN(n450) );
  INV_X1 U415 ( .A(G143), .ZN(n407) );
  XOR2_X1 U416 ( .A(G146), .B(G125), .Z(n499) );
  XOR2_X1 U417 ( .A(G110), .B(G104), .Z(n493) );
  INV_X1 U418 ( .A(n695), .ZN(n352) );
  NOR2_X1 U419 ( .A1(n623), .A2(n676), .ZN(n353) );
  NOR2_X1 U420 ( .A1(n623), .A2(n676), .ZN(n354) );
  INV_X1 U421 ( .A(n387), .ZN(n355) );
  NOR2_X2 U422 ( .A1(n623), .A2(n676), .ZN(n724) );
  NOR2_X2 U423 ( .A1(n630), .A2(G902), .ZN(n498) );
  XNOR2_X2 U424 ( .A(n524), .B(n497), .ZN(n630) );
  INV_X1 U425 ( .A(n452), .ZN(n400) );
  NOR2_X1 U426 ( .A1(n598), .A2(n429), .ZN(n428) );
  XNOR2_X1 U427 ( .A(n441), .B(n363), .ZN(n612) );
  AND2_X1 U428 ( .A1(n591), .A2(n440), .ZN(n412) );
  XNOR2_X1 U429 ( .A(n377), .B(n431), .ZN(n376) );
  INV_X1 U430 ( .A(KEYINPUT98), .ZN(n431) );
  XOR2_X1 U431 ( .A(KEYINPUT80), .B(KEYINPUT8), .Z(n506) );
  INV_X1 U432 ( .A(n538), .ZN(n410) );
  NAND2_X1 U433 ( .A1(n460), .A2(n483), .ZN(n484) );
  NAND2_X1 U434 ( .A1(G898), .A2(n408), .ZN(n483) );
  INV_X1 U435 ( .A(KEYINPUT72), .ZN(n402) );
  XNOR2_X1 U436 ( .A(n503), .B(n358), .ZN(n414) );
  XOR2_X1 U437 ( .A(KEYINPUT79), .B(KEYINPUT24), .Z(n503) );
  INV_X1 U438 ( .A(n585), .ZN(n436) );
  NOR2_X1 U439 ( .A1(n398), .A2(n413), .ZN(n555) );
  INV_X1 U440 ( .A(KEYINPUT22), .ZN(n551) );
  XNOR2_X1 U441 ( .A(n443), .B(n442), .ZN(n589) );
  INV_X1 U442 ( .A(KEYINPUT30), .ZN(n442) );
  NOR2_X1 U443 ( .A1(n638), .A2(G902), .ZN(n406) );
  NOR2_X1 U444 ( .A1(n685), .A2(n582), .ZN(n567) );
  XOR2_X1 U445 ( .A(KEYINPUT6), .B(n588), .Z(n572) );
  BUF_X1 U446 ( .A(n682), .Z(n413) );
  OR2_X1 U447 ( .A1(G902), .A2(G237), .ZN(n474) );
  XNOR2_X1 U448 ( .A(G116), .B(KEYINPUT93), .ZN(n517) );
  NAND2_X1 U449 ( .A1(G237), .A2(G234), .ZN(n478) );
  INV_X1 U450 ( .A(KEYINPUT34), .ZN(n392) );
  AND2_X1 U451 ( .A1(n447), .A2(n446), .ZN(n454) );
  NAND2_X1 U452 ( .A1(n357), .A2(KEYINPUT82), .ZN(n444) );
  INV_X1 U453 ( .A(G134), .ZN(n488) );
  XNOR2_X1 U454 ( .A(G143), .B(G122), .ZN(n529) );
  XOR2_X1 U455 ( .A(G104), .B(G113), .Z(n530) );
  XNOR2_X1 U456 ( .A(KEYINPUT95), .B(KEYINPUT11), .ZN(n531) );
  XOR2_X1 U457 ( .A(KEYINPUT12), .B(KEYINPUT96), .Z(n532) );
  INV_X1 U458 ( .A(KEYINPUT17), .ZN(n461) );
  XNOR2_X1 U459 ( .A(n420), .B(KEYINPUT41), .ZN(n711) );
  NOR2_X1 U460 ( .A1(n422), .A2(n421), .ZN(n420) );
  NOR2_X1 U461 ( .A1(n438), .A2(n484), .ZN(n434) );
  XNOR2_X1 U462 ( .A(n565), .B(KEYINPUT94), .ZN(n391) );
  NAND2_X1 U463 ( .A1(n417), .A2(n416), .ZN(n565) );
  NAND2_X1 U464 ( .A1(n436), .A2(n435), .ZN(n382) );
  NOR2_X1 U465 ( .A1(n698), .A2(n477), .ZN(n435) );
  NAND2_X1 U466 ( .A1(n381), .A2(n580), .ZN(n380) );
  XNOR2_X1 U467 ( .A(n569), .B(KEYINPUT100), .ZN(n381) );
  BUF_X1 U468 ( .A(G953), .Z(n408) );
  XNOR2_X1 U469 ( .A(n397), .B(n508), .ZN(n726) );
  XNOR2_X1 U470 ( .A(n507), .B(n539), .ZN(n397) );
  NOR2_X1 U471 ( .A1(G952), .A2(n733), .ZN(n728) );
  NOR2_X1 U472 ( .A1(n612), .A2(n593), .ZN(n594) );
  XNOR2_X1 U473 ( .A(n415), .B(KEYINPUT36), .ZN(n578) );
  OR2_X1 U474 ( .A1(n604), .A2(n571), .ZN(n415) );
  XNOR2_X1 U475 ( .A(n558), .B(n364), .ZN(n452) );
  XNOR2_X1 U476 ( .A(n419), .B(n418), .ZN(n665) );
  INV_X1 U477 ( .A(KEYINPUT31), .ZN(n418) );
  NOR2_X1 U478 ( .A1(n391), .A2(n563), .ZN(n419) );
  NOR2_X1 U479 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U480 ( .A(KEYINPUT97), .B(n562), .Z(n664) );
  XNOR2_X1 U481 ( .A(n570), .B(KEYINPUT86), .ZN(n405) );
  XNOR2_X1 U482 ( .A(n452), .B(n399), .ZN(G21) );
  INV_X1 U483 ( .A(G119), .ZN(n399) );
  AND2_X1 U484 ( .A1(n400), .A2(KEYINPUT44), .ZN(n356) );
  NAND2_X1 U485 ( .A1(KEYINPUT2), .A2(n617), .ZN(n357) );
  XOR2_X1 U486 ( .A(G140), .B(KEYINPUT23), .Z(n358) );
  OR2_X1 U487 ( .A1(n661), .A2(n664), .ZN(n359) );
  INV_X1 U488 ( .A(n698), .ZN(n476) );
  XOR2_X1 U489 ( .A(n601), .B(KEYINPUT76), .Z(n360) );
  AND2_X1 U490 ( .A1(n401), .A2(n356), .ZN(n361) );
  INV_X1 U491 ( .A(n438), .ZN(n437) );
  NOR2_X1 U492 ( .A1(n476), .A2(KEYINPUT19), .ZN(n438) );
  BUF_X1 U493 ( .A(n588), .Z(n580) );
  INV_X1 U494 ( .A(n580), .ZN(n416) );
  AND2_X1 U495 ( .A1(n439), .A2(n437), .ZN(n362) );
  XOR2_X1 U496 ( .A(KEYINPUT70), .B(KEYINPUT39), .Z(n363) );
  XOR2_X1 U497 ( .A(KEYINPUT77), .B(KEYINPUT32), .Z(n364) );
  XNOR2_X1 U498 ( .A(KEYINPUT35), .B(KEYINPUT75), .ZN(n365) );
  AND2_X1 U499 ( .A1(n575), .A2(n432), .ZN(n366) );
  XOR2_X1 U500 ( .A(KEYINPUT46), .B(KEYINPUT64), .Z(n367) );
  INV_X1 U501 ( .A(KEYINPUT82), .ZN(n457) );
  AND2_X1 U502 ( .A1(n357), .A2(n617), .ZN(n368) );
  NAND2_X1 U503 ( .A1(n401), .A2(n400), .ZN(n373) );
  NAND2_X1 U504 ( .A1(n372), .A2(n369), .ZN(n378) );
  NAND2_X1 U505 ( .A1(n379), .A2(n366), .ZN(n370) );
  NAND2_X1 U506 ( .A1(n373), .A2(n432), .ZN(n371) );
  NAND2_X1 U507 ( .A1(n361), .A2(n654), .ZN(n372) );
  NAND2_X1 U508 ( .A1(n379), .A2(n575), .ZN(n654) );
  NAND2_X1 U509 ( .A1(n405), .A2(n413), .ZN(n375) );
  NAND2_X1 U510 ( .A1(n388), .A2(n359), .ZN(n377) );
  XNOR2_X1 U511 ( .A(n380), .B(KEYINPUT67), .ZN(n379) );
  NAND2_X1 U512 ( .A1(n362), .A2(n382), .ZN(n596) );
  NAND2_X1 U513 ( .A1(n385), .A2(n383), .ZN(n394) );
  NAND2_X1 U514 ( .A1(n386), .A2(n392), .ZN(n385) );
  NAND2_X1 U515 ( .A1(n352), .A2(n566), .ZN(n386) );
  INV_X1 U516 ( .A(n695), .ZN(n387) );
  NAND2_X1 U517 ( .A1(n390), .A2(n389), .ZN(n388) );
  INV_X1 U518 ( .A(n649), .ZN(n389) );
  INV_X1 U519 ( .A(n665), .ZN(n390) );
  NAND2_X1 U520 ( .A1(n691), .A2(n391), .ZN(n692) );
  XNOR2_X2 U521 ( .A(n393), .B(n365), .ZN(n401) );
  NAND2_X1 U522 ( .A1(n394), .A2(n360), .ZN(n393) );
  NAND2_X1 U523 ( .A1(n423), .A2(n426), .ZN(n395) );
  INV_X1 U524 ( .A(n757), .ZN(n396) );
  XNOR2_X1 U525 ( .A(n594), .B(KEYINPUT40), .ZN(n757) );
  NAND2_X1 U526 ( .A1(n585), .A2(n477), .ZN(n439) );
  NOR2_X1 U527 ( .A1(n578), .A2(n398), .ZN(n668) );
  XNOR2_X1 U528 ( .A(n684), .B(KEYINPUT88), .ZN(n398) );
  XNOR2_X1 U529 ( .A(n401), .B(G122), .ZN(G24) );
  XNOR2_X2 U530 ( .A(n498), .B(G469), .ZN(n582) );
  INV_X1 U531 ( .A(n756), .ZN(n429) );
  XNOR2_X1 U532 ( .A(n602), .B(KEYINPUT103), .ZN(n756) );
  AND2_X1 U533 ( .A1(n427), .A2(n428), .ZN(n426) );
  NOR2_X1 U534 ( .A1(n711), .A2(n595), .ZN(n587) );
  XNOR2_X2 U535 ( .A(n407), .B(G128), .ZN(n489) );
  XNOR2_X1 U536 ( .A(n493), .B(n494), .ZN(n411) );
  XNOR2_X1 U537 ( .A(n411), .B(n410), .ZN(n495) );
  NAND2_X1 U538 ( .A1(n412), .A2(n592), .ZN(n441) );
  XNOR2_X1 U539 ( .A(n414), .B(n504), .ZN(n508) );
  NOR2_X2 U540 ( .A1(n590), .A2(n589), .ZN(n592) );
  XNOR2_X2 U541 ( .A(n743), .B(n492), .ZN(n524) );
  NOR2_X1 U542 ( .A1(n588), .A2(n698), .ZN(n443) );
  NAND2_X1 U543 ( .A1(n751), .A2(n368), .ZN(n445) );
  NAND2_X1 U544 ( .A1(n619), .A2(n457), .ZN(n447) );
  INV_X1 U545 ( .A(n564), .ZN(n417) );
  INV_X1 U546 ( .A(n560), .ZN(n559) );
  NAND2_X1 U547 ( .A1(n751), .A2(n617), .ZN(n616) );
  INV_X1 U548 ( .A(n422), .ZN(n696) );
  INV_X1 U549 ( .A(n700), .ZN(n421) );
  INV_X1 U550 ( .A(n758), .ZN(n425) );
  XNOR2_X1 U551 ( .A(n668), .B(KEYINPUT85), .ZN(n427) );
  INV_X1 U552 ( .A(KEYINPUT44), .ZN(n432) );
  NAND2_X1 U553 ( .A1(n436), .A2(n476), .ZN(n571) );
  NOR2_X2 U554 ( .A1(n622), .A2(n621), .ZN(n676) );
  NAND2_X1 U555 ( .A1(n456), .A2(n455), .ZN(n453) );
  NAND2_X1 U556 ( .A1(n592), .A2(n591), .ZN(n599) );
  INV_X1 U557 ( .A(n699), .ZN(n440) );
  XNOR2_X2 U558 ( .A(n525), .B(G472), .ZN(n588) );
  NAND2_X1 U559 ( .A1(n445), .A2(n444), .ZN(n446) );
  NOR2_X1 U560 ( .A1(n616), .A2(n457), .ZN(n456) );
  INV_X2 U561 ( .A(G953), .ZN(n479) );
  AND2_X1 U562 ( .A1(n572), .A2(n569), .ZN(n570) );
  XNOR2_X2 U563 ( .A(n514), .B(n513), .ZN(n682) );
  XNOR2_X1 U564 ( .A(KEYINPUT104), .B(KEYINPUT62), .ZN(n459) );
  AND2_X1 U565 ( .A1(n680), .A2(n482), .ZN(n460) );
  XNOR2_X1 U566 ( .A(n463), .B(n462), .ZN(n465) );
  XNOR2_X1 U567 ( .A(n491), .B(G146), .ZN(n492) );
  INV_X1 U568 ( .A(KEYINPUT19), .ZN(n477) );
  XNOR2_X1 U569 ( .A(n642), .B(n459), .ZN(n643) );
  XOR2_X1 U570 ( .A(KEYINPUT74), .B(KEYINPUT18), .Z(n462) );
  XNOR2_X1 U571 ( .A(n491), .B(n499), .ZN(n464) );
  XNOR2_X1 U572 ( .A(n465), .B(n464), .ZN(n467) );
  XOR2_X1 U573 ( .A(n489), .B(n487), .Z(n466) );
  XNOR2_X1 U574 ( .A(n467), .B(n466), .ZN(n471) );
  XOR2_X1 U575 ( .A(n493), .B(KEYINPUT16), .Z(n470) );
  XNOR2_X1 U576 ( .A(G116), .B(G107), .ZN(n468) );
  XNOR2_X1 U577 ( .A(n468), .B(G122), .ZN(n543) );
  XNOR2_X1 U578 ( .A(n520), .B(n543), .ZN(n469) );
  XNOR2_X1 U579 ( .A(n470), .B(n469), .ZN(n734) );
  XNOR2_X1 U580 ( .A(n734), .B(n471), .ZN(n625) );
  OR2_X2 U581 ( .A1(n625), .A2(n617), .ZN(n473) );
  NAND2_X1 U582 ( .A1(G210), .A2(n474), .ZN(n472) );
  XNOR2_X2 U583 ( .A(n473), .B(n472), .ZN(n585) );
  NAND2_X1 U584 ( .A1(G214), .A2(n474), .ZN(n475) );
  XNOR2_X1 U585 ( .A(KEYINPUT89), .B(n475), .ZN(n698) );
  XNOR2_X1 U586 ( .A(n478), .B(KEYINPUT14), .ZN(n680) );
  NOR2_X1 U587 ( .A1(G902), .A2(n733), .ZN(n481) );
  NOR2_X1 U588 ( .A1(n408), .A2(G952), .ZN(n480) );
  NOR2_X1 U589 ( .A1(n481), .A2(n480), .ZN(n482) );
  XNOR2_X2 U590 ( .A(n485), .B(KEYINPUT0), .ZN(n563) );
  INV_X1 U591 ( .A(KEYINPUT90), .ZN(n486) );
  XNOR2_X1 U592 ( .A(n563), .B(n486), .ZN(n566) );
  INV_X1 U593 ( .A(n566), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n487), .B(G137), .ZN(n490) );
  XNOR2_X1 U595 ( .A(G107), .B(KEYINPUT91), .ZN(n496) );
  XOR2_X1 U596 ( .A(G140), .B(G131), .Z(n538) );
  NAND2_X1 U597 ( .A1(G227), .A2(n733), .ZN(n494) );
  XNOR2_X1 U598 ( .A(n496), .B(n495), .ZN(n497) );
  INV_X1 U599 ( .A(n499), .ZN(n500) );
  XNOR2_X1 U600 ( .A(KEYINPUT10), .B(n500), .ZN(n539) );
  XOR2_X1 U601 ( .A(G110), .B(G119), .Z(n502) );
  XNOR2_X1 U602 ( .A(G128), .B(G137), .ZN(n501) );
  XNOR2_X1 U603 ( .A(n502), .B(n501), .ZN(n504) );
  NAND2_X1 U604 ( .A1(G234), .A2(n479), .ZN(n505) );
  XNOR2_X1 U605 ( .A(n505), .B(n506), .ZN(n545) );
  NAND2_X1 U606 ( .A1(G221), .A2(n545), .ZN(n507) );
  XOR2_X1 U607 ( .A(KEYINPUT25), .B(KEYINPUT73), .Z(n512) );
  INV_X1 U608 ( .A(n617), .ZN(n509) );
  NAND2_X1 U609 ( .A1(n509), .A2(G234), .ZN(n510) );
  XNOR2_X1 U610 ( .A(n510), .B(KEYINPUT20), .ZN(n515) );
  NAND2_X1 U611 ( .A1(n515), .A2(G217), .ZN(n511) );
  XNOR2_X1 U612 ( .A(n512), .B(n511), .ZN(n513) );
  NAND2_X1 U613 ( .A1(G221), .A2(n515), .ZN(n516) );
  XOR2_X1 U614 ( .A(KEYINPUT21), .B(n516), .Z(n681) );
  NAND2_X1 U615 ( .A1(n682), .A2(n681), .ZN(n685) );
  XOR2_X1 U616 ( .A(G131), .B(KEYINPUT5), .Z(n518) );
  XNOR2_X1 U617 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U618 ( .A(n520), .B(n519), .Z(n522) );
  NOR2_X1 U619 ( .A1(n408), .A2(G237), .ZN(n535) );
  NAND2_X1 U620 ( .A1(n535), .A2(G210), .ZN(n521) );
  XNOR2_X1 U621 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U622 ( .A(n524), .B(n523), .ZN(n642) );
  NOR2_X1 U623 ( .A1(n642), .A2(G902), .ZN(n525) );
  XOR2_X1 U624 ( .A(KEYINPUT87), .B(KEYINPUT33), .Z(n526) );
  XNOR2_X1 U625 ( .A(n527), .B(n526), .ZN(n695) );
  XNOR2_X1 U626 ( .A(KEYINPUT13), .B(G475), .ZN(n542) );
  XNOR2_X1 U627 ( .A(n530), .B(n529), .ZN(n534) );
  XNOR2_X1 U628 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U629 ( .A(n534), .B(n533), .Z(n537) );
  NAND2_X1 U630 ( .A1(G214), .A2(n535), .ZN(n536) );
  XNOR2_X1 U631 ( .A(n537), .B(n536), .ZN(n540) );
  XNOR2_X1 U632 ( .A(n539), .B(n538), .ZN(n746) );
  XNOR2_X1 U633 ( .A(n540), .B(n746), .ZN(n719) );
  NOR2_X1 U634 ( .A1(G902), .A2(n719), .ZN(n541) );
  XNOR2_X1 U635 ( .A(n542), .B(n541), .ZN(n561) );
  XNOR2_X1 U636 ( .A(n544), .B(n543), .ZN(n549) );
  XOR2_X1 U637 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n547) );
  NAND2_X1 U638 ( .A1(n545), .A2(G217), .ZN(n546) );
  XNOR2_X1 U639 ( .A(n547), .B(n546), .ZN(n548) );
  NAND2_X1 U640 ( .A1(n561), .A2(n559), .ZN(n601) );
  NAND2_X1 U641 ( .A1(n700), .A2(n681), .ZN(n550) );
  NOR2_X1 U642 ( .A1(n563), .A2(n550), .ZN(n552) );
  XNOR2_X1 U643 ( .A(n552), .B(n551), .ZN(n557) );
  BUF_X1 U644 ( .A(n553), .Z(n684) );
  INV_X1 U645 ( .A(n684), .ZN(n554) );
  INV_X1 U646 ( .A(n682), .ZN(n575) );
  NAND2_X1 U647 ( .A1(n555), .A2(n572), .ZN(n556) );
  NOR2_X1 U648 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U649 ( .A1(n560), .A2(n561), .ZN(n593) );
  INV_X1 U650 ( .A(n593), .ZN(n661) );
  NOR2_X1 U651 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U652 ( .A(n567), .B(KEYINPUT92), .ZN(n591) );
  NAND2_X1 U653 ( .A1(n566), .A2(n591), .ZN(n568) );
  NOR2_X1 U654 ( .A1(n416), .A2(n568), .ZN(n649) );
  INV_X1 U655 ( .A(n572), .ZN(n577) );
  INV_X1 U656 ( .A(n681), .ZN(n573) );
  NAND2_X1 U657 ( .A1(n408), .A2(G900), .ZN(n748) );
  NAND2_X1 U658 ( .A1(n460), .A2(n748), .ZN(n590) );
  NOR2_X1 U659 ( .A1(n573), .A2(n590), .ZN(n574) );
  NAND2_X1 U660 ( .A1(n575), .A2(n574), .ZN(n579) );
  NOR2_X1 U661 ( .A1(n593), .A2(n579), .ZN(n576) );
  NAND2_X1 U662 ( .A1(n577), .A2(n576), .ZN(n604) );
  NOR2_X1 U663 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U664 ( .A(KEYINPUT28), .B(n581), .ZN(n584) );
  INV_X1 U665 ( .A(n582), .ZN(n583) );
  NAND2_X1 U666 ( .A1(n584), .A2(n583), .ZN(n595) );
  XNOR2_X1 U667 ( .A(KEYINPUT38), .B(KEYINPUT71), .ZN(n586) );
  BUF_X2 U668 ( .A(n585), .Z(n609) );
  XNOR2_X1 U669 ( .A(n587), .B(KEYINPUT42), .ZN(n758) );
  NOR2_X1 U670 ( .A1(n596), .A2(n595), .ZN(n658) );
  NAND2_X1 U671 ( .A1(n658), .A2(n359), .ZN(n597) );
  XNOR2_X1 U672 ( .A(KEYINPUT47), .B(n597), .ZN(n598) );
  XOR2_X1 U673 ( .A(KEYINPUT84), .B(KEYINPUT48), .Z(n603) );
  NOR2_X1 U674 ( .A1(n698), .A2(n604), .ZN(n605) );
  NAND2_X1 U675 ( .A1(n605), .A2(n684), .ZN(n608) );
  XOR2_X1 U676 ( .A(KEYINPUT43), .B(KEYINPUT101), .Z(n606) );
  XNOR2_X1 U677 ( .A(KEYINPUT102), .B(n606), .ZN(n607) );
  XNOR2_X1 U678 ( .A(n608), .B(n607), .ZN(n610) );
  NAND2_X1 U679 ( .A1(n610), .A2(n609), .ZN(n672) );
  INV_X1 U680 ( .A(n664), .ZN(n611) );
  NOR2_X1 U681 ( .A1(n612), .A2(n611), .ZN(n670) );
  INV_X1 U682 ( .A(n670), .ZN(n613) );
  AND2_X1 U683 ( .A1(n672), .A2(n613), .ZN(n614) );
  AND2_X2 U684 ( .A1(n615), .A2(n614), .ZN(n751) );
  INV_X1 U685 ( .A(KEYINPUT66), .ZN(n618) );
  INV_X1 U686 ( .A(n455), .ZN(n622) );
  NAND2_X1 U687 ( .A1(n751), .A2(KEYINPUT2), .ZN(n620) );
  XOR2_X1 U688 ( .A(KEYINPUT83), .B(n620), .Z(n621) );
  NAND2_X1 U689 ( .A1(n354), .A2(G210), .ZN(n627) );
  XOR2_X1 U690 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n624) );
  XNOR2_X1 U691 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U692 ( .A(n627), .B(n626), .ZN(n628) );
  NOR2_X2 U693 ( .A1(n628), .A2(n728), .ZN(n629) );
  XNOR2_X1 U694 ( .A(n629), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U695 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n632) );
  XNOR2_X1 U696 ( .A(n630), .B(KEYINPUT57), .ZN(n631) );
  XNOR2_X1 U697 ( .A(n632), .B(n631), .ZN(n634) );
  NAND2_X1 U698 ( .A1(n724), .A2(G469), .ZN(n633) );
  XNOR2_X1 U699 ( .A(n634), .B(n633), .ZN(n635) );
  XNOR2_X1 U700 ( .A(n636), .B(KEYINPUT120), .ZN(G54) );
  NAND2_X1 U701 ( .A1(n353), .A2(G478), .ZN(n637) );
  INV_X1 U702 ( .A(KEYINPUT121), .ZN(n640) );
  XNOR2_X1 U703 ( .A(n641), .B(n640), .ZN(G63) );
  NAND2_X1 U704 ( .A1(n354), .A2(G472), .ZN(n644) );
  XNOR2_X1 U705 ( .A(n644), .B(n643), .ZN(n645) );
  NOR2_X2 U706 ( .A1(n645), .A2(n728), .ZN(n647) );
  XNOR2_X1 U707 ( .A(KEYINPUT63), .B(KEYINPUT105), .ZN(n646) );
  XNOR2_X1 U708 ( .A(n647), .B(n646), .ZN(G57) );
  NAND2_X1 U709 ( .A1(n649), .A2(n661), .ZN(n648) );
  XNOR2_X1 U710 ( .A(n648), .B(G104), .ZN(G6) );
  XOR2_X1 U711 ( .A(KEYINPUT26), .B(KEYINPUT107), .Z(n651) );
  NAND2_X1 U712 ( .A1(n649), .A2(n664), .ZN(n650) );
  XNOR2_X1 U713 ( .A(n651), .B(n650), .ZN(n653) );
  XOR2_X1 U714 ( .A(G107), .B(KEYINPUT27), .Z(n652) );
  XNOR2_X1 U715 ( .A(n653), .B(n652), .ZN(G9) );
  XNOR2_X1 U716 ( .A(n654), .B(G110), .ZN(G12) );
  XOR2_X1 U717 ( .A(KEYINPUT108), .B(KEYINPUT29), .Z(n656) );
  NAND2_X1 U718 ( .A1(n658), .A2(n664), .ZN(n655) );
  XNOR2_X1 U719 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U720 ( .A(G128), .B(n657), .ZN(G30) );
  XOR2_X1 U721 ( .A(G146), .B(KEYINPUT109), .Z(n660) );
  NAND2_X1 U722 ( .A1(n658), .A2(n661), .ZN(n659) );
  XNOR2_X1 U723 ( .A(n660), .B(n659), .ZN(G48) );
  NAND2_X1 U724 ( .A1(n665), .A2(n661), .ZN(n662) );
  XNOR2_X1 U725 ( .A(n662), .B(KEYINPUT110), .ZN(n663) );
  XNOR2_X1 U726 ( .A(G113), .B(n663), .ZN(G15) );
  XOR2_X1 U727 ( .A(G116), .B(KEYINPUT111), .Z(n667) );
  NAND2_X1 U728 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U729 ( .A(n667), .B(n666), .ZN(G18) );
  XNOR2_X1 U730 ( .A(G125), .B(n668), .ZN(n669) );
  XNOR2_X1 U731 ( .A(n669), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U732 ( .A(G134), .B(n670), .Z(n671) );
  XNOR2_X1 U733 ( .A(KEYINPUT112), .B(n671), .ZN(G36) );
  XNOR2_X1 U734 ( .A(G140), .B(n672), .ZN(G42) );
  XNOR2_X1 U735 ( .A(KEYINPUT2), .B(KEYINPUT78), .ZN(n673) );
  OR2_X1 U736 ( .A1(n751), .A2(n673), .ZN(n678) );
  NOR2_X1 U737 ( .A1(n455), .A2(n673), .ZN(n674) );
  XOR2_X1 U738 ( .A(KEYINPUT81), .B(n674), .Z(n675) );
  NOR2_X1 U739 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U740 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U741 ( .A1(n679), .A2(n733), .ZN(n717) );
  NAND2_X1 U742 ( .A1(G952), .A2(n680), .ZN(n710) );
  XNOR2_X1 U743 ( .A(KEYINPUT51), .B(KEYINPUT114), .ZN(n693) );
  NOR2_X1 U744 ( .A1(n413), .A2(n681), .ZN(n683) );
  XNOR2_X1 U745 ( .A(KEYINPUT49), .B(n683), .ZN(n690) );
  NAND2_X1 U746 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U747 ( .A(n686), .B(KEYINPUT113), .ZN(n687) );
  XNOR2_X1 U748 ( .A(n687), .B(KEYINPUT50), .ZN(n688) );
  NOR2_X1 U749 ( .A1(n416), .A2(n688), .ZN(n689) );
  NAND2_X1 U750 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U751 ( .A(n693), .B(n692), .ZN(n694) );
  NOR2_X1 U752 ( .A1(n711), .A2(n694), .ZN(n706) );
  NAND2_X1 U753 ( .A1(n696), .A2(n359), .ZN(n697) );
  XNOR2_X1 U754 ( .A(KEYINPUT115), .B(n697), .ZN(n703) );
  NAND2_X1 U755 ( .A1(n699), .A2(n698), .ZN(n701) );
  AND2_X1 U756 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U757 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U758 ( .A1(n355), .A2(n704), .ZN(n705) );
  NOR2_X1 U759 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U760 ( .A(KEYINPUT52), .B(n707), .ZN(n708) );
  XNOR2_X1 U761 ( .A(KEYINPUT116), .B(n708), .ZN(n709) );
  NOR2_X1 U762 ( .A1(n710), .A2(n709), .ZN(n714) );
  NOR2_X1 U763 ( .A1(n355), .A2(n711), .ZN(n712) );
  XOR2_X1 U764 ( .A(KEYINPUT117), .B(n712), .Z(n713) );
  NOR2_X1 U765 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U766 ( .A(KEYINPUT118), .B(n715), .Z(n716) );
  NOR2_X1 U767 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U768 ( .A(KEYINPUT53), .B(n718), .ZN(G75) );
  NAND2_X1 U769 ( .A1(n724), .A2(G475), .ZN(n720) );
  XNOR2_X1 U770 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X1 U771 ( .A(n723), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U772 ( .A1(G217), .A2(n353), .ZN(n725) );
  XNOR2_X1 U773 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U774 ( .A1(n728), .A2(n727), .ZN(G66) );
  NAND2_X1 U775 ( .A1(n733), .A2(n455), .ZN(n732) );
  NAND2_X1 U776 ( .A1(n408), .A2(G224), .ZN(n729) );
  XNOR2_X1 U777 ( .A(KEYINPUT61), .B(n729), .ZN(n730) );
  NAND2_X1 U778 ( .A1(n730), .A2(G898), .ZN(n731) );
  NAND2_X1 U779 ( .A1(n732), .A2(n731), .ZN(n742) );
  NOR2_X1 U780 ( .A1(G898), .A2(n733), .ZN(n738) );
  BUF_X1 U781 ( .A(n734), .Z(n735) );
  XOR2_X1 U782 ( .A(G101), .B(n735), .Z(n736) );
  XNOR2_X1 U783 ( .A(KEYINPUT123), .B(n736), .ZN(n737) );
  NOR2_X1 U784 ( .A1(n738), .A2(n737), .ZN(n740) );
  XNOR2_X1 U785 ( .A(KEYINPUT122), .B(KEYINPUT124), .ZN(n739) );
  XNOR2_X1 U786 ( .A(n740), .B(n739), .ZN(n741) );
  XNOR2_X1 U787 ( .A(n742), .B(n741), .ZN(G69) );
  BUF_X1 U788 ( .A(n743), .Z(n744) );
  XOR2_X1 U789 ( .A(n744), .B(KEYINPUT91), .Z(n745) );
  XNOR2_X1 U790 ( .A(n746), .B(n745), .ZN(n749) );
  XOR2_X1 U791 ( .A(G227), .B(n749), .Z(n747) );
  NOR2_X1 U792 ( .A1(n748), .A2(n747), .ZN(n754) );
  XNOR2_X1 U793 ( .A(KEYINPUT125), .B(n749), .ZN(n750) );
  XNOR2_X1 U794 ( .A(n751), .B(n750), .ZN(n752) );
  NOR2_X1 U795 ( .A1(n408), .A2(n752), .ZN(n753) );
  NOR2_X1 U796 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U797 ( .A(KEYINPUT126), .B(n755), .ZN(G72) );
  XNOR2_X1 U798 ( .A(G143), .B(n756), .ZN(G45) );
  XOR2_X1 U799 ( .A(n757), .B(G131), .Z(G33) );
  XOR2_X1 U800 ( .A(n758), .B(G137), .Z(G39) );
  XOR2_X1 U801 ( .A(G101), .B(n759), .Z(n760) );
  XNOR2_X1 U802 ( .A(KEYINPUT106), .B(n760), .ZN(G3) );
endmodule

