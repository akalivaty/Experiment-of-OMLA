//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1321,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1387, new_n1388, new_n1389,
    new_n1390, new_n1391, new_n1392, new_n1393;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT64), .Z(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(KEYINPUT65), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n220), .A2(KEYINPUT65), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n209), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n212), .B(new_n217), .C1(new_n226), .C2(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  NOR2_X1   g0044(.A1(G20), .A2(G33), .ZN(new_n245));
  AOI22_X1  g0045(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT8), .B(G58), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n207), .A2(G33), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n215), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n202), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n254), .A2(new_n251), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n206), .A2(G20), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G50), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n252), .B(new_n255), .C1(new_n257), .C2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(KEYINPUT9), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n262), .A2(G222), .ZN(new_n263));
  XOR2_X1   g0063(.A(KEYINPUT68), .B(G223), .Z(new_n264));
  AOI21_X1  g0064(.A(new_n263), .B1(new_n264), .B2(G1698), .ZN(new_n265));
  INV_X1    g0065(.A(G77), .ZN(new_n266));
  AND2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  OAI21_X1  g0068(.A(KEYINPUT67), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT3), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT67), .ZN(new_n273));
  NAND2_X1  g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n269), .A2(new_n275), .ZN(new_n276));
  MUX2_X1   g0076(.A(new_n265), .B(new_n266), .S(new_n276), .Z(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(G1), .A3(G13), .ZN(new_n279));
  OR2_X1    g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n206), .B(G274), .C1(G41), .C2(G45), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G226), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n281), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(G200), .B1(new_n280), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n277), .A2(new_n279), .ZN(new_n288));
  NOR3_X1   g0088(.A1(new_n288), .A2(G190), .A3(new_n285), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n261), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT72), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT10), .ZN(new_n292));
  OR2_X1    g0092(.A1(new_n291), .A2(KEYINPUT10), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n290), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n280), .A2(new_n295), .A3(new_n286), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n288), .A2(new_n285), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n296), .B1(G200), .B2(new_n297), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n298), .A2(new_n291), .A3(KEYINPUT10), .A4(new_n261), .ZN(new_n299));
  INV_X1    g0099(.A(G169), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G179), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n288), .A2(new_n302), .A3(new_n285), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n260), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n294), .A2(new_n299), .A3(new_n304), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n269), .A2(new_n275), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n262), .A2(G232), .ZN(new_n307));
  NAND2_X1  g0107(.A1(G238), .A2(G1698), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(KEYINPUT69), .A2(G107), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(KEYINPUT69), .A2(G107), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n269), .B2(new_n275), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n279), .B1(new_n310), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G244), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n281), .B1(new_n283), .B2(new_n318), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n317), .A2(G179), .A3(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n300), .B1(new_n317), .B2(new_n319), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n320), .B1(KEYINPUT71), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n279), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n276), .B1(new_n308), .B2(new_n307), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(new_n315), .ZN(new_n325));
  INV_X1    g0125(.A(new_n319), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n325), .A2(KEYINPUT71), .A3(new_n302), .A4(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(G20), .A2(G77), .ZN(new_n328));
  INV_X1    g0128(.A(new_n245), .ZN(new_n329));
  XOR2_X1   g0129(.A(KEYINPUT15), .B(G87), .Z(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  OAI221_X1 g0131(.A(new_n328), .B1(new_n329), .B2(new_n247), .C1(new_n331), .C2(new_n248), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n251), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT70), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n258), .A2(G77), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n334), .B1(new_n257), .B2(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n256), .A2(KEYINPUT70), .A3(G77), .A4(new_n258), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n254), .A2(new_n266), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n333), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n327), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n322), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n325), .A2(new_n295), .A3(new_n326), .ZN(new_n343));
  INV_X1    g0143(.A(G200), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n344), .B1(new_n317), .B2(new_n319), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n340), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  OR3_X1    g0146(.A1(new_n305), .A2(new_n342), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n247), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n258), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n257), .A2(new_n349), .B1(new_n253), .B2(new_n348), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n267), .A2(new_n268), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n352), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n353));
  AOI21_X1  g0153(.A(G20), .B1(new_n269), .B2(new_n275), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n353), .B1(new_n354), .B2(KEYINPUT7), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G68), .ZN(new_n356));
  INV_X1    g0156(.A(G58), .ZN(new_n357));
  INV_X1    g0157(.A(G68), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(G20), .B1(new_n359), .B2(new_n201), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n245), .A2(G159), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT16), .B1(new_n356), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n272), .A2(new_n274), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT7), .ZN(new_n366));
  NOR3_X1   g0166(.A1(new_n365), .A2(new_n366), .A3(G20), .ZN(new_n367));
  AOI21_X1  g0167(.A(KEYINPUT7), .B1(new_n352), .B2(new_n207), .ZN(new_n368));
  OAI21_X1  g0168(.A(G68), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n363), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT16), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n251), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n351), .B1(new_n364), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n279), .A2(G232), .A3(new_n282), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n281), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT75), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n262), .A2(G223), .ZN(new_n377));
  NAND2_X1  g0177(.A1(G226), .A2(G1698), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n272), .A2(new_n274), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G87), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n271), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n323), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT75), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n374), .A2(new_n383), .A3(new_n281), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n376), .A2(new_n302), .A3(new_n382), .A4(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n377), .A2(new_n378), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n365), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n381), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n279), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n300), .B1(new_n389), .B2(new_n375), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n385), .A2(KEYINPUT76), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT76), .B1(new_n385), .B2(new_n390), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n373), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT18), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT18), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n373), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  OR2_X1    g0197(.A1(new_n364), .A2(new_n372), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n344), .B1(new_n389), .B2(new_n375), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n376), .A2(new_n384), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n382), .A2(new_n295), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n398), .A2(KEYINPUT17), .A3(new_n351), .A4(new_n402), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n351), .B(new_n402), .C1(new_n364), .C2(new_n372), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT17), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n395), .A2(new_n397), .A3(new_n403), .A4(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(KEYINPUT73), .B1(new_n254), .B2(new_n358), .ZN(new_n408));
  XNOR2_X1  g0208(.A(new_n408), .B(KEYINPUT12), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT11), .ZN(new_n410));
  OAI22_X1  g0210(.A1(new_n329), .A2(new_n202), .B1(new_n207), .B2(G68), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n248), .A2(new_n266), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n251), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n409), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n410), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n256), .A2(G68), .A3(new_n258), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT13), .ZN(new_n420));
  INV_X1    g0220(.A(G238), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n281), .B1(new_n283), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(G232), .A2(G1698), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(new_n284), .B2(G1698), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n269), .A2(new_n275), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G97), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n420), .B(new_n423), .C1(new_n428), .C2(new_n279), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n279), .B1(new_n426), .B2(new_n427), .ZN(new_n430));
  OAI21_X1  g0230(.A(KEYINPUT13), .B1(new_n430), .B2(new_n422), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n429), .A2(G179), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT14), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n429), .A2(new_n431), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n300), .A2(KEYINPUT74), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n432), .A2(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n434), .A2(new_n433), .A3(new_n435), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n419), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n434), .A2(G190), .ZN(new_n439));
  AOI21_X1  g0239(.A(G200), .B1(new_n429), .B2(new_n431), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n418), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n347), .A2(new_n407), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT84), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT24), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT23), .ZN(new_n446));
  INV_X1    g0246(.A(G107), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n446), .A2(new_n447), .A3(G20), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n448), .B1(G20), .B2(new_n449), .ZN(new_n450));
  OR2_X1    g0250(.A1(KEYINPUT69), .A2(G107), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n446), .B1(new_n451), .B2(new_n311), .ZN(new_n452));
  OAI21_X1  g0252(.A(KEYINPUT81), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT23), .B1(new_n312), .B2(new_n313), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G116), .ZN(new_n455));
  AOI21_X1  g0255(.A(G20), .B1(new_n455), .B2(new_n446), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT81), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n454), .A2(new_n457), .A3(new_n458), .A4(new_n448), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT80), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n380), .A2(KEYINPUT22), .A3(G20), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n269), .A2(new_n275), .A3(new_n462), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n207), .B(G87), .C1(new_n267), .C2(new_n268), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT22), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n460), .A2(new_n461), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n461), .B1(new_n460), .B2(new_n466), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n445), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n450), .A2(new_n452), .A3(KEYINPUT81), .ZN(new_n470));
  NOR3_X1   g0270(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n456), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n458), .B1(new_n472), .B2(new_n454), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n466), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT80), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n460), .A2(new_n461), .A3(new_n466), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n475), .A2(KEYINPUT24), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n469), .A2(new_n477), .A3(new_n251), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n254), .A2(new_n447), .ZN(new_n479));
  XNOR2_X1  g0279(.A(new_n479), .B(KEYINPUT25), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n206), .A2(G33), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n253), .A2(new_n481), .A3(new_n215), .A4(new_n250), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n480), .B1(new_n483), .B2(G107), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT82), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n262), .A2(G250), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n486), .B1(new_n352), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G294), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n271), .A2(new_n489), .ZN(new_n490));
  AND2_X1   g0290(.A1(G257), .A2(G1698), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n490), .B1(new_n365), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n365), .A2(KEYINPUT82), .A3(G250), .A4(new_n262), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n488), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n323), .ZN(new_n495));
  INV_X1    g0295(.A(G45), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(G1), .ZN(new_n497));
  AND2_X1   g0297(.A1(KEYINPUT5), .A2(G41), .ZN(new_n498));
  NOR2_X1   g0298(.A1(KEYINPUT5), .A2(G41), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AND3_X1   g0300(.A1(new_n500), .A2(G264), .A3(new_n279), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n497), .B(G274), .C1(new_n499), .C2(new_n498), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n495), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n504), .A2(new_n302), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n501), .B1(new_n494), .B2(new_n323), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n300), .B1(new_n506), .B2(new_n503), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n485), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n503), .ZN(new_n511));
  AOI211_X1 g0311(.A(new_n511), .B(new_n501), .C1(new_n494), .C2(new_n323), .ZN(new_n512));
  OAI21_X1  g0312(.A(KEYINPUT83), .B1(new_n512), .B2(G200), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT83), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n504), .A2(new_n514), .A3(new_n344), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n512), .A2(new_n295), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n513), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n517), .A2(new_n478), .A3(new_n484), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n444), .B1(new_n510), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n510), .A2(new_n444), .A3(new_n518), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n269), .A2(new_n275), .A3(G250), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n262), .B1(new_n523), .B2(KEYINPUT4), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT4), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n352), .B2(new_n318), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G283), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n262), .A2(KEYINPUT4), .A3(G244), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n526), .B(new_n527), .C1(new_n276), .C2(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n323), .B1(new_n524), .B2(new_n529), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n500), .A2(new_n279), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n511), .B1(new_n531), .B2(G257), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n302), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT77), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT77), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n530), .A2(new_n535), .A3(new_n302), .A4(new_n532), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n314), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n355), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n447), .A2(KEYINPUT6), .A3(G97), .ZN(new_n540));
  INV_X1    g0340(.A(G97), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n541), .A2(new_n447), .ZN(new_n542));
  NOR2_X1   g0342(.A1(G97), .A2(G107), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n540), .B1(new_n544), .B2(KEYINPUT6), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n545), .A2(G20), .B1(G77), .B2(new_n245), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n539), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n251), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n253), .A2(G97), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n483), .B2(G97), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n530), .A2(new_n532), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n548), .A2(new_n550), .B1(new_n551), .B2(new_n300), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n537), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(G244), .A2(G1698), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n421), .B2(G1698), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n365), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n279), .B1(new_n556), .B2(new_n455), .ZN(new_n557));
  OAI21_X1  g0357(.A(G250), .B1(new_n496), .B2(G1), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n497), .A2(G274), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n323), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n344), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n558), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n279), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n365), .A2(new_n555), .B1(G33), .B2(G116), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n563), .B(new_n295), .C1(new_n564), .C2(new_n279), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n330), .A2(new_n253), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n482), .A2(new_n380), .ZN(new_n568));
  NOR2_X1   g0368(.A1(G87), .A2(G97), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n451), .A2(new_n569), .A3(new_n311), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT19), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n207), .B1(new_n427), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n207), .B(G68), .C1(new_n267), .C2(new_n268), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n571), .B1(new_n427), .B2(G20), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  AOI211_X1 g0376(.A(new_n567), .B(new_n568), .C1(new_n576), .C2(new_n251), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n566), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n567), .B1(new_n576), .B2(new_n251), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n483), .A2(new_n330), .ZN(new_n580));
  OAI21_X1  g0380(.A(G169), .B1(new_n557), .B2(new_n560), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n563), .B(G179), .C1(new_n564), .C2(new_n279), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n579), .A2(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(KEYINPUT78), .B1(new_n578), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n579), .A2(new_n580), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n581), .A2(new_n582), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n566), .A2(new_n577), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT78), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n550), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(new_n547), .B2(new_n251), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n551), .A2(G190), .ZN(new_n594));
  AOI21_X1  g0394(.A(G200), .B1(new_n530), .B2(new_n532), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n553), .A2(new_n591), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n271), .A2(G97), .ZN(new_n598));
  AOI21_X1  g0398(.A(G20), .B1(new_n598), .B2(new_n527), .ZN(new_n599));
  INV_X1    g0399(.A(G116), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n207), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n251), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT20), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(KEYINPUT20), .B(new_n251), .C1(new_n599), .C2(new_n601), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n253), .A2(new_n600), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n483), .B2(new_n600), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n511), .B1(new_n531), .B2(G270), .ZN(new_n611));
  INV_X1    g0411(.A(G303), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n612), .B1(new_n269), .B2(new_n275), .ZN(new_n613));
  NAND2_X1  g0413(.A1(G264), .A2(G1698), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n262), .A2(G257), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n352), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n323), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT79), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n611), .A2(new_n617), .A3(KEYINPUT79), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n620), .A2(new_n344), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(G190), .B1(new_n620), .B2(new_n621), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n610), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n300), .B1(new_n606), .B2(new_n608), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n620), .A2(new_n621), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT21), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n618), .A2(new_n302), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n626), .A2(new_n627), .B1(new_n609), .B2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n620), .A2(new_n625), .A3(KEYINPUT21), .A4(new_n621), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n624), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n597), .A2(new_n631), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n443), .A2(new_n522), .A3(new_n632), .ZN(G372));
  AND3_X1   g0433(.A1(new_n373), .A2(new_n393), .A3(new_n396), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n396), .B1(new_n373), .B2(new_n393), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n342), .A2(new_n441), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n438), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n638), .A2(KEYINPUT85), .ZN(new_n639));
  XNOR2_X1  g0439(.A(new_n404), .B(KEYINPUT17), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n638), .B2(KEYINPUT85), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n636), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n642), .A2(new_n299), .A3(new_n294), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n643), .A2(new_n304), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n588), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n508), .B1(new_n478), .B2(new_n484), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n626), .A2(new_n627), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n628), .A2(new_n609), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(new_n649), .A3(new_n630), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n518), .B(new_n596), .C1(new_n647), .C2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n646), .B1(new_n651), .B2(new_n553), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n589), .B1(new_n587), .B2(new_n588), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n537), .B(new_n552), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n587), .B1(new_n656), .B2(new_n645), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n443), .B1(new_n652), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n644), .A2(new_n658), .ZN(G369));
  NAND3_X1  g0459(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(G213), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT86), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n664), .A2(G343), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(G343), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n668), .B1(new_n478), .B2(new_n484), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n669), .B1(new_n520), .B2(new_n521), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n647), .A2(new_n667), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n631), .B1(new_n610), .B2(new_n668), .ZN(new_n674));
  INV_X1    g0474(.A(new_n650), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n675), .A2(new_n609), .A3(new_n667), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(G330), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n673), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n510), .A2(new_n667), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n675), .A2(new_n667), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n681), .B1(new_n670), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n680), .A2(new_n683), .ZN(G399));
  INV_X1    g0484(.A(new_n210), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(G41), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n570), .A2(G116), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G1), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n214), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n689), .B1(new_n690), .B2(new_n687), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT28), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n655), .A2(new_n645), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n537), .A2(new_n552), .A3(KEYINPUT26), .A4(new_n588), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n583), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n517), .A2(new_n478), .A3(new_n484), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n696), .B1(new_n510), .B2(new_n675), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n587), .A2(new_n588), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n553), .A2(new_n596), .A3(new_n699), .ZN(new_n700));
  AOI22_X1  g0500(.A1(new_n695), .A2(KEYINPUT88), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n537), .A2(new_n552), .ZN(new_n702));
  AOI21_X1  g0502(.A(KEYINPUT26), .B1(new_n702), .B2(new_n591), .ZN(new_n703));
  INV_X1    g0503(.A(new_n694), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n587), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT88), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n667), .B1(new_n701), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT29), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n668), .B1(new_n652), .B2(new_n657), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT29), .ZN(new_n711));
  AOI21_X1  g0511(.A(KEYINPUT87), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n710), .A2(KEYINPUT87), .A3(new_n711), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n709), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n696), .A2(new_n647), .A3(KEYINPUT84), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n632), .B(new_n668), .C1(new_n715), .C2(new_n519), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT30), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n557), .A2(new_n560), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n506), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n628), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n717), .B1(new_n720), .B2(new_n551), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n512), .A2(G179), .A3(new_n718), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n722), .A2(new_n620), .A3(new_n621), .A4(new_n551), .ZN(new_n723));
  INV_X1    g0523(.A(new_n551), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n724), .A2(KEYINPUT30), .A3(new_n628), .A4(new_n719), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n721), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n726), .A2(KEYINPUT31), .A3(new_n667), .ZN(new_n727));
  AOI21_X1  g0527(.A(KEYINPUT31), .B1(new_n726), .B2(new_n667), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n716), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G330), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n714), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n692), .B1(new_n733), .B2(G1), .ZN(G364));
  INV_X1    g0534(.A(new_n679), .ZN(new_n735));
  INV_X1    g0535(.A(G13), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G20), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G45), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n687), .A2(G1), .A3(new_n738), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n739), .A2(KEYINPUT89), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(KEYINPUT89), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n677), .A2(new_n678), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n735), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n215), .B1(G20), .B2(new_n300), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n207), .A2(G190), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n747), .A2(new_n302), .A3(new_n344), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n748), .A2(KEYINPUT91), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(KEYINPUT91), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(G159), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT32), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n295), .A2(G179), .A3(G200), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n207), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G97), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n302), .A2(new_n344), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n747), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n302), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n747), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n760), .A2(new_n358), .B1(new_n762), .B2(new_n266), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n276), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n344), .A2(G179), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n747), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n447), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n207), .A2(new_n295), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n759), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n767), .B1(G50), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n768), .A2(new_n761), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n771), .B1(new_n357), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n768), .A2(new_n765), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n774), .A2(KEYINPUT92), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(KEYINPUT92), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n773), .B1(G87), .B2(new_n778), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n754), .A2(new_n758), .A3(new_n764), .A4(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n760), .ZN(new_n781));
  XNOR2_X1  g0581(.A(KEYINPUT33), .B(G317), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G326), .A2(new_n770), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G283), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n783), .B1(new_n784), .B2(new_n766), .ZN(new_n785));
  INV_X1    g0585(.A(new_n751), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n785), .B1(G329), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G322), .ZN(new_n788));
  INV_X1    g0588(.A(G311), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n772), .A2(new_n788), .B1(new_n762), .B2(new_n789), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n306), .B(new_n790), .C1(G294), .C2(new_n757), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n787), .B(new_n791), .C1(new_n612), .C2(new_n777), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n746), .B1(new_n780), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G13), .A2(G33), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(G20), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n745), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n685), .A2(new_n276), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n798), .A2(G355), .B1(new_n600), .B2(new_n685), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n685), .A2(new_n365), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(new_n214), .B2(new_n496), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(KEYINPUT90), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(new_n496), .B2(new_n243), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n802), .A2(KEYINPUT90), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n799), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n742), .B(new_n793), .C1(new_n797), .C2(new_n806), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT93), .Z(new_n808));
  INV_X1    g0608(.A(new_n677), .ZN(new_n809));
  INV_X1    g0609(.A(new_n796), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n744), .B1(new_n808), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n812), .A2(KEYINPUT94), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n812), .A2(KEYINPUT94), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(G396));
  NAND2_X1  g0616(.A1(new_n343), .A2(new_n345), .ZN(new_n817));
  INV_X1    g0617(.A(new_n340), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n340), .A2(new_n667), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n327), .A2(new_n340), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n325), .A2(new_n302), .A3(new_n326), .ZN(new_n822));
  AOI21_X1  g0622(.A(G169), .B1(new_n325), .B2(new_n326), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT71), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n819), .A2(new_n820), .B1(new_n821), .B2(new_n825), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n322), .A2(new_n341), .A3(new_n667), .ZN(new_n827));
  OAI21_X1  g0627(.A(KEYINPUT96), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n821), .A2(new_n825), .A3(new_n668), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT96), .ZN(new_n830));
  INV_X1    g0630(.A(new_n820), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n346), .A2(new_n831), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n829), .B(new_n830), .C1(new_n342), .C2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n828), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n668), .B(new_n834), .C1(new_n652), .C2(new_n657), .ZN(new_n835));
  INV_X1    g0635(.A(new_n710), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT97), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n834), .B(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n835), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n742), .B1(new_n839), .B2(new_n731), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n839), .A2(new_n731), .ZN(new_n842));
  INV_X1    g0642(.A(new_n834), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n794), .ZN(new_n844));
  INV_X1    g0644(.A(new_n742), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n745), .A2(new_n794), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n845), .B1(G77), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n762), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n770), .A2(G137), .B1(new_n849), .B2(G159), .ZN(new_n850));
  INV_X1    g0650(.A(G143), .ZN(new_n851));
  INV_X1    g0651(.A(G150), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n850), .B1(new_n851), .B2(new_n772), .C1(new_n852), .C2(new_n760), .ZN(new_n853));
  XNOR2_X1  g0653(.A(KEYINPUT95), .B(KEYINPUT34), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n853), .B(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n365), .B1(new_n766), .B2(new_n358), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(G58), .B2(new_n757), .ZN(new_n857));
  INV_X1    g0657(.A(G132), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n857), .B1(new_n777), .B2(new_n202), .C1(new_n858), .C2(new_n751), .ZN(new_n859));
  AOI22_X1  g0659(.A1(G303), .A2(new_n770), .B1(new_n781), .B2(G283), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n489), .B2(new_n772), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(G311), .B2(new_n786), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n447), .B2(new_n777), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n849), .A2(G116), .ZN(new_n864));
  INV_X1    g0664(.A(new_n766), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(G87), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n758), .A2(new_n276), .A3(new_n864), .A4(new_n866), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n855), .A2(new_n859), .B1(new_n863), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n848), .B1(new_n868), .B2(new_n745), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n841), .A2(new_n842), .B1(new_n844), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(G384));
  OR2_X1    g0671(.A1(new_n545), .A2(KEYINPUT35), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(G116), .A3(new_n216), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(KEYINPUT35), .B2(new_n545), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n874), .A2(KEYINPUT36), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(KEYINPUT36), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n690), .A2(new_n266), .A3(new_n359), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n358), .A2(G50), .ZN(new_n878));
  OAI211_X1 g0678(.A(G1), .B(new_n736), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n875), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT98), .Z(new_n881));
  NAND2_X1  g0681(.A1(new_n432), .A2(new_n433), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n434), .A2(new_n435), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n434), .A2(new_n433), .A3(new_n435), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n418), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n668), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n251), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n366), .B1(new_n365), .B2(G20), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n353), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n362), .B1(new_n891), .B2(G68), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n889), .B1(new_n892), .B2(KEYINPUT16), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n370), .A2(new_n371), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n350), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n895), .A2(new_n663), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n407), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n663), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT76), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n381), .B1(new_n365), .B2(new_n386), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n302), .B1(new_n900), .B2(new_n279), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n374), .A2(new_n383), .A3(new_n281), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n383), .B1(new_n374), .B2(new_n281), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n375), .ZN(new_n905));
  AOI21_X1  g0705(.A(G169), .B1(new_n905), .B2(new_n382), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n899), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n385), .A2(KEYINPUT76), .A3(new_n390), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n898), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n404), .B1(new_n909), .B2(new_n895), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(KEYINPUT37), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n373), .A2(new_n898), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT37), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n394), .A2(new_n912), .A3(new_n913), .A4(new_n404), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n897), .A2(KEYINPUT38), .A3(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT39), .ZN(new_n917));
  INV_X1    g0717(.A(new_n912), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n394), .A2(new_n912), .A3(new_n404), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(KEYINPUT37), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n407), .A2(new_n918), .B1(new_n920), .B2(new_n914), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n916), .B(new_n917), .C1(new_n921), .C2(KEYINPUT38), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT100), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT38), .ZN(new_n924));
  INV_X1    g0724(.A(new_n896), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n636), .B2(new_n640), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n911), .A2(new_n914), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n916), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n922), .A2(new_n923), .B1(new_n929), .B2(KEYINPUT39), .ZN(new_n930));
  AOI211_X1 g0730(.A(KEYINPUT100), .B(new_n917), .C1(new_n928), .C2(new_n916), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n888), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n438), .B(new_n441), .C1(new_n418), .C2(new_n668), .ZN(new_n933));
  OAI21_X1  g0733(.A(KEYINPUT99), .B1(new_n438), .B2(new_n668), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT99), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n886), .A2(new_n935), .A3(new_n667), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n933), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n835), .B2(new_n829), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n929), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n636), .A2(new_n898), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n932), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n709), .B(new_n443), .C1(new_n712), .C2(new_n713), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n644), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n943), .B(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n937), .A2(new_n834), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n929), .A2(new_n730), .A3(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT40), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n920), .A2(new_n914), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n912), .B1(new_n636), .B2(new_n640), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n924), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n950), .B1(new_n953), .B2(new_n916), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n947), .B1(new_n716), .B2(new_n729), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n949), .A2(new_n950), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n443), .A2(new_n730), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n956), .B(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(G330), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n946), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n206), .B2(new_n737), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n946), .A2(new_n959), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n881), .B1(new_n961), .B2(new_n962), .ZN(G367));
  OR2_X1    g0763(.A1(new_n577), .A2(new_n668), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n964), .A2(new_n587), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n965), .A2(KEYINPUT101), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n699), .A2(new_n964), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(KEYINPUT101), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n796), .ZN(new_n971));
  AOI21_X1  g0771(.A(KEYINPUT106), .B1(new_n778), .B2(G116), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT46), .Z(new_n973));
  OAI22_X1  g0773(.A1(new_n541), .A2(new_n766), .B1(new_n762), .B2(new_n784), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n365), .B(new_n974), .C1(G294), .C2(new_n781), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n786), .A2(G317), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n769), .A2(new_n789), .B1(new_n772), .B2(new_n612), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT105), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n757), .A2(new_n538), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n975), .A2(new_n976), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n772), .ZN(new_n981));
  AOI22_X1  g0781(.A1(G150), .A2(new_n981), .B1(new_n781), .B2(G159), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n757), .A2(G68), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n982), .A2(new_n306), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n865), .A2(G77), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n202), .B2(new_n762), .C1(new_n851), .C2(new_n769), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(G58), .B2(new_n778), .ZN(new_n987));
  INV_X1    g0787(.A(G137), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n987), .B1(new_n988), .B2(new_n751), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n973), .A2(new_n980), .B1(new_n984), .B2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT47), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n990), .A2(new_n991), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n992), .A2(new_n745), .A3(new_n993), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n801), .A2(new_n235), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n796), .B(new_n745), .C1(new_n685), .C2(new_n330), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n742), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n971), .A2(new_n994), .A3(new_n997), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n553), .A2(new_n596), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n593), .A2(new_n668), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n670), .A2(new_n682), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1003), .A2(KEYINPUT42), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1002), .B1(new_n1004), .B2(new_n681), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n670), .A2(new_n682), .A3(new_n1002), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n1006), .A2(KEYINPUT42), .B1(new_n702), .B2(new_n668), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT43), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n970), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1008), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1005), .A2(new_n1009), .A3(new_n970), .A4(new_n1007), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n680), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1002), .B1(new_n702), .B2(new_n667), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(KEYINPUT102), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT102), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1014), .A2(new_n1021), .A3(new_n1018), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1020), .B(new_n1022), .C1(new_n1018), .C2(new_n1014), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n738), .A2(G1), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT104), .Z(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n683), .A2(new_n1017), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT45), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n683), .A2(new_n1017), .A3(KEYINPUT45), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n683), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT44), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1032), .A2(new_n1033), .A3(new_n1016), .ZN(new_n1034));
  OAI21_X1  g0834(.A(KEYINPUT44), .B1(new_n683), .B2(new_n1017), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1015), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(new_n680), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1003), .A2(KEYINPUT103), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT103), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n670), .A2(new_n1042), .A3(new_n682), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n671), .B(new_n672), .C1(new_n675), .C2(new_n667), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n735), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1044), .A2(new_n735), .A3(new_n1045), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1037), .A2(new_n1040), .A3(new_n1049), .A4(new_n733), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n733), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n686), .B(KEYINPUT41), .Z(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1026), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n998), .B1(new_n1023), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT107), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1055), .B(new_n1056), .ZN(G387));
  INV_X1    g0857(.A(new_n688), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n798), .A2(new_n1058), .B1(new_n447), .B2(new_n685), .ZN(new_n1059));
  AOI211_X1 g0859(.A(G45), .B(new_n1058), .C1(G68), .C2(G77), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(KEYINPUT109), .ZN(new_n1061));
  OAI21_X1  g0861(.A(KEYINPUT50), .B1(new_n247), .B2(G50), .ZN(new_n1062));
  OR3_X1    g0862(.A1(new_n247), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1060), .A2(KEYINPUT109), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n800), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n232), .A2(new_n496), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1059), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n742), .B1(new_n1068), .B2(new_n797), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n778), .A2(G294), .B1(G283), .B2(new_n757), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT48), .ZN(new_n1071));
  INV_X1    g0871(.A(G317), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n789), .A2(new_n760), .B1(new_n772), .B2(new_n1072), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n769), .A2(new_n788), .B1(new_n762), .B2(new_n612), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1070), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT111), .Z(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(KEYINPUT48), .B2(new_n1075), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  OR2_X1    g0880(.A1(new_n1080), .A2(KEYINPUT49), .ZN(new_n1081));
  INV_X1    g0881(.A(G326), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n352), .B1(new_n600), .B2(new_n766), .C1(new_n751), .C2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n1080), .B2(KEYINPUT49), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n757), .A2(new_n330), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1085), .B(new_n365), .C1(new_n541), .C2(new_n766), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n760), .A2(new_n247), .B1(new_n762), .B2(new_n358), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n769), .A2(new_n752), .B1(new_n772), .B2(new_n202), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  XOR2_X1   g0889(.A(KEYINPUT110), .B(G150), .Z(new_n1090));
  AOI22_X1  g0890(.A1(new_n786), .A2(new_n1090), .B1(new_n778), .B2(G77), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1081), .A2(new_n1084), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1069), .B1(new_n673), .B2(new_n810), .C1(new_n746), .C2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1048), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1026), .B1(new_n1095), .B2(new_n1046), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(KEYINPUT108), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT108), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1049), .A2(new_n1098), .A3(new_n1026), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1094), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1095), .A2(new_n1046), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n732), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1049), .A2(new_n733), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1102), .A2(new_n1103), .A3(new_n686), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1100), .A2(new_n1104), .ZN(G393));
  NAND2_X1  g0905(.A1(new_n1037), .A2(new_n1040), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n1103), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1107), .A2(new_n686), .A3(new_n1050), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1016), .A2(new_n796), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n240), .A2(new_n801), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n797), .B1(new_n541), .B2(new_n210), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n845), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n781), .A2(G50), .B1(new_n849), .B2(new_n348), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n757), .A2(G77), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1113), .A2(new_n1114), .A3(new_n365), .A4(new_n866), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n769), .A2(new_n852), .B1(new_n772), .B2(new_n752), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT51), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n1117), .B1(new_n358), .B2(new_n777), .C1(new_n851), .C2(new_n751), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n769), .A2(new_n1072), .B1(new_n772), .B2(new_n789), .ZN(new_n1119));
  XOR2_X1   g0919(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n1120));
  XNOR2_X1  g0920(.A(new_n1119), .B(new_n1120), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1121), .B1(new_n784), .B2(new_n777), .C1(new_n788), .C2(new_n751), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n306), .B1(G116), .B2(new_n757), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n767), .B1(G294), .B2(new_n849), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1123), .B(new_n1124), .C1(new_n612), .C2(new_n760), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n1115), .A2(new_n1118), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1112), .B1(new_n1126), .B2(new_n745), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1109), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n1106), .B2(new_n1025), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1108), .A2(new_n1130), .ZN(G390));
  AOI21_X1  g0931(.A(new_n678), .B1(new_n716), .B2(new_n729), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n948), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n835), .A2(new_n829), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n888), .B1(new_n1135), .B2(new_n937), .ZN(new_n1136));
  NOR3_X1   g0936(.A1(new_n1136), .A2(new_n930), .A3(new_n931), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n888), .B1(new_n953), .B2(new_n916), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  OAI211_X1 g0939(.A(KEYINPUT88), .B(new_n587), .C1(new_n703), .C2(new_n704), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n697), .A2(new_n700), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n695), .A2(KEYINPUT88), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n668), .B(new_n834), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n829), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1139), .B1(new_n1145), .B2(new_n937), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1134), .B1(new_n1137), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n929), .A2(KEYINPUT39), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n922), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1148), .B1(new_n1149), .B2(KEYINPUT100), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n931), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(new_n939), .C2(new_n888), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n827), .B1(new_n708), .B2(new_n834), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1138), .B1(new_n1153), .B2(new_n938), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1152), .A2(new_n1154), .A3(new_n1133), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1147), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n938), .B1(new_n731), .B2(new_n843), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1158), .A2(new_n1133), .B1(new_n829), .B2(new_n835), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1133), .A2(new_n1144), .A3(new_n829), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n937), .B1(new_n838), .B2(new_n1132), .ZN(new_n1161));
  OAI21_X1  g0961(.A(KEYINPUT113), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n838), .A2(new_n1132), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n938), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT113), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1164), .A2(new_n1153), .A3(new_n1165), .A4(new_n1133), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1159), .B1(new_n1162), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n443), .A2(G330), .A3(new_n730), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n944), .A2(new_n644), .A3(new_n1168), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n686), .B1(new_n1157), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1162), .A2(new_n1166), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1159), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1169), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1176), .A2(new_n1156), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1171), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1150), .A2(new_n794), .A3(new_n1151), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n742), .B1(new_n247), .B2(new_n846), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1114), .B(new_n276), .C1(new_n600), .C2(new_n772), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n769), .A2(new_n784), .B1(new_n762), .B2(new_n541), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n538), .B2(new_n781), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT115), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1181), .B(new_n1184), .C1(G87), .C2(new_n778), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n751), .A2(new_n489), .B1(new_n358), .B2(new_n766), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT116), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n778), .A2(new_n1090), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT53), .Z(new_n1189));
  AOI22_X1  g0989(.A1(new_n770), .A2(G128), .B1(new_n865), .B2(G50), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1190), .B1(new_n858), .B2(new_n772), .C1(new_n988), .C2(new_n760), .ZN(new_n1191));
  INV_X1    g0991(.A(G125), .ZN(new_n1192));
  XOR2_X1   g0992(.A(KEYINPUT54), .B(G143), .Z(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT114), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n751), .A2(new_n1192), .B1(new_n1194), .B2(new_n762), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n306), .B1(new_n752), .B2(new_n756), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n1191), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1185), .A2(new_n1187), .B1(new_n1189), .B2(new_n1197), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1179), .B(new_n1180), .C1(new_n746), .C2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n1156), .B2(new_n1025), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1178), .A2(new_n1200), .ZN(G378));
  INV_X1    g1001(.A(KEYINPUT121), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n260), .A2(new_n898), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n305), .A2(new_n1204), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n294), .A2(new_n299), .A3(new_n304), .A4(new_n1203), .ZN(new_n1206));
  XOR2_X1   g1006(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1205), .A2(new_n1206), .A3(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1208), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT120), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n949), .A2(new_n950), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n954), .A2(new_n955), .ZN(new_n1215));
  AND4_X1   g1015(.A1(new_n1213), .A2(new_n1214), .A3(G330), .A4(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1213), .B1(new_n956), .B2(G330), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1212), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(KEYINPUT118), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n1207), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT118), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1221), .A2(new_n1222), .A3(new_n1209), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1219), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1214), .A2(G330), .A3(new_n1215), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1218), .A2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1202), .B1(new_n1229), .B2(new_n943), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1226), .A2(KEYINPUT120), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n956), .A2(new_n1213), .A3(G330), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1227), .B1(new_n1233), .B2(new_n1212), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n943), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT122), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1212), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT122), .ZN(new_n1239));
  NOR4_X1   g1039(.A1(new_n1238), .A2(new_n943), .A3(new_n1239), .A4(new_n1227), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1230), .B1(new_n1236), .B2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n943), .B1(new_n1238), .B2(new_n1227), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(KEYINPUT121), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1218), .A2(new_n1235), .A3(new_n1228), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1239), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1234), .A2(KEYINPUT122), .A3(new_n1235), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1243), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1241), .A2(new_n1247), .A3(new_n1026), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1225), .A2(new_n794), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n845), .B1(G50), .B2(new_n847), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n365), .A2(G41), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n766), .A2(new_n357), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(G97), .B2(new_n781), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n770), .A2(G116), .B1(new_n849), .B2(new_n330), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1255), .A2(new_n1256), .A3(new_n983), .A4(new_n1251), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n772), .A2(new_n447), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT117), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1259), .B1(new_n266), .B2(new_n777), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1257), .B(new_n1260), .C1(G283), .C2(new_n786), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1253), .B1(new_n1261), .B2(KEYINPUT58), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n769), .A2(new_n1192), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n760), .A2(new_n858), .B1(new_n762), .B2(new_n988), .ZN(new_n1264));
  AOI211_X1 g1064(.A(new_n1263), .B(new_n1264), .C1(G128), .C2(new_n981), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n1265), .B1(new_n852), .B2(new_n756), .C1(new_n777), .C2(new_n1194), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(KEYINPUT59), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n786), .A2(G124), .ZN(new_n1268));
  AOI211_X1 g1068(.A(G33), .B(G41), .C1(new_n865), .C2(G159), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1267), .A2(new_n1268), .A3(new_n1269), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1266), .A2(KEYINPUT59), .ZN(new_n1271));
  OAI221_X1 g1071(.A(new_n1262), .B1(KEYINPUT58), .B2(new_n1261), .C1(new_n1270), .C2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1250), .B1(new_n1272), .B2(new_n745), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1249), .A2(new_n1273), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1274), .B(KEYINPUT119), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1248), .A2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1175), .B1(new_n1156), .B2(new_n1167), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(KEYINPUT123), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT123), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1279), .B(new_n1175), .C1(new_n1156), .C2(new_n1167), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1281), .A2(new_n1241), .A3(new_n1247), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT57), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1283), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n687), .B1(new_n1281), .B2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1276), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(G375));
  NAND2_X1  g1088(.A1(new_n938), .A2(new_n794), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n845), .B1(G68), .B2(new_n847), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n786), .A2(G128), .ZN(new_n1291));
  OAI221_X1 g1091(.A(new_n1291), .B1(new_n752), .B2(new_n777), .C1(new_n760), .C2(new_n1194), .ZN(new_n1292));
  AOI211_X1 g1092(.A(new_n352), .B(new_n1254), .C1(G50), .C2(new_n757), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(G137), .A2(new_n981), .B1(new_n849), .B2(G150), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1293), .B(new_n1294), .C1(new_n858), .C2(new_n769), .ZN(new_n1295));
  OAI22_X1  g1095(.A1(new_n769), .A2(new_n489), .B1(new_n772), .B2(new_n784), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1296), .B1(G116), .B2(new_n781), .ZN(new_n1297));
  OAI221_X1 g1097(.A(new_n1297), .B1(new_n541), .B2(new_n777), .C1(new_n612), .C2(new_n751), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n849), .A2(new_n538), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1085), .A2(new_n276), .A3(new_n985), .A4(new_n1299), .ZN(new_n1300));
  OAI22_X1  g1100(.A1(new_n1292), .A2(new_n1295), .B1(new_n1298), .B2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1290), .B1(new_n1301), .B2(new_n745), .ZN(new_n1302));
  AOI22_X1  g1102(.A1(new_n1174), .A2(new_n1026), .B1(new_n1289), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1176), .A2(new_n1053), .A3(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT124), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1304), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1308), .B1(new_n1307), .B2(new_n1306), .ZN(G381));
  INV_X1    g1109(.A(G378), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1287), .A2(new_n1310), .ZN(new_n1311));
  NOR3_X1   g1111(.A1(new_n1031), .A2(new_n1015), .A3(new_n1036), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n680), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1101), .A2(new_n732), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n687), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1129), .B1(new_n1316), .B2(new_n1107), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1100), .A2(new_n815), .A3(new_n1104), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1317), .A2(new_n1318), .A3(new_n870), .ZN(new_n1319));
  OR4_X1    g1119(.A1(G387), .A2(new_n1311), .A3(G381), .A4(new_n1319), .ZN(G407));
  NAND3_X1  g1120(.A1(new_n665), .A2(new_n666), .A3(G213), .ZN(new_n1321));
  OAI211_X1 g1121(.A(G407), .B(G213), .C1(new_n1311), .C2(new_n1321), .ZN(G409));
  AOI21_X1  g1122(.A(new_n815), .B1(new_n1100), .B2(new_n1104), .ZN(new_n1323));
  OAI211_X1 g1123(.A(new_n1317), .B(new_n1056), .C1(new_n1318), .C2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(G393), .A2(G396), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1100), .A2(new_n815), .A3(new_n1104), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1325), .A2(G390), .A3(new_n1326), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1324), .A2(new_n1055), .A3(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1055), .B1(new_n1324), .B2(new_n1327), .ZN(new_n1329));
  OAI21_X1  g1129(.A(KEYINPUT127), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1324), .A2(new_n1327), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1055), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT127), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1324), .A2(new_n1055), .A3(new_n1327), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1333), .A2(new_n1334), .A3(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1330), .A2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1276), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1338), .A2(G378), .A3(new_n1339), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1281), .A2(new_n1241), .A3(new_n1247), .A4(new_n1053), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1025), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1342), .B1(new_n1249), .B2(new_n1273), .ZN(new_n1343));
  AOI21_X1  g1143(.A(G378), .B1(new_n1341), .B2(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1340), .A2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT62), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1305), .A2(KEYINPUT60), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT60), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1167), .A2(new_n1169), .A3(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1348), .A2(new_n1350), .ZN(new_n1351));
  NOR2_X1   g1151(.A1(new_n1170), .A2(new_n687), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1304), .B1(new_n1351), .B2(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT125), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1353), .A2(new_n1354), .A3(G384), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1176), .A2(new_n686), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1356), .B1(new_n1348), .B2(new_n1350), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n870), .B1(new_n1357), .B2(new_n1304), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1355), .A2(new_n1358), .ZN(new_n1359));
  AOI21_X1  g1159(.A(new_n1354), .B1(new_n1353), .B2(G384), .ZN(new_n1360));
  NOR2_X1   g1160(.A1(new_n1359), .A2(new_n1360), .ZN(new_n1361));
  NAND4_X1  g1161(.A1(new_n1346), .A2(new_n1347), .A3(new_n1321), .A4(new_n1361), .ZN(new_n1362));
  INV_X1    g1162(.A(new_n1321), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1363), .A2(G2897), .ZN(new_n1364));
  INV_X1    g1164(.A(new_n1364), .ZN(new_n1365));
  OAI21_X1  g1165(.A(new_n1365), .B1(new_n1359), .B2(new_n1360), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1353), .A2(G384), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1367), .A2(KEYINPUT125), .ZN(new_n1368));
  NAND4_X1  g1168(.A1(new_n1368), .A2(new_n1355), .A3(new_n1358), .A4(new_n1364), .ZN(new_n1369));
  AND2_X1   g1169(.A1(new_n1366), .A2(new_n1369), .ZN(new_n1370));
  AOI21_X1  g1170(.A(new_n1344), .B1(new_n1287), .B2(G378), .ZN(new_n1371));
  OAI21_X1  g1171(.A(new_n1370), .B1(new_n1371), .B2(new_n1363), .ZN(new_n1372));
  INV_X1    g1172(.A(KEYINPUT61), .ZN(new_n1373));
  NAND3_X1  g1173(.A1(new_n1362), .A2(new_n1372), .A3(new_n1373), .ZN(new_n1374));
  AOI21_X1  g1174(.A(new_n1363), .B1(new_n1340), .B2(new_n1345), .ZN(new_n1375));
  AOI21_X1  g1175(.A(new_n1347), .B1(new_n1375), .B2(new_n1361), .ZN(new_n1376));
  OAI21_X1  g1176(.A(new_n1337), .B1(new_n1374), .B2(new_n1376), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1346), .A2(new_n1321), .ZN(new_n1378));
  AOI21_X1  g1178(.A(KEYINPUT61), .B1(new_n1378), .B2(new_n1370), .ZN(new_n1379));
  NAND3_X1  g1179(.A1(new_n1346), .A2(new_n1321), .A3(new_n1361), .ZN(new_n1380));
  XOR2_X1   g1180(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1381));
  NAND2_X1  g1181(.A1(new_n1380), .A2(new_n1381), .ZN(new_n1382));
  NAND2_X1  g1182(.A1(new_n1333), .A2(new_n1335), .ZN(new_n1383));
  NAND3_X1  g1183(.A1(new_n1375), .A2(KEYINPUT63), .A3(new_n1361), .ZN(new_n1384));
  NAND4_X1  g1184(.A1(new_n1379), .A2(new_n1382), .A3(new_n1383), .A4(new_n1384), .ZN(new_n1385));
  NAND2_X1  g1185(.A1(new_n1377), .A2(new_n1385), .ZN(G405));
  NAND2_X1  g1186(.A1(G375), .A2(G378), .ZN(new_n1387));
  NAND2_X1  g1187(.A1(new_n1387), .A2(new_n1311), .ZN(new_n1388));
  AND2_X1   g1188(.A1(new_n1330), .A2(new_n1336), .ZN(new_n1389));
  NAND2_X1  g1189(.A1(new_n1388), .A2(new_n1389), .ZN(new_n1390));
  NAND3_X1  g1190(.A1(new_n1337), .A2(new_n1387), .A3(new_n1311), .ZN(new_n1391));
  AND3_X1   g1191(.A1(new_n1390), .A2(new_n1361), .A3(new_n1391), .ZN(new_n1392));
  AOI21_X1  g1192(.A(new_n1361), .B1(new_n1390), .B2(new_n1391), .ZN(new_n1393));
  NOR2_X1   g1193(.A1(new_n1392), .A2(new_n1393), .ZN(G402));
endmodule


