

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733;

  XNOR2_X1 U371 ( .A(G113), .B(KEYINPUT3), .ZN(n440) );
  XNOR2_X1 U372 ( .A(n440), .B(G119), .ZN(n370) );
  NOR2_X1 U373 ( .A1(n588), .A2(n585), .ZN(n591) );
  NOR2_X2 U374 ( .A1(n599), .A2(n403), .ZN(n406) );
  XOR2_X2 U375 ( .A(G125), .B(G146), .Z(n524) );
  NAND2_X1 U376 ( .A1(n557), .A2(n613), .ZN(n548) );
  NOR2_X1 U377 ( .A1(n640), .A2(n549), .ZN(n547) );
  NOR2_X1 U378 ( .A1(n549), .A2(n550), .ZN(n399) );
  INV_X1 U379 ( .A(n589), .ZN(n624) );
  XNOR2_X1 U380 ( .A(n463), .B(n411), .ZN(n690) );
  INV_X1 U381 ( .A(KEYINPUT78), .ZN(n398) );
  AND2_X2 U382 ( .A1(n382), .A2(n417), .ZN(n445) );
  NAND2_X1 U383 ( .A1(n418), .A2(n362), .ZN(n417) );
  NOR2_X1 U384 ( .A1(n649), .A2(KEYINPUT2), .ZN(n651) );
  AND2_X1 U385 ( .A1(n426), .A2(n424), .ZN(n428) );
  OR2_X1 U386 ( .A1(n368), .A2(n729), .ZN(n395) );
  XNOR2_X1 U387 ( .A(n419), .B(KEYINPUT73), .ZN(n427) );
  XNOR2_X1 U388 ( .A(n547), .B(KEYINPUT42), .ZN(n731) );
  XNOR2_X1 U389 ( .A(n367), .B(n580), .ZN(n729) );
  XNOR2_X1 U390 ( .A(n429), .B(n584), .ZN(n588) );
  XNOR2_X1 U391 ( .A(n399), .B(n398), .ZN(n674) );
  NAND2_X1 U392 ( .A1(n431), .A2(n430), .ZN(n429) );
  AND2_X1 U393 ( .A1(n573), .A2(n589), .ZN(n402) );
  NOR2_X1 U394 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X1 U395 ( .A1(n623), .A2(n544), .ZN(n595) );
  INV_X1 U396 ( .A(n540), .ZN(n350) );
  XNOR2_X1 U397 ( .A(n626), .B(n492), .ZN(n581) );
  NOR2_X1 U398 ( .A1(G902), .A2(n690), .ZN(n467) );
  XNOR2_X1 U399 ( .A(n691), .B(n364), .ZN(n692) );
  XNOR2_X1 U400 ( .A(n463), .B(n412), .ZN(n490) );
  XNOR2_X1 U401 ( .A(n414), .B(n413), .ZN(n412) );
  XNOR2_X1 U402 ( .A(n456), .B(n454), .ZN(n414) );
  XNOR2_X1 U403 ( .A(n407), .B(n355), .ZN(n462) );
  XNOR2_X1 U404 ( .A(n460), .B(n461), .ZN(n407) );
  XOR2_X1 U405 ( .A(G116), .B(G107), .Z(n519) );
  XNOR2_X2 U406 ( .A(n548), .B(KEYINPUT19), .ZN(n570) );
  XNOR2_X2 U407 ( .A(n572), .B(KEYINPUT0), .ZN(n600) );
  AND2_X1 U408 ( .A1(n629), .A2(n447), .ZN(n541) );
  INV_X1 U409 ( .A(n600), .ZN(n431) );
  INV_X1 U410 ( .A(KEYINPUT75), .ZN(n371) );
  NAND2_X1 U411 ( .A1(n375), .A2(n373), .ZN(n640) );
  AND2_X1 U412 ( .A1(n377), .A2(n376), .ZN(n375) );
  NAND2_X1 U413 ( .A1(n374), .A2(n354), .ZN(n373) );
  AND2_X1 U414 ( .A1(n731), .A2(KEYINPUT46), .ZN(n425) );
  XNOR2_X1 U415 ( .A(n395), .B(n394), .ZN(n605) );
  INV_X1 U416 ( .A(KEYINPUT44), .ZN(n394) );
  NOR2_X1 U417 ( .A1(G953), .A2(G237), .ZN(n502) );
  INV_X1 U418 ( .A(G134), .ZN(n459) );
  XOR2_X1 U419 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n506) );
  XNOR2_X1 U420 ( .A(G140), .B(KEYINPUT99), .ZN(n505) );
  XNOR2_X1 U421 ( .A(n450), .B(n449), .ZN(n448) );
  XNOR2_X1 U422 ( .A(KEYINPUT23), .B(KEYINPUT92), .ZN(n450) );
  XNOR2_X1 U423 ( .A(G110), .B(KEYINPUT91), .ZN(n449) );
  XNOR2_X1 U424 ( .A(n480), .B(KEYINPUT24), .ZN(n451) );
  XNOR2_X1 U425 ( .A(G119), .B(G128), .ZN(n480) );
  XNOR2_X1 U426 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n481) );
  NAND2_X1 U427 ( .A1(n546), .A2(n545), .ZN(n549) );
  XNOR2_X1 U428 ( .A(n583), .B(KEYINPUT65), .ZN(n584) );
  XNOR2_X1 U429 ( .A(n468), .B(KEYINPUT66), .ZN(n469) );
  INV_X1 U430 ( .A(KEYINPUT1), .ZN(n468) );
  XNOR2_X1 U431 ( .A(G478), .B(n500), .ZN(n554) );
  NAND2_X1 U432 ( .A1(n383), .A2(n382), .ZN(n381) );
  NOR2_X1 U433 ( .A1(n655), .A2(n654), .ZN(n656) );
  INV_X1 U434 ( .A(n733), .ZN(n423) );
  NOR2_X1 U435 ( .A1(n674), .A2(n617), .ZN(n552) );
  XOR2_X1 U436 ( .A(KEYINPUT20), .B(KEYINPUT93), .Z(n478) );
  INV_X1 U437 ( .A(KEYINPUT48), .ZN(n435) );
  NAND2_X1 U438 ( .A1(G234), .A2(G237), .ZN(n470) );
  INV_X1 U439 ( .A(KEYINPUT45), .ZN(n390) );
  OR2_X1 U440 ( .A1(G237), .A2(G902), .ZN(n530) );
  NOR2_X1 U441 ( .A1(n615), .A2(n628), .ZN(n430) );
  INV_X1 U442 ( .A(KEYINPUT94), .ZN(n452) );
  XNOR2_X1 U443 ( .A(n439), .B(n438), .ZN(n437) );
  XNOR2_X1 U444 ( .A(KEYINPUT5), .B(KEYINPUT95), .ZN(n439) );
  XNOR2_X1 U445 ( .A(G137), .B(KEYINPUT74), .ZN(n438) );
  XNOR2_X1 U446 ( .A(n370), .B(KEYINPUT16), .ZN(n520) );
  INV_X1 U447 ( .A(KEYINPUT9), .ZN(n401) );
  XOR2_X1 U448 ( .A(G122), .B(G104), .Z(n518) );
  XOR2_X1 U449 ( .A(KEYINPUT11), .B(KEYINPUT101), .Z(n504) );
  XNOR2_X1 U450 ( .A(G902), .B(KEYINPUT15), .ZN(n607) );
  XNOR2_X1 U451 ( .A(n432), .B(n465), .ZN(n372) );
  XNOR2_X1 U452 ( .A(n464), .B(G110), .ZN(n432) );
  INV_X1 U453 ( .A(KEYINPUT71), .ZN(n464) );
  XNOR2_X1 U454 ( .A(G104), .B(G107), .ZN(n461) );
  NOR2_X1 U455 ( .A1(n623), .A2(n581), .ZN(n573) );
  XNOR2_X1 U456 ( .A(n416), .B(n361), .ZN(n564) );
  INV_X1 U457 ( .A(KEYINPUT98), .ZN(n405) );
  BUF_X1 U458 ( .A(n626), .Z(n403) );
  XNOR2_X1 U459 ( .A(n451), .B(n448), .ZN(n483) );
  NOR2_X1 U460 ( .A1(n558), .A2(n548), .ZN(n531) );
  NOR2_X1 U461 ( .A1(n576), .A2(n577), .ZN(n367) );
  XNOR2_X1 U462 ( .A(KEYINPUT32), .B(KEYINPUT64), .ZN(n433) );
  XNOR2_X1 U463 ( .A(n695), .B(n387), .ZN(n697) );
  XNOR2_X1 U464 ( .A(n696), .B(KEYINPUT122), .ZN(n387) );
  XNOR2_X1 U465 ( .A(n384), .B(n365), .ZN(G51) );
  XNOR2_X1 U466 ( .A(n379), .B(n659), .ZN(G75) );
  NAND2_X1 U467 ( .A1(n381), .A2(n380), .ZN(n379) );
  AND2_X1 U468 ( .A1(n658), .A2(n723), .ZN(n380) );
  AND2_X1 U469 ( .A1(n554), .A2(KEYINPUT41), .ZN(n351) );
  XOR2_X1 U470 ( .A(n687), .B(n366), .Z(n352) );
  XOR2_X1 U471 ( .A(KEYINPUT96), .B(G472), .Z(n353) );
  AND2_X1 U472 ( .A1(n553), .A2(n351), .ZN(n354) );
  XNOR2_X1 U473 ( .A(G137), .B(G140), .ZN(n355) );
  AND2_X1 U474 ( .A1(G221), .A2(n493), .ZN(n356) );
  XOR2_X1 U475 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n357) );
  AND2_X1 U476 ( .A1(G224), .A2(n723), .ZN(n358) );
  AND2_X1 U477 ( .A1(n403), .A2(n629), .ZN(n359) );
  XOR2_X1 U478 ( .A(n539), .B(KEYINPUT40), .Z(n360) );
  XOR2_X1 U479 ( .A(n538), .B(KEYINPUT39), .Z(n361) );
  INV_X1 U480 ( .A(KEYINPUT46), .ZN(n441) );
  INV_X1 U481 ( .A(KEYINPUT41), .ZN(n378) );
  OR2_X1 U482 ( .A1(n608), .A2(n607), .ZN(n362) );
  XOR2_X1 U483 ( .A(n490), .B(KEYINPUT62), .Z(n363) );
  XNOR2_X1 U484 ( .A(KEYINPUT121), .B(KEYINPUT59), .ZN(n364) );
  XOR2_X1 U485 ( .A(KEYINPUT56), .B(KEYINPUT120), .Z(n365) );
  XNOR2_X1 U486 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n366) );
  NOR2_X1 U487 ( .A1(G952), .A2(n723), .ZN(n701) );
  INV_X1 U488 ( .A(n701), .ZN(n385) );
  NAND2_X1 U489 ( .A1(n728), .A2(n668), .ZN(n368) );
  NAND2_X1 U490 ( .A1(n369), .A2(n359), .ZN(n668) );
  XNOR2_X1 U491 ( .A(n590), .B(KEYINPUT104), .ZN(n369) );
  XNOR2_X2 U492 ( .A(n587), .B(n433), .ZN(n728) );
  XNOR2_X1 U493 ( .A(n437), .B(n370), .ZN(n413) );
  XNOR2_X2 U494 ( .A(n611), .B(n371), .ZN(n382) );
  XNOR2_X1 U495 ( .A(n523), .B(n372), .ZN(n526) );
  XNOR2_X1 U496 ( .A(n462), .B(n372), .ZN(n411) );
  NAND2_X1 U497 ( .A1(n616), .A2(n378), .ZN(n377) );
  NAND2_X1 U498 ( .A1(n350), .A2(n613), .ZN(n616) );
  INV_X1 U499 ( .A(n616), .ZN(n374) );
  NAND2_X1 U500 ( .A1(n615), .A2(n378), .ZN(n376) );
  NAND2_X1 U501 ( .A1(n553), .A2(n554), .ZN(n615) );
  INV_X1 U502 ( .A(n657), .ZN(n383) );
  NAND2_X1 U503 ( .A1(n386), .A2(n385), .ZN(n384) );
  XNOR2_X1 U504 ( .A(n688), .B(n352), .ZN(n386) );
  INV_X1 U505 ( .A(n542), .ZN(n626) );
  XNOR2_X1 U506 ( .A(n388), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U507 ( .A1(n396), .A2(n385), .ZN(n388) );
  NAND2_X1 U508 ( .A1(n428), .A2(n427), .ZN(n436) );
  XNOR2_X1 U509 ( .A(n389), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U510 ( .A1(n694), .A2(n701), .ZN(n389) );
  XNOR2_X2 U511 ( .A(n391), .B(n390), .ZN(n652) );
  NAND2_X1 U512 ( .A1(n605), .A2(n604), .ZN(n391) );
  XNOR2_X2 U513 ( .A(n392), .B(n360), .ZN(n733) );
  NAND2_X1 U514 ( .A1(n564), .A2(n676), .ZN(n392) );
  XNOR2_X1 U515 ( .A(n561), .B(n537), .ZN(n540) );
  XNOR2_X1 U516 ( .A(n436), .B(n435), .ZN(n408) );
  NOR2_X1 U517 ( .A1(n609), .A2(n652), .ZN(n610) );
  NAND2_X1 U518 ( .A1(n565), .A2(n686), .ZN(n609) );
  NAND2_X1 U519 ( .A1(n393), .A2(n423), .ZN(n422) );
  NAND2_X1 U520 ( .A1(n397), .A2(n441), .ZN(n393) );
  XNOR2_X1 U521 ( .A(n612), .B(n363), .ZN(n396) );
  INV_X1 U522 ( .A(n731), .ZN(n397) );
  XOR2_X1 U523 ( .A(n446), .B(n543), .Z(n546) );
  XNOR2_X1 U524 ( .A(n400), .B(n497), .ZN(n498) );
  XNOR2_X1 U525 ( .A(n496), .B(n401), .ZN(n400) );
  XNOR2_X2 U526 ( .A(n402), .B(KEYINPUT33), .ZN(n622) );
  NAND2_X1 U527 ( .A1(n404), .A2(n649), .ZN(n418) );
  XNOR2_X1 U528 ( .A(n606), .B(KEYINPUT82), .ZN(n404) );
  XNOR2_X1 U529 ( .A(n406), .B(n405), .ZN(n634) );
  XNOR2_X1 U530 ( .A(n509), .B(n355), .ZN(n716) );
  XNOR2_X1 U531 ( .A(n716), .B(n484), .ZN(n699) );
  XNOR2_X1 U532 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U533 ( .A(n527), .B(n710), .ZN(n687) );
  NOR2_X1 U534 ( .A1(n425), .A2(n683), .ZN(n424) );
  NOR2_X2 U535 ( .A1(G902), .A2(n490), .ZN(n491) );
  NOR2_X1 U536 ( .A1(n535), .A2(n628), .ZN(n447) );
  XNOR2_X2 U537 ( .A(n491), .B(n353), .ZN(n542) );
  XNOR2_X1 U538 ( .A(n574), .B(n575), .ZN(n576) );
  NOR2_X2 U539 ( .A1(n652), .A2(n607), .ZN(n606) );
  XNOR2_X2 U540 ( .A(n609), .B(KEYINPUT83), .ZN(n649) );
  INV_X4 U541 ( .A(G953), .ZN(n723) );
  XNOR2_X1 U542 ( .A(n522), .B(n358), .ZN(n523) );
  XNOR2_X1 U543 ( .A(n434), .B(KEYINPUT85), .ZN(n565) );
  NAND2_X1 U544 ( .A1(n408), .A2(n730), .ZN(n434) );
  NAND2_X1 U545 ( .A1(n420), .A2(n672), .ZN(n419) );
  XNOR2_X2 U546 ( .A(n522), .B(n459), .ZN(n496) );
  XNOR2_X2 U547 ( .A(n458), .B(G128), .ZN(n522) );
  NAND2_X1 U548 ( .A1(n409), .A2(n602), .ZN(n603) );
  INV_X1 U549 ( .A(n410), .ZN(n409) );
  NOR2_X1 U550 ( .A1(n680), .A2(n664), .ZN(n410) );
  XNOR2_X2 U551 ( .A(n717), .B(G146), .ZN(n463) );
  XNOR2_X2 U552 ( .A(n496), .B(n510), .ZN(n717) );
  NAND2_X1 U553 ( .A1(n536), .A2(n595), .ZN(n555) );
  NAND2_X1 U554 ( .A1(n415), .A2(n536), .ZN(n416) );
  AND2_X1 U555 ( .A1(n595), .A2(n350), .ZN(n415) );
  XNOR2_X1 U556 ( .A(n552), .B(KEYINPUT47), .ZN(n420) );
  NAND2_X1 U557 ( .A1(n422), .A2(n421), .ZN(n426) );
  NAND2_X1 U558 ( .A1(n733), .A2(n441), .ZN(n421) );
  NAND2_X1 U559 ( .A1(n570), .A2(n571), .ZN(n572) );
  XNOR2_X2 U560 ( .A(n529), .B(n528), .ZN(n557) );
  XNOR2_X2 U561 ( .A(KEYINPUT4), .B(G101), .ZN(n465) );
  INV_X2 U562 ( .A(G143), .ZN(n458) );
  NOR2_X1 U563 ( .A1(n442), .A2(n701), .ZN(G54) );
  XNOR2_X1 U564 ( .A(n444), .B(n443), .ZN(n442) );
  XNOR2_X1 U565 ( .A(n690), .B(n689), .ZN(n443) );
  NAND2_X1 U566 ( .A1(n445), .A2(G469), .ZN(n444) );
  NAND2_X1 U567 ( .A1(n445), .A2(G475), .ZN(n693) );
  NAND2_X1 U568 ( .A1(n445), .A2(G472), .ZN(n612) );
  NAND2_X1 U569 ( .A1(n445), .A2(G210), .ZN(n688) );
  NAND2_X1 U570 ( .A1(n445), .A2(G478), .ZN(n695) );
  NAND2_X1 U571 ( .A1(n445), .A2(G217), .ZN(n698) );
  NAND2_X1 U572 ( .A1(n541), .A2(n542), .ZN(n446) );
  XNOR2_X1 U573 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U574 ( .A(n483), .B(n356), .ZN(n484) );
  XNOR2_X1 U575 ( .A(n453), .B(n452), .ZN(n454) );
  INV_X1 U576 ( .A(KEYINPUT81), .ZN(n650) );
  XNOR2_X1 U577 ( .A(n524), .B(n357), .ZN(n525) );
  XNOR2_X1 U578 ( .A(KEYINPUT103), .B(KEYINPUT6), .ZN(n492) );
  INV_X1 U579 ( .A(KEYINPUT77), .ZN(n578) );
  XNOR2_X1 U580 ( .A(n579), .B(n578), .ZN(n580) );
  NAND2_X1 U581 ( .A1(n502), .A2(G210), .ZN(n453) );
  INV_X1 U582 ( .A(n465), .ZN(n455) );
  XNOR2_X1 U583 ( .A(G116), .B(n455), .ZN(n456) );
  XNOR2_X1 U584 ( .A(G131), .B(KEYINPUT69), .ZN(n457) );
  XNOR2_X1 U585 ( .A(n457), .B(KEYINPUT68), .ZN(n510) );
  NAND2_X1 U586 ( .A1(n723), .A2(G227), .ZN(n460) );
  XNOR2_X1 U587 ( .A(KEYINPUT70), .B(G469), .ZN(n466) );
  XNOR2_X2 U588 ( .A(n467), .B(n466), .ZN(n544) );
  XNOR2_X2 U589 ( .A(n544), .B(n469), .ZN(n589) );
  XNOR2_X1 U590 ( .A(n470), .B(KEYINPUT87), .ZN(n471) );
  XOR2_X1 U591 ( .A(KEYINPUT14), .B(n471), .Z(n474) );
  AND2_X1 U592 ( .A1(n474), .A2(G953), .ZN(n472) );
  NAND2_X1 U593 ( .A1(G902), .A2(n472), .ZN(n566) );
  XOR2_X1 U594 ( .A(n566), .B(KEYINPUT105), .Z(n473) );
  NOR2_X1 U595 ( .A1(G900), .A2(n473), .ZN(n476) );
  NAND2_X1 U596 ( .A1(n474), .A2(G952), .ZN(n646) );
  NOR2_X1 U597 ( .A1(G953), .A2(n646), .ZN(n475) );
  XNOR2_X1 U598 ( .A(KEYINPUT88), .B(n475), .ZN(n567) );
  NOR2_X1 U599 ( .A1(n476), .A2(n567), .ZN(n535) );
  NAND2_X1 U600 ( .A1(G234), .A2(n607), .ZN(n477) );
  XNOR2_X1 U601 ( .A(n478), .B(n477), .ZN(n485) );
  NAND2_X1 U602 ( .A1(G221), .A2(n485), .ZN(n479) );
  XNOR2_X1 U603 ( .A(n479), .B(KEYINPUT21), .ZN(n628) );
  INV_X1 U604 ( .A(n628), .ZN(n582) );
  XOR2_X1 U605 ( .A(KEYINPUT10), .B(n524), .Z(n509) );
  NAND2_X1 U606 ( .A1(n723), .A2(G234), .ZN(n482) );
  XNOR2_X1 U607 ( .A(n482), .B(n481), .ZN(n493) );
  NOR2_X1 U608 ( .A1(n699), .A2(G902), .ZN(n489) );
  XOR2_X1 U609 ( .A(KEYINPUT25), .B(KEYINPUT76), .Z(n487) );
  NAND2_X1 U610 ( .A1(G217), .A2(n485), .ZN(n486) );
  XNOR2_X1 U611 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U612 ( .A(n489), .B(n488), .ZN(n629) );
  XOR2_X1 U613 ( .A(KEYINPUT7), .B(KEYINPUT102), .Z(n495) );
  NAND2_X1 U614 ( .A1(G217), .A2(n493), .ZN(n494) );
  XNOR2_X1 U615 ( .A(n495), .B(n494), .ZN(n499) );
  XNOR2_X1 U616 ( .A(G122), .B(n519), .ZN(n497) );
  XOR2_X1 U617 ( .A(n499), .B(n498), .Z(n696) );
  NOR2_X1 U618 ( .A1(G902), .A2(n696), .ZN(n500) );
  XNOR2_X1 U619 ( .A(G113), .B(n518), .ZN(n501) );
  XNOR2_X1 U620 ( .A(n501), .B(G143), .ZN(n514) );
  NAND2_X1 U621 ( .A1(G214), .A2(n502), .ZN(n503) );
  XNOR2_X1 U622 ( .A(n504), .B(n503), .ZN(n508) );
  XNOR2_X1 U623 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U624 ( .A(n508), .B(n507), .Z(n512) );
  XNOR2_X1 U625 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U626 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U627 ( .A(n514), .B(n513), .ZN(n691) );
  NOR2_X1 U628 ( .A1(G902), .A2(n691), .ZN(n516) );
  XNOR2_X1 U629 ( .A(KEYINPUT13), .B(G475), .ZN(n515) );
  XNOR2_X1 U630 ( .A(n516), .B(n515), .ZN(n551) );
  NAND2_X1 U631 ( .A1(n554), .A2(n551), .ZN(n673) );
  NOR2_X1 U632 ( .A1(n581), .A2(n673), .ZN(n517) );
  NAND2_X1 U633 ( .A1(n541), .A2(n517), .ZN(n558) );
  XOR2_X1 U634 ( .A(n519), .B(n518), .Z(n521) );
  XNOR2_X1 U635 ( .A(n521), .B(n520), .ZN(n710) );
  NAND2_X1 U636 ( .A1(n687), .A2(n607), .ZN(n529) );
  AND2_X1 U637 ( .A1(G210), .A2(n530), .ZN(n528) );
  NAND2_X1 U638 ( .A1(G214), .A2(n530), .ZN(n613) );
  XOR2_X1 U639 ( .A(KEYINPUT36), .B(n531), .Z(n532) );
  NOR2_X1 U640 ( .A1(n624), .A2(n532), .ZN(n683) );
  INV_X1 U641 ( .A(KEYINPUT109), .ZN(n539) );
  INV_X1 U642 ( .A(n629), .ZN(n593) );
  NAND2_X1 U643 ( .A1(n582), .A2(n593), .ZN(n623) );
  NAND2_X1 U644 ( .A1(n542), .A2(n613), .ZN(n533) );
  XNOR2_X1 U645 ( .A(KEYINPUT30), .B(n533), .ZN(n534) );
  INV_X1 U646 ( .A(KEYINPUT38), .ZN(n537) );
  INV_X1 U647 ( .A(n557), .ZN(n561) );
  INV_X1 U648 ( .A(KEYINPUT86), .ZN(n538) );
  INV_X1 U649 ( .A(n673), .ZN(n676) );
  INV_X1 U650 ( .A(n551), .ZN(n553) );
  XNOR2_X1 U651 ( .A(KEYINPUT28), .B(KEYINPUT108), .ZN(n543) );
  XNOR2_X1 U652 ( .A(n544), .B(KEYINPUT107), .ZN(n545) );
  INV_X1 U653 ( .A(n570), .ZN(n550) );
  NOR2_X1 U654 ( .A1(n551), .A2(n554), .ZN(n679) );
  NOR2_X1 U655 ( .A1(n679), .A2(n676), .ZN(n617) );
  OR2_X1 U656 ( .A1(n554), .A2(n553), .ZN(n577) );
  NOR2_X1 U657 ( .A1(n555), .A2(n577), .ZN(n556) );
  NAND2_X1 U658 ( .A1(n557), .A2(n556), .ZN(n672) );
  NOR2_X1 U659 ( .A1(n558), .A2(n589), .ZN(n559) );
  NAND2_X1 U660 ( .A1(n559), .A2(n613), .ZN(n560) );
  XNOR2_X1 U661 ( .A(n560), .B(KEYINPUT43), .ZN(n562) );
  NAND2_X1 U662 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U663 ( .A(KEYINPUT106), .B(n563), .ZN(n730) );
  NAND2_X1 U664 ( .A1(n679), .A2(n564), .ZN(n686) );
  INV_X1 U665 ( .A(n649), .ZN(n719) );
  INV_X1 U666 ( .A(KEYINPUT34), .ZN(n575) );
  NOR2_X1 U667 ( .A1(G898), .A2(n566), .ZN(n568) );
  NOR2_X1 U668 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U669 ( .A(KEYINPUT89), .B(n569), .ZN(n571) );
  XNOR2_X1 U670 ( .A(n600), .B(KEYINPUT90), .ZN(n594) );
  NOR2_X1 U671 ( .A1(n594), .A2(n622), .ZN(n574) );
  XOR2_X1 U672 ( .A(KEYINPUT84), .B(KEYINPUT35), .Z(n579) );
  INV_X1 U673 ( .A(n581), .ZN(n585) );
  XOR2_X1 U674 ( .A(KEYINPUT22), .B(KEYINPUT72), .Z(n583) );
  NOR2_X1 U675 ( .A1(n593), .A2(n624), .ZN(n586) );
  NAND2_X1 U676 ( .A1(n591), .A2(n586), .ZN(n587) );
  NOR2_X1 U677 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U678 ( .A1(n591), .A2(n624), .ZN(n592) );
  NAND2_X1 U679 ( .A1(n593), .A2(n592), .ZN(n660) );
  INV_X1 U680 ( .A(n617), .ZN(n602) );
  INV_X1 U681 ( .A(n594), .ZN(n597) );
  AND2_X1 U682 ( .A1(n403), .A2(n595), .ZN(n596) );
  NAND2_X1 U683 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U684 ( .A(KEYINPUT97), .B(n598), .ZN(n664) );
  OR2_X1 U685 ( .A1(n623), .A2(n624), .ZN(n599) );
  NOR2_X1 U686 ( .A1(n600), .A2(n634), .ZN(n601) );
  XOR2_X1 U687 ( .A(KEYINPUT31), .B(n601), .Z(n680) );
  AND2_X1 U688 ( .A1(n660), .A2(n603), .ZN(n604) );
  INV_X1 U689 ( .A(KEYINPUT2), .ZN(n608) );
  NAND2_X1 U690 ( .A1(KEYINPUT2), .A2(n610), .ZN(n611) );
  NOR2_X1 U691 ( .A1(n640), .A2(n622), .ZN(n648) );
  NOR2_X1 U692 ( .A1(n350), .A2(n613), .ZN(n614) );
  NOR2_X1 U693 ( .A1(n615), .A2(n614), .ZN(n619) );
  NOR2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U696 ( .A(n620), .B(KEYINPUT118), .ZN(n621) );
  NOR2_X1 U697 ( .A1(n622), .A2(n621), .ZN(n643) );
  NAND2_X1 U698 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U699 ( .A(KEYINPUT50), .B(n625), .ZN(n627) );
  NAND2_X1 U700 ( .A1(n627), .A2(n403), .ZN(n633) );
  XNOR2_X1 U701 ( .A(KEYINPUT49), .B(KEYINPUT115), .ZN(n631) );
  NAND2_X1 U702 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U703 ( .A(n631), .B(n630), .Z(n632) );
  NOR2_X1 U704 ( .A1(n633), .A2(n632), .ZN(n636) );
  INV_X1 U705 ( .A(n634), .ZN(n635) );
  NOR2_X1 U706 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U707 ( .A(KEYINPUT116), .B(n637), .Z(n638) );
  XNOR2_X1 U708 ( .A(n638), .B(KEYINPUT51), .ZN(n639) );
  NOR2_X1 U709 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U710 ( .A(KEYINPUT117), .B(n641), .Z(n642) );
  NOR2_X1 U711 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U712 ( .A(n644), .B(KEYINPUT52), .ZN(n645) );
  NOR2_X1 U713 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U714 ( .A1(n648), .A2(n647), .ZN(n658) );
  XNOR2_X1 U715 ( .A(n651), .B(n650), .ZN(n655) );
  INV_X1 U716 ( .A(n652), .ZN(n702) );
  NOR2_X1 U717 ( .A1(n702), .A2(KEYINPUT2), .ZN(n653) );
  XNOR2_X1 U718 ( .A(KEYINPUT80), .B(n653), .ZN(n654) );
  XNOR2_X1 U719 ( .A(n656), .B(KEYINPUT79), .ZN(n657) );
  XNOR2_X1 U720 ( .A(KEYINPUT53), .B(KEYINPUT119), .ZN(n659) );
  XNOR2_X1 U721 ( .A(G101), .B(KEYINPUT110), .ZN(n661) );
  XNOR2_X1 U722 ( .A(n661), .B(n660), .ZN(G3) );
  XOR2_X1 U723 ( .A(G104), .B(KEYINPUT111), .Z(n663) );
  NAND2_X1 U724 ( .A1(n664), .A2(n676), .ZN(n662) );
  XNOR2_X1 U725 ( .A(n663), .B(n662), .ZN(G6) );
  XOR2_X1 U726 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n666) );
  NAND2_X1 U727 ( .A1(n664), .A2(n679), .ZN(n665) );
  XNOR2_X1 U728 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U729 ( .A(G107), .B(n667), .ZN(G9) );
  XNOR2_X1 U730 ( .A(G110), .B(n668), .ZN(G12) );
  INV_X1 U731 ( .A(n679), .ZN(n669) );
  NOR2_X1 U732 ( .A1(n674), .A2(n669), .ZN(n671) );
  XNOR2_X1 U733 ( .A(G128), .B(KEYINPUT29), .ZN(n670) );
  XNOR2_X1 U734 ( .A(n671), .B(n670), .ZN(G30) );
  XNOR2_X1 U735 ( .A(G143), .B(n672), .ZN(G45) );
  NOR2_X1 U736 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U737 ( .A(G146), .B(n675), .Z(G48) );
  NAND2_X1 U738 ( .A1(n680), .A2(n676), .ZN(n677) );
  XNOR2_X1 U739 ( .A(n677), .B(KEYINPUT112), .ZN(n678) );
  XNOR2_X1 U740 ( .A(G113), .B(n678), .ZN(G15) );
  XOR2_X1 U741 ( .A(G116), .B(KEYINPUT113), .Z(n682) );
  NAND2_X1 U742 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U743 ( .A(n682), .B(n681), .ZN(G18) );
  XNOR2_X1 U744 ( .A(n683), .B(KEYINPUT37), .ZN(n684) );
  XNOR2_X1 U745 ( .A(n684), .B(KEYINPUT114), .ZN(n685) );
  XNOR2_X1 U746 ( .A(G125), .B(n685), .ZN(G27) );
  XNOR2_X1 U747 ( .A(G134), .B(n686), .ZN(G36) );
  XOR2_X1 U748 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n689) );
  NOR2_X1 U749 ( .A1(n701), .A2(n697), .ZN(G63) );
  XNOR2_X1 U750 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U751 ( .A1(n701), .A2(n700), .ZN(G66) );
  NAND2_X1 U752 ( .A1(n723), .A2(n702), .ZN(n706) );
  NAND2_X1 U753 ( .A1(G953), .A2(G224), .ZN(n703) );
  XNOR2_X1 U754 ( .A(KEYINPUT61), .B(n703), .ZN(n704) );
  NAND2_X1 U755 ( .A1(n704), .A2(G898), .ZN(n705) );
  NAND2_X1 U756 ( .A1(n706), .A2(n705), .ZN(n714) );
  XOR2_X1 U757 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n708) );
  XNOR2_X1 U758 ( .A(G101), .B(G110), .ZN(n707) );
  XNOR2_X1 U759 ( .A(n708), .B(n707), .ZN(n709) );
  XOR2_X1 U760 ( .A(n710), .B(n709), .Z(n712) );
  NOR2_X1 U761 ( .A1(G898), .A2(n723), .ZN(n711) );
  NOR2_X1 U762 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U763 ( .A(n714), .B(n713), .ZN(n715) );
  XOR2_X1 U764 ( .A(KEYINPUT125), .B(n715), .Z(G69) );
  XNOR2_X1 U765 ( .A(KEYINPUT4), .B(n716), .ZN(n718) );
  XOR2_X1 U766 ( .A(n717), .B(n718), .Z(n721) );
  XNOR2_X1 U767 ( .A(n721), .B(n719), .ZN(n720) );
  NAND2_X1 U768 ( .A1(n720), .A2(n723), .ZN(n726) );
  XNOR2_X1 U769 ( .A(n721), .B(G227), .ZN(n722) );
  NOR2_X1 U770 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U771 ( .A1(G900), .A2(n724), .ZN(n725) );
  NAND2_X1 U772 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U773 ( .A(KEYINPUT126), .B(n727), .Z(G72) );
  XNOR2_X1 U774 ( .A(n728), .B(G119), .ZN(G21) );
  XOR2_X1 U775 ( .A(n729), .B(G122), .Z(G24) );
  XNOR2_X1 U776 ( .A(G140), .B(n730), .ZN(G42) );
  XNOR2_X1 U777 ( .A(G137), .B(KEYINPUT127), .ZN(n732) );
  XNOR2_X1 U778 ( .A(n732), .B(n731), .ZN(G39) );
  XOR2_X1 U779 ( .A(n733), .B(G131), .Z(G33) );
endmodule

