//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1297,
    new_n1298, new_n1299, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1357, new_n1358, new_n1359,
    new_n1360;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT65), .Z(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT0), .Z(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n209), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n203), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n214), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G107), .ZN(new_n223));
  INV_X1    g0023(.A(G264), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n226));
  INV_X1    g0026(.A(G58), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  INV_X1    g0028(.A(G97), .ZN(new_n229));
  INV_X1    g0029(.A(G257), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n226), .B1(new_n227), .B2(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n211), .B1(new_n225), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT66), .ZN(new_n233));
  INV_X1    g0033(.A(KEYINPUT1), .ZN(new_n234));
  OR2_X1    g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n233), .A2(new_n234), .ZN(new_n236));
  AND3_X1   g0036(.A1(new_n219), .A2(new_n235), .A3(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XOR2_X1   g0046(.A(G50), .B(G58), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(KEYINPUT73), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G1), .A3(G13), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G223), .A2(G1698), .ZN(new_n256));
  INV_X1    g0056(.A(G226), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n256), .B1(new_n257), .B2(G1698), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT72), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n261), .B1(new_n259), .B2(KEYINPUT3), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(KEYINPUT72), .A3(G33), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n258), .A2(new_n260), .A3(new_n262), .A4(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G87), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n255), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(new_n255), .A3(G274), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n255), .A2(G232), .A3(new_n268), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n267), .A2(G190), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n262), .A2(new_n260), .A3(new_n264), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n257), .A2(G1698), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n275), .B1(G223), .B2(G1698), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n266), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n255), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n270), .A2(new_n271), .ZN(new_n280));
  AOI21_X1  g0080(.A(G200), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n253), .B1(new_n273), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G200), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n283), .B1(new_n267), .B2(new_n272), .ZN(new_n284));
  INV_X1    g0084(.A(G190), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n279), .A2(new_n280), .A3(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(KEYINPUT73), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n289), .A2(KEYINPUT67), .B1(G1), .B2(G13), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT67), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n291), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n290), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT69), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n290), .A2(KEYINPUT69), .A3(new_n292), .A4(new_n293), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g0098(.A(KEYINPUT8), .B(G58), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n299), .B1(new_n208), .B2(G20), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n293), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n290), .A2(new_n292), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n263), .A2(G33), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n260), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT7), .B1(new_n308), .B2(new_n209), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT7), .ZN(new_n310));
  AOI211_X1 g0110(.A(new_n310), .B(G20), .C1(new_n260), .C2(new_n307), .ZN(new_n311));
  OAI21_X1  g0111(.A(G68), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G68), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n227), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(G20), .B1(new_n314), .B2(new_n202), .ZN(new_n315));
  NOR2_X1   g0115(.A1(G20), .A2(G33), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G159), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT16), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n306), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n274), .A2(new_n209), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT7), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n274), .A2(new_n310), .A3(new_n209), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n323), .A2(G68), .A3(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n325), .A2(KEYINPUT16), .A3(new_n318), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n304), .B1(new_n321), .B2(new_n326), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n288), .A2(KEYINPUT17), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT17), .B1(new_n288), .B2(new_n327), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n294), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n208), .A2(G20), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n331), .A2(G68), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT11), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n313), .A2(G20), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n209), .A2(G33), .ZN(new_n336));
  INV_X1    g0136(.A(new_n316), .ZN(new_n337));
  INV_X1    g0137(.A(G50), .ZN(new_n338));
  OAI221_X1 g0138(.A(new_n335), .B1(new_n336), .B2(new_n221), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n305), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n333), .B1(new_n334), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n334), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n302), .A2(new_n313), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n343), .B(KEYINPUT12), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT14), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT13), .ZN(new_n349));
  XNOR2_X1  g0149(.A(KEYINPUT3), .B(G33), .ZN(new_n350));
  INV_X1    g0150(.A(G1698), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n257), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n228), .A2(G1698), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n350), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(G33), .A2(G97), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n255), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n255), .A2(new_n268), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G274), .ZN(new_n360));
  INV_X1    g0160(.A(new_n215), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n360), .B1(new_n361), .B2(new_n254), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n359), .A2(G238), .B1(new_n362), .B2(new_n269), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n349), .B1(new_n357), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G238), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n270), .B1(new_n365), .B2(new_n358), .ZN(new_n366));
  NOR3_X1   g0166(.A1(new_n356), .A2(new_n366), .A3(KEYINPUT13), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n348), .B(G169), .C1(new_n364), .C2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n357), .A2(new_n349), .A3(new_n363), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT13), .B1(new_n356), .B2(new_n366), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n369), .A2(G179), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n369), .A2(new_n370), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n348), .B1(new_n373), .B2(G169), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n347), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(G200), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n376), .B(new_n346), .C1(new_n285), .C2(new_n373), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT18), .ZN(new_n380));
  OAI21_X1  g0180(.A(G169), .B1(new_n267), .B2(new_n272), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n279), .A2(new_n280), .A3(G179), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n380), .B1(new_n327), .B2(new_n384), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n298), .A2(new_n300), .B1(new_n302), .B2(new_n299), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n310), .B1(new_n350), .B2(G20), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n308), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n313), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n315), .A2(new_n317), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n320), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n305), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n318), .A2(KEYINPUT16), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n310), .B1(new_n274), .B2(new_n209), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n394), .A2(new_n313), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n393), .B1(new_n324), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n386), .B1(new_n392), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n397), .A2(KEYINPUT18), .A3(new_n383), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n385), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G20), .A2(G77), .ZN(new_n400));
  XNOR2_X1  g0200(.A(KEYINPUT15), .B(G87), .ZN(new_n401));
  OAI221_X1 g0201(.A(new_n400), .B1(new_n299), .B2(new_n337), .C1(new_n336), .C2(new_n401), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n402), .A2(new_n305), .B1(new_n221), .B2(new_n302), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n331), .A2(G77), .A3(new_n332), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n270), .B1(new_n222), .B2(new_n358), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n350), .A2(G238), .A3(G1698), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n350), .A2(G232), .A3(new_n351), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n407), .B(new_n408), .C1(new_n223), .C2(new_n350), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n406), .B1(new_n409), .B2(new_n278), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n405), .B1(G190), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(new_n283), .B2(new_n410), .ZN(new_n412));
  INV_X1    g0212(.A(G150), .ZN(new_n413));
  OAI22_X1  g0213(.A1(new_n299), .A2(new_n336), .B1(new_n413), .B2(new_n337), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT68), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT68), .ZN(new_n416));
  OAI221_X1 g0216(.A(new_n416), .B1(new_n337), .B2(new_n413), .C1(new_n299), .C2(new_n336), .ZN(new_n417));
  OAI21_X1  g0217(.A(G20), .B1(new_n201), .B2(new_n203), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n415), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n305), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n298), .A2(G50), .A3(new_n332), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n302), .A2(new_n338), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(G222), .A2(G1698), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n351), .A2(G223), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n350), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n426), .B(new_n278), .C1(G77), .C2(new_n350), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n359), .A2(G226), .B1(new_n362), .B2(new_n269), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(G179), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n423), .B(new_n431), .C1(G169), .C2(new_n429), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n410), .A2(new_n430), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n405), .B(new_n433), .C1(G169), .C2(new_n410), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n412), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n330), .A2(new_n379), .A3(new_n399), .A4(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT9), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT70), .B1(new_n423), .B2(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n429), .A2(new_n283), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n439), .B1(G190), .B2(new_n429), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n423), .A2(new_n437), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT71), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n420), .A2(new_n422), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT70), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n444), .A2(new_n445), .A3(KEYINPUT9), .A4(new_n421), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n442), .A2(new_n443), .A3(KEYINPUT10), .A4(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n446), .A2(new_n438), .A3(new_n440), .A4(new_n441), .ZN(new_n448));
  OR2_X1    g0248(.A1(new_n443), .A2(KEYINPUT10), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n443), .A2(KEYINPUT10), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n436), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT81), .ZN(new_n454));
  INV_X1    g0254(.A(G169), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n224), .A2(G1698), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(G257), .B2(G1698), .ZN(new_n457));
  INV_X1    g0257(.A(G303), .ZN(new_n458));
  OAI22_X1  g0258(.A1(new_n274), .A2(new_n457), .B1(new_n458), .B2(new_n350), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n278), .ZN(new_n460));
  XNOR2_X1  g0260(.A(KEYINPUT5), .B(G41), .ZN(new_n461));
  INV_X1    g0261(.A(G45), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(G1), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n461), .A2(new_n463), .B1(new_n361), .B2(new_n254), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n208), .A2(G45), .ZN(new_n465));
  NOR2_X1   g0265(.A1(KEYINPUT5), .A2(G41), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n464), .A2(G270), .B1(new_n362), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n455), .B1(new_n460), .B2(new_n470), .ZN(new_n471));
  AND2_X1   g0271(.A1(KEYINPUT5), .A2(G41), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n463), .B1(new_n472), .B2(new_n466), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(G270), .A3(new_n255), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n461), .A2(G274), .A3(new_n255), .A4(new_n463), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n476), .B1(new_n278), .B2(new_n459), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n471), .A2(KEYINPUT21), .B1(new_n477), .B2(G179), .ZN(new_n478));
  AOI21_X1  g0278(.A(G20), .B1(G33), .B2(G283), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n259), .A2(G97), .ZN(new_n480));
  INV_X1    g0280(.A(G116), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n479), .A2(new_n480), .B1(G20), .B2(new_n481), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n305), .A2(KEYINPUT20), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(KEYINPUT20), .B1(new_n305), .B2(new_n482), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n302), .A2(new_n481), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n208), .A2(G33), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n290), .A2(new_n292), .A3(new_n293), .A4(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n486), .B1(new_n488), .B2(new_n481), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n454), .B1(new_n478), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n460), .A2(new_n470), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(KEYINPUT21), .A3(G169), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n477), .A2(G179), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n490), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(KEYINPUT81), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n491), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT21), .ZN(new_n499));
  INV_X1    g0299(.A(new_n471), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n499), .B1(new_n500), .B2(new_n490), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n492), .A2(G200), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n490), .B(new_n502), .C1(new_n285), .C2(new_n492), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n498), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT77), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n351), .A2(KEYINPUT4), .A3(G244), .ZN(new_n507));
  INV_X1    g0307(.A(G283), .ZN(new_n508));
  OAI22_X1  g0308(.A1(new_n308), .A2(new_n507), .B1(new_n259), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT4), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n222), .A2(G1698), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n262), .A2(new_n264), .A3(new_n511), .A4(new_n260), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n509), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n260), .A2(new_n307), .A3(G250), .A4(G1698), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT75), .ZN(new_n515));
  XNOR2_X1  g0315(.A(new_n514), .B(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n255), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n473), .A2(G257), .A3(new_n255), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n475), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT76), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n518), .A2(KEYINPUT76), .A3(new_n475), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n455), .B1(new_n517), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT6), .ZN(new_n525));
  NOR3_X1   g0325(.A1(new_n525), .A2(new_n229), .A3(G107), .ZN(new_n526));
  XNOR2_X1  g0326(.A(G97), .B(G107), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n526), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  OAI22_X1  g0328(.A1(new_n528), .A2(new_n209), .B1(new_n221), .B2(new_n337), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n223), .B1(new_n387), .B2(new_n388), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n305), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n488), .A2(G97), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n293), .A2(new_n229), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n532), .A2(KEYINPUT74), .A3(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(KEYINPUT74), .B1(new_n532), .B2(new_n533), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n531), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n518), .A2(KEYINPUT76), .A3(new_n475), .ZN(new_n538));
  AOI21_X1  g0338(.A(KEYINPUT76), .B1(new_n518), .B2(new_n475), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g0340(.A(new_n514), .B(KEYINPUT75), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n512), .A2(new_n510), .ZN(new_n542));
  INV_X1    g0342(.A(new_n507), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n350), .A2(new_n543), .B1(G33), .B2(G283), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n278), .B1(new_n541), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n540), .A2(new_n546), .A3(new_n430), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n524), .A2(new_n537), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n540), .A2(new_n546), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n283), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n540), .A2(new_n546), .A3(new_n285), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n537), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n506), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n527), .A2(new_n525), .ZN(new_n554));
  INV_X1    g0354(.A(new_n526), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n556), .A2(G20), .B1(G77), .B2(new_n316), .ZN(new_n557));
  OAI21_X1  g0357(.A(G107), .B1(new_n309), .B2(new_n311), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n306), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n536), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n559), .B1(new_n560), .B2(new_n534), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n540), .A2(new_n546), .A3(new_n285), .ZN(new_n562));
  AOI21_X1  g0362(.A(G200), .B1(new_n540), .B2(new_n546), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n524), .A2(new_n537), .A3(new_n547), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(new_n565), .A3(KEYINPUT77), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n553), .A2(new_n566), .ZN(new_n567));
  AND2_X1   g0367(.A1(KEYINPUT83), .A2(KEYINPUT24), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT82), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n223), .A2(G20), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n569), .B1(new_n570), .B2(KEYINPUT23), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT23), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n572), .A2(new_n223), .A3(G20), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n209), .A2(G33), .A3(G116), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT22), .ZN(new_n577));
  INV_X1    g0377(.A(G87), .ZN(new_n578));
  NOR3_X1   g0378(.A1(new_n577), .A2(new_n578), .A3(G20), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n579), .A2(new_n260), .A3(new_n262), .A4(new_n264), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n578), .A2(G20), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n581), .A2(new_n260), .A3(new_n307), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n577), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n570), .A2(new_n569), .A3(KEYINPUT23), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n576), .A2(new_n580), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(KEYINPUT83), .A2(KEYINPUT24), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n584), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n588), .A2(new_n571), .A3(new_n575), .ZN(new_n589));
  INV_X1    g0389(.A(new_n586), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n589), .A2(new_n590), .A3(new_n580), .A4(new_n583), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n568), .B1(new_n587), .B2(new_n591), .ZN(new_n592));
  OR2_X1    g0392(.A1(new_n592), .A2(new_n306), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT84), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n293), .A2(G107), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT25), .ZN(new_n596));
  XNOR2_X1  g0396(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n488), .A2(new_n223), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n594), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  XNOR2_X1  g0399(.A(new_n595), .B(KEYINPUT25), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n600), .B(KEYINPUT84), .C1(new_n223), .C2(new_n488), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(G33), .A2(G294), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n230), .A2(G1698), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(G250), .B2(G1698), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n603), .B1(new_n274), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n278), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n464), .A2(G264), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n607), .A2(new_n475), .A3(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT85), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n606), .A2(new_n278), .B1(G264), .B2(new_n464), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n612), .A2(KEYINPUT85), .A3(new_n475), .ZN(new_n613));
  AOI21_X1  g0413(.A(G190), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n609), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n615), .A2(G200), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n593), .B(new_n602), .C1(new_n614), .C2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n611), .A2(G169), .A3(new_n613), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n615), .A2(G179), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n602), .B1(new_n592), .B2(new_n306), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT80), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n264), .A2(new_n260), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT79), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n313), .A2(G20), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n625), .A2(new_n626), .A3(new_n262), .A4(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n262), .A2(new_n264), .A3(new_n627), .A4(new_n260), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT79), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT19), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n355), .B2(new_n209), .ZN(new_n632));
  NOR4_X1   g0432(.A1(KEYINPUT78), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT78), .ZN(new_n634));
  NOR2_X1   g0434(.A1(G87), .A2(G97), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n634), .B1(new_n635), .B2(new_n223), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n632), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n631), .B1(new_n336), .B2(new_n229), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n628), .A2(new_n630), .A3(new_n637), .A4(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n305), .ZN(new_n640));
  INV_X1    g0440(.A(new_n401), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n641), .A2(new_n293), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n624), .B1(new_n640), .B2(new_n643), .ZN(new_n644));
  AOI211_X1 g0444(.A(KEYINPUT80), .B(new_n642), .C1(new_n639), .C2(new_n305), .ZN(new_n645));
  OAI22_X1  g0445(.A1(new_n644), .A2(new_n645), .B1(new_n401), .B2(new_n488), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n463), .A2(G250), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n465), .A2(G274), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n647), .A2(new_n278), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n222), .A2(G1698), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n650), .B1(G238), .B2(G1698), .ZN(new_n651));
  OAI22_X1  g0451(.A1(new_n274), .A2(new_n651), .B1(new_n259), .B2(new_n481), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n649), .B1(new_n652), .B2(new_n278), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n653), .A2(G169), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n654), .B1(new_n430), .B2(new_n653), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n646), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n653), .A2(new_n285), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(G200), .B2(new_n653), .ZN(new_n658));
  INV_X1    g0458(.A(new_n488), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G87), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n658), .B(new_n660), .C1(new_n644), .C2(new_n645), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n623), .A2(new_n662), .ZN(new_n663));
  AND4_X1   g0463(.A1(new_n453), .A2(new_n505), .A3(new_n567), .A4(new_n663), .ZN(G372));
  NAND2_X1  g0464(.A1(new_n375), .A2(new_n434), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n330), .A2(new_n377), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g0466(.A(KEYINPUT86), .B(KEYINPUT87), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n274), .A2(new_n310), .A3(new_n209), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n669), .A2(new_n394), .A3(new_n313), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n391), .B(new_n305), .C1(new_n670), .C2(new_n393), .ZN(new_n671));
  AOI221_X4 g0471(.A(new_n380), .B1(new_n381), .B2(new_n382), .C1(new_n671), .C2(new_n386), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT18), .B1(new_n397), .B2(new_n383), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n668), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n385), .A2(new_n398), .A3(new_n667), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n451), .B(new_n447), .C1(new_n666), .C2(new_n676), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n677), .A2(new_n432), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n488), .A2(new_n401), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n640), .A2(new_n643), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(KEYINPUT80), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n640), .A2(new_n624), .A3(new_n643), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n679), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n655), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n548), .B(new_n661), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT26), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n656), .A2(KEYINPUT26), .A3(new_n548), .A4(new_n661), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n564), .A2(new_n565), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n611), .A2(new_n613), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n285), .ZN(new_n692));
  INV_X1    g0492(.A(new_n616), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n621), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n681), .A2(new_n682), .B1(G87), .B2(new_n659), .ZN(new_n696));
  AOI22_X1  g0496(.A1(new_n696), .A2(new_n658), .B1(new_n646), .B2(new_n655), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n495), .A2(new_n496), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n622), .A2(new_n698), .A3(new_n501), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n695), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n689), .A2(new_n656), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n453), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n678), .B1(new_n702), .B2(new_n703), .ZN(G369));
  NAND2_X1  g0504(.A1(new_n698), .A2(new_n501), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n706), .A2(KEYINPUT27), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(KEYINPUT27), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(new_n708), .A3(G213), .ZN(new_n709));
  XOR2_X1   g0509(.A(KEYINPUT88), .B(G343), .Z(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n490), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n705), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n504), .B2(new_n713), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n715), .A2(KEYINPUT89), .A3(G330), .ZN(new_n716));
  AOI21_X1  g0516(.A(KEYINPUT89), .B1(new_n715), .B2(G330), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n623), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n621), .A2(new_n711), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n620), .A2(new_n621), .A3(new_n711), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n718), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n711), .B1(new_n498), .B2(new_n501), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(new_n622), .B2(new_n711), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g0527(.A(new_n727), .B(KEYINPUT90), .Z(G399));
  NOR3_X1   g0528(.A1(new_n633), .A2(new_n636), .A3(G116), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT91), .ZN(new_n730));
  INV_X1    g0530(.A(new_n212), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G41), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n730), .A2(G1), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(new_n217), .B2(new_n733), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT28), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT29), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n701), .A2(new_n737), .A3(new_n712), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n498), .A2(new_n501), .A3(new_n622), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n695), .A2(new_n739), .A3(new_n697), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n689), .A2(new_n656), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n737), .B1(new_n741), .B2(new_n712), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n477), .A2(G179), .A3(new_n612), .A4(new_n653), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT30), .ZN(new_n745));
  OR3_X1    g0545(.A1(new_n744), .A2(new_n549), .A3(new_n745), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n615), .A2(G179), .A3(new_n477), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT92), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n653), .B(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n747), .A2(new_n749), .A3(new_n549), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n745), .B1(new_n744), .B2(new_n549), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n746), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  AND3_X1   g0552(.A1(new_n752), .A2(KEYINPUT31), .A3(new_n711), .ZN(new_n753));
  AOI21_X1  g0553(.A(KEYINPUT31), .B1(new_n752), .B2(new_n711), .ZN(new_n754));
  OR3_X1    g0554(.A1(new_n753), .A2(new_n754), .A3(KEYINPUT93), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n663), .A2(new_n505), .A3(new_n567), .A4(new_n712), .ZN(new_n756));
  OAI21_X1  g0556(.A(KEYINPUT93), .B1(new_n753), .B2(new_n754), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G330), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n743), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n736), .B1(new_n761), .B2(G1), .ZN(G364));
  AND2_X1   g0562(.A1(new_n209), .A2(G13), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n208), .B1(new_n763), .B2(G45), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n732), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI211_X1 g0567(.A(new_n718), .B(new_n767), .C1(G330), .C2(new_n715), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n212), .A2(new_n350), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n769), .A2(new_n206), .B1(G116), .B2(new_n212), .ZN(new_n770));
  INV_X1    g0570(.A(new_n274), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n731), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(new_n462), .B2(new_n218), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n248), .A2(G45), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n770), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G13), .A2(G33), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n215), .B1(G20), .B2(new_n455), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n766), .B1(new_n776), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n209), .A2(new_n430), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G190), .A2(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n784), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n787), .A2(new_n285), .A3(G200), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n350), .B1(new_n221), .B2(new_n786), .C1(new_n789), .C2(new_n227), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n787), .A2(new_n285), .A3(new_n283), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(KEYINPUT94), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n791), .A2(KEYINPUT94), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n790), .B1(new_n796), .B2(G50), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n209), .A2(G179), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n798), .A2(G190), .A3(G200), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n578), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n798), .A2(new_n285), .A3(G200), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n800), .B1(G107), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n798), .A2(new_n785), .ZN(new_n804));
  INV_X1    g0604(.A(G159), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT32), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n797), .A2(new_n803), .A3(new_n807), .ZN(new_n808));
  NOR3_X1   g0608(.A1(new_n285), .A2(G179), .A3(G200), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n209), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(new_n229), .ZN(new_n811));
  NOR3_X1   g0611(.A1(new_n787), .A2(new_n283), .A3(G190), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n811), .B1(G68), .B2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT95), .Z(new_n814));
  NAND2_X1  g0614(.A1(new_n796), .A2(G326), .ZN(new_n815));
  INV_X1    g0615(.A(new_n786), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n788), .A2(G322), .B1(G311), .B2(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(KEYINPUT33), .B(G317), .ZN(new_n818));
  INV_X1    g0618(.A(new_n804), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n812), .A2(new_n818), .B1(G329), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n810), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n821), .A2(G294), .B1(new_n802), .B2(G283), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n815), .A2(new_n817), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n308), .B1(new_n799), .B2(new_n458), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT96), .Z(new_n825));
  OAI22_X1  g0625(.A1(new_n808), .A2(new_n814), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n826), .A2(KEYINPUT97), .ZN(new_n827));
  INV_X1    g0627(.A(new_n780), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(new_n826), .B2(KEYINPUT97), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n783), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n779), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n830), .B1(new_n715), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n768), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(G396));
  NAND2_X1  g0634(.A1(new_n405), .A2(new_n711), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n412), .A2(new_n434), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(KEYINPUT99), .B1(new_n434), .B2(new_n712), .ZN(new_n837));
  INV_X1    g0637(.A(new_n410), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n838), .A2(new_n455), .B1(new_n404), .B2(new_n403), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT99), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n839), .A2(new_n840), .A3(new_n433), .A4(new_n711), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n836), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(new_n701), .B2(new_n712), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n712), .ZN(new_n845));
  INV_X1    g0645(.A(new_n656), .ZN(new_n846));
  NOR3_X1   g0646(.A1(new_n662), .A2(new_n690), .A3(new_n694), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n846), .B1(new_n847), .B2(new_n699), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n845), .B1(new_n848), .B2(new_n689), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n850), .A2(new_n759), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n766), .B1(new_n850), .B2(new_n759), .ZN(new_n853));
  INV_X1    g0653(.A(G137), .ZN(new_n854));
  INV_X1    g0654(.A(new_n812), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n795), .A2(new_n854), .B1(new_n413), .B2(new_n855), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT98), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n788), .A2(G143), .B1(G159), .B2(new_n816), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT34), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n274), .B1(new_n819), .B2(G132), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n810), .A2(new_n227), .B1(new_n799), .B2(new_n338), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(G68), .B2(new_n802), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n860), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n796), .A2(G303), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n350), .B(new_n811), .C1(G283), .C2(new_n812), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n801), .A2(new_n578), .ZN(new_n867));
  INV_X1    g0667(.A(new_n799), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n867), .B1(G107), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(G311), .ZN(new_n870));
  OAI22_X1  g0670(.A1(new_n786), .A2(new_n481), .B1(new_n804), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(G294), .B2(new_n788), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n865), .A2(new_n866), .A3(new_n869), .A4(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n828), .B1(new_n864), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n780), .A2(new_n777), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n767), .B(new_n874), .C1(new_n221), .C2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n843), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n777), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n852), .A2(new_n853), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(G384));
  OR2_X1    g0680(.A1(new_n556), .A2(KEYINPUT35), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n556), .A2(KEYINPUT35), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n881), .A2(G116), .A3(new_n216), .A4(new_n882), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n883), .B(KEYINPUT36), .Z(new_n884));
  OR3_X1    g0684(.A1(new_n217), .A2(new_n221), .A3(new_n314), .ZN(new_n885));
  INV_X1    g0685(.A(new_n201), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(G68), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n208), .B(G13), .C1(new_n885), .C2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n434), .A2(new_n711), .ZN(new_n890));
  INV_X1    g0690(.A(new_n845), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n890), .B1(new_n701), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n347), .A2(new_n711), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n375), .A2(new_n377), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n893), .B1(new_n375), .B2(new_n377), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT38), .ZN(new_n898));
  NOR3_X1   g0698(.A1(new_n273), .A2(new_n281), .A3(new_n253), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT73), .B1(new_n284), .B2(new_n286), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n671), .B(new_n386), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n305), .B1(new_n670), .B2(new_n393), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT16), .B1(new_n325), .B2(new_n318), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n386), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n709), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n904), .A2(new_n383), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n901), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT37), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n709), .B1(new_n671), .B2(new_n386), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n327), .B2(new_n288), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT37), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n397), .A2(new_n383), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n909), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n906), .B1(new_n330), .B2(new_n399), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n898), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n906), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT17), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n901), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n288), .A2(KEYINPUT17), .A3(new_n327), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n672), .A2(new_n673), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n918), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n909), .A2(new_n914), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n924), .A2(new_n925), .A3(KEYINPUT38), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n917), .A2(new_n926), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n897), .A2(new_n927), .B1(new_n676), .B2(new_n709), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n924), .A2(KEYINPUT38), .A3(new_n925), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT38), .B1(new_n924), .B2(new_n925), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT39), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT101), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n927), .A2(KEYINPUT101), .A3(KEYINPUT39), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT39), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n674), .A2(new_n675), .A3(new_n920), .A4(new_n921), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n910), .ZN(new_n937));
  INV_X1    g0737(.A(new_n910), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n901), .A2(new_n938), .A3(new_n913), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT102), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n911), .A2(KEYINPUT102), .A3(new_n913), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT86), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n901), .A2(new_n938), .A3(new_n943), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n941), .A2(new_n942), .A3(KEYINPUT37), .A4(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(KEYINPUT37), .ZN(new_n946));
  AOI21_X1  g0746(.A(KEYINPUT102), .B1(new_n911), .B2(new_n913), .ZN(new_n947));
  AND4_X1   g0747(.A1(KEYINPUT102), .A2(new_n901), .A3(new_n938), .A4(new_n913), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n937), .A2(new_n945), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n929), .B1(new_n950), .B2(new_n898), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n933), .A2(new_n934), .B1(new_n935), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT100), .ZN(new_n953));
  OR3_X1    g0753(.A1(new_n375), .A2(new_n953), .A3(new_n711), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n953), .B1(new_n375), .B2(new_n711), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n928), .B1(new_n952), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n453), .B1(new_n738), .B2(new_n742), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n678), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n957), .B(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n950), .A2(new_n898), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n926), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT40), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n843), .B1(new_n894), .B2(new_n895), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n753), .A2(new_n754), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n963), .B(new_n964), .C1(new_n756), .C2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n756), .A2(new_n965), .ZN(new_n967));
  INV_X1    g0767(.A(new_n964), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n967), .B(new_n968), .C1(new_n929), .C2(new_n930), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n962), .A2(new_n966), .B1(new_n969), .B2(new_n963), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n970), .A2(new_n453), .A3(new_n967), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(G330), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n970), .B1(new_n453), .B2(new_n967), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n960), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n208), .B2(new_n763), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n960), .A2(new_n974), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n889), .B1(new_n976), .B2(new_n977), .ZN(G367));
  NOR2_X1   g0778(.A1(new_n561), .A2(new_n712), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n690), .A2(new_n979), .B1(new_n565), .B2(new_n712), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT103), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n981), .A2(new_n719), .A3(new_n724), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT42), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n981), .A2(new_n621), .A3(new_n620), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n711), .B1(new_n984), .B2(new_n565), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT43), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n696), .A2(new_n712), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n662), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(new_n846), .B2(new_n988), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n986), .A2(new_n987), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n987), .ZN(new_n992));
  INV_X1    g0792(.A(new_n990), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n992), .B(new_n994), .C1(new_n983), .C2(new_n985), .ZN(new_n995));
  AND4_X1   g0795(.A1(new_n723), .A2(new_n991), .A3(new_n981), .A4(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n991), .A2(new_n995), .B1(new_n723), .B2(new_n981), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n732), .B(KEYINPUT41), .Z(new_n999));
  INV_X1    g0799(.A(new_n981), .ZN(new_n1000));
  AOI21_X1  g0800(.A(KEYINPUT44), .B1(new_n1000), .B2(new_n726), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n726), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT44), .ZN(new_n1003));
  NOR3_X1   g0803(.A1(new_n1002), .A2(new_n981), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT45), .ZN(new_n1005));
  NOR3_X1   g0805(.A1(new_n1000), .A2(new_n1005), .A3(new_n726), .ZN(new_n1006));
  AOI21_X1  g0806(.A(KEYINPUT45), .B1(new_n1002), .B2(new_n981), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n1001), .A2(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT104), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n723), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1008), .B(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n761), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n721), .A2(new_n722), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n725), .B1(new_n1013), .B2(new_n724), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n718), .B(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(KEYINPUT105), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1015), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT105), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1017), .A2(new_n761), .A3(new_n1018), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1011), .A2(new_n1016), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n999), .B1(new_n1020), .B2(new_n761), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n998), .B1(new_n1021), .B2(new_n765), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n781), .B1(new_n212), .B2(new_n401), .C1(new_n773), .C2(new_n244), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n796), .A2(G143), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n350), .B1(new_n789), .B2(new_n413), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G58), .B2(new_n868), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n801), .A2(new_n221), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(G68), .B2(new_n821), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n886), .A2(new_n786), .B1(new_n804), .B2(new_n854), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(G159), .B2(new_n812), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1024), .A2(new_n1026), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n795), .A2(new_n870), .B1(new_n458), .B2(new_n789), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT106), .Z(new_n1033));
  AOI22_X1  g0833(.A1(new_n812), .A2(G294), .B1(G283), .B2(new_n816), .ZN(new_n1034));
  INV_X1    g0834(.A(G317), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1034), .B1(new_n1035), .B2(new_n804), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n799), .A2(new_n481), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1036), .B1(KEYINPUT46), .B2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n801), .A2(new_n229), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n771), .B(new_n1039), .C1(G107), .C2(new_n821), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1038), .B(new_n1040), .C1(KEYINPUT46), .C2(new_n1037), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1031), .B1(new_n1033), .B2(new_n1041), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT47), .Z(new_n1043));
  OAI211_X1 g0843(.A(new_n766), .B(new_n1023), .C1(new_n1043), .C2(new_n828), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT107), .Z(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n831), .B2(new_n993), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1022), .A2(new_n1046), .ZN(G387));
  INV_X1    g0847(.A(KEYINPUT110), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n732), .B(KEYINPUT109), .Z(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n1017), .B2(new_n761), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1017), .A2(new_n765), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n772), .B1(new_n241), .B2(new_n462), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n730), .B2(new_n769), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n299), .A2(G50), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT50), .ZN(new_n1056));
  AOI21_X1  g0856(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n730), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1054), .A2(new_n1058), .B1(new_n223), .B2(new_n731), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n766), .B1(new_n1059), .B2(new_n782), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n812), .A2(G311), .B1(G303), .B2(new_n816), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n1035), .B2(new_n789), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n796), .B2(G322), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1063), .A2(KEYINPUT48), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(KEYINPUT48), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n821), .A2(G283), .B1(new_n868), .B2(G294), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT49), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n801), .A2(new_n481), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n771), .B(new_n1071), .C1(G326), .C2(new_n819), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1069), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n795), .A2(new_n805), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1039), .A2(new_n274), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n821), .A2(new_n641), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1075), .B(new_n1076), .C1(new_n221), .C2(new_n799), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n786), .A2(new_n313), .B1(new_n804), .B2(new_n413), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n338), .A2(new_n789), .B1(new_n855), .B2(new_n299), .ZN(new_n1079));
  NOR4_X1   g0879(.A1(new_n1074), .A2(new_n1077), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT108), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1073), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1060), .B1(new_n1082), .B2(new_n780), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n1013), .B2(new_n831), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1052), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1048), .B1(new_n1051), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n1051), .A2(new_n1048), .A3(new_n1085), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(G393));
  OAI22_X1  g0890(.A1(new_n795), .A2(new_n413), .B1(new_n805), .B2(new_n789), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT51), .Z(new_n1092));
  NAND2_X1  g0892(.A1(new_n819), .A2(G143), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1093), .B1(new_n299), .B2(new_n786), .C1(new_n855), .C2(new_n886), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n810), .A2(new_n221), .B1(new_n799), .B2(new_n313), .ZN(new_n1095));
  OR4_X1    g0895(.A1(new_n274), .A2(new_n1094), .A3(new_n867), .A4(new_n1095), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n795), .A2(new_n1035), .B1(new_n870), .B2(new_n789), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT52), .Z(new_n1098));
  AOI22_X1  g0898(.A1(new_n812), .A2(G303), .B1(G294), .B2(new_n816), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n481), .B2(new_n810), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT112), .Z(new_n1101));
  AOI21_X1  g0901(.A(new_n350), .B1(new_n819), .B2(G322), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1102), .B1(new_n223), .B2(new_n801), .C1(new_n508), .C2(new_n799), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n1103), .A2(KEYINPUT111), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(KEYINPUT111), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1101), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1092), .A2(new_n1096), .B1(new_n1098), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n780), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n772), .A2(new_n251), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n782), .B1(G97), .B2(new_n731), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n767), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1108), .B(new_n1111), .C1(new_n981), .C2(new_n831), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1008), .B(new_n723), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1112), .B1(new_n1113), .B2(new_n764), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n1020), .A2(new_n1049), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n1113), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1114), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(G390));
  NAND2_X1  g0919(.A1(new_n967), .A2(G330), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n896), .B1(new_n1120), .B2(new_n877), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n896), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n758), .A2(G330), .A3(new_n843), .A4(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n741), .A2(new_n712), .A3(new_n843), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n890), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1121), .A2(new_n1123), .A3(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1120), .A2(new_n964), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n758), .A2(G330), .A3(new_n843), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1128), .B1(new_n1129), .B2(new_n896), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1127), .B1(new_n1130), .B2(new_n892), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1120), .A2(new_n703), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n959), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n951), .A2(new_n935), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n956), .B1(new_n892), .B2(new_n896), .ZN(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT101), .B1(new_n927), .B2(KEYINPUT39), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n932), .B(new_n935), .C1(new_n917), .C2(new_n926), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1135), .B(new_n1136), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT113), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n954), .A2(new_n1140), .A3(new_n955), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1140), .B1(new_n954), .B2(new_n955), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n962), .B(new_n1144), .C1(new_n1126), .C2(new_n896), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1139), .A2(new_n1145), .A3(new_n1123), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1139), .A2(new_n1145), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n1128), .ZN(new_n1148));
  AND4_X1   g0948(.A1(KEYINPUT114), .A2(new_n1134), .A3(new_n1146), .A4(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(KEYINPUT114), .A2(new_n1134), .B1(new_n1148), .B2(new_n1146), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1049), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1148), .A2(new_n765), .A3(new_n1146), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n767), .B1(new_n299), .B2(new_n875), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT54), .B(G143), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n812), .A2(G137), .B1(new_n816), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(G132), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1156), .B1(new_n1157), .B2(new_n789), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n796), .B2(G128), .ZN(new_n1159));
  INV_X1    g0959(.A(G125), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n350), .B1(new_n804), .B2(new_n1160), .C1(new_n810), .C2(new_n805), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n201), .B2(new_n802), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n799), .A2(new_n413), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1163), .B(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1159), .A2(new_n1162), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n796), .A2(G283), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n350), .B(new_n800), .C1(G107), .C2(new_n812), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n821), .A2(G77), .B1(new_n802), .B2(G68), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n789), .A2(new_n481), .B1(new_n786), .B2(new_n229), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(G294), .B2(new_n819), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .A4(new_n1171), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1166), .A2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1135), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1153), .B1(new_n828), .B2(new_n1173), .C1(new_n1174), .C2(new_n778), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n1152), .A2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1176), .A2(KEYINPUT116), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1152), .A2(KEYINPUT116), .A3(new_n1175), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1151), .B1(new_n1177), .B2(new_n1178), .ZN(G378));
  INV_X1    g0979(.A(KEYINPUT118), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n447), .A2(new_n451), .A3(new_n432), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n423), .A2(new_n905), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n447), .A2(new_n451), .A3(new_n432), .A4(new_n1182), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1186), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1180), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1189), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1191), .A2(KEYINPUT118), .A3(new_n1187), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n777), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n795), .A2(new_n481), .B1(new_n313), .B2(new_n810), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT117), .ZN(new_n1196));
  OR2_X1    g0996(.A1(new_n771), .A2(G41), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n641), .A2(new_n816), .B1(new_n819), .B2(G283), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1198), .B1(new_n789), .B2(new_n223), .C1(new_n229), .C2(new_n855), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n799), .A2(new_n221), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n801), .A2(new_n227), .ZN(new_n1201));
  OR3_X1    g1001(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  NOR3_X1   g1002(.A1(new_n1196), .A2(new_n1197), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(KEYINPUT58), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1197), .B(new_n338), .C1(G33), .C2(G41), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n855), .A2(new_n1157), .B1(new_n786), .B2(new_n854), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G128), .B2(new_n788), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n821), .A2(G150), .B1(new_n868), .B2(new_n1155), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1208), .B(new_n1209), .C1(new_n1160), .C2(new_n795), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1210), .A2(KEYINPUT59), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(KEYINPUT59), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n802), .A2(G159), .ZN(new_n1213));
  AOI211_X1 g1013(.A(G33), .B(G41), .C1(new_n819), .C2(G124), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n1203), .A2(KEYINPUT58), .B1(new_n1211), .B2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n780), .B1(new_n1206), .B2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n767), .B1(new_n886), .B2(new_n875), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1194), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n941), .A2(new_n942), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n946), .A2(new_n1221), .B1(new_n936), .B2(new_n910), .ZN(new_n1222));
  AOI21_X1  g1022(.A(KEYINPUT38), .B1(new_n1222), .B2(new_n945), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n966), .B1(new_n1223), .B2(new_n929), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n969), .A2(new_n963), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1224), .A2(new_n1225), .A3(G330), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1226), .A2(new_n1193), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n970), .B2(G330), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n957), .B1(new_n1227), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n676), .A2(new_n709), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1122), .B1(new_n849), .B2(new_n890), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n927), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1232), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n956), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1235), .B1(new_n1174), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n970), .A2(G330), .A3(new_n1192), .A4(new_n1190), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT119), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1231), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  OAI211_X1 g1042(.A(KEYINPUT119), .B(new_n957), .C1(new_n1227), .C2(new_n1230), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1220), .B1(new_n1244), .B2(new_n765), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n896), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(new_n1247), .A2(new_n951), .A3(new_n1143), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n952), .B2(new_n1136), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1128), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1131), .B(new_n1146), .C1(new_n1249), .C2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1133), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1252), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1049), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT57), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(new_n1231), .B2(new_n1240), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1254), .B1(new_n1256), .B2(new_n1252), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n1253), .A2(KEYINPUT57), .B1(new_n1257), .B2(KEYINPUT120), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1257), .A2(KEYINPUT120), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1246), .B1(new_n1259), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(G375));
  OR2_X1    g1063(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n999), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1264), .A2(new_n1265), .A3(new_n1134), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n896), .A2(new_n777), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n780), .A2(G68), .A3(new_n777), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(G107), .A2(new_n816), .B1(new_n819), .B2(G303), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n508), .B2(new_n789), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n350), .B(new_n1027), .C1(G116), .C2(new_n812), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1271), .B(new_n1076), .C1(new_n229), .C2(new_n799), .ZN(new_n1272));
  AOI211_X1 g1072(.A(new_n1270), .B(new_n1272), .C1(G294), .C2(new_n796), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT121), .ZN(new_n1274));
  OR2_X1    g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n786), .A2(new_n413), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n854), .A2(new_n789), .B1(new_n855), .B2(new_n1154), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n1277), .B(new_n1278), .C1(G128), .C2(new_n819), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1201), .A2(new_n274), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1280), .B(KEYINPUT122), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n796), .A2(G132), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n821), .A2(G50), .B1(new_n868), .B2(G159), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1279), .A2(new_n1281), .A3(new_n1282), .A4(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1275), .A2(new_n1276), .A3(new_n1284), .ZN(new_n1285));
  AOI211_X1 g1085(.A(new_n767), .B(new_n1268), .C1(new_n1285), .C2(new_n780), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(new_n1131), .A2(new_n765), .B1(new_n1267), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1266), .A2(new_n1287), .ZN(G381));
  AND3_X1   g1088(.A1(new_n1118), .A2(new_n1022), .A3(new_n1046), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1151), .A2(new_n1176), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  OR3_X1    g1091(.A1(new_n1051), .A2(new_n1048), .A3(new_n1085), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(new_n1086), .A3(new_n833), .ZN(new_n1293));
  NOR3_X1   g1093(.A1(new_n1293), .A2(G384), .A3(G381), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1262), .A2(new_n1289), .A3(new_n1291), .A4(new_n1294), .ZN(new_n1295));
  XOR2_X1   g1095(.A(new_n1295), .B(KEYINPUT123), .Z(G407));
  NAND2_X1  g1096(.A1(new_n710), .A2(G213), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1262), .A2(new_n1291), .A3(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(G407), .A2(G213), .A3(new_n1299), .ZN(G409));
  OAI211_X1 g1100(.A(G378), .B(new_n1245), .C1(new_n1258), .C2(new_n1260), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT125), .ZN(new_n1302));
  AND2_X1   g1102(.A1(new_n1231), .A2(new_n1240), .ZN(new_n1303));
  OAI211_X1 g1103(.A(new_n1302), .B(new_n1219), .C1(new_n1303), .C2(new_n764), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n764), .B1(new_n1231), .B2(new_n1240), .ZN(new_n1305));
  OAI21_X1  g1105(.A(KEYINPUT125), .B1(new_n1305), .B2(new_n1220), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1252), .A2(new_n1242), .A3(new_n1265), .A4(new_n1243), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT124), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1304), .B(new_n1306), .C1(new_n1307), .C2(new_n1308), .ZN(new_n1309));
  AND2_X1   g1109(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1291), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1301), .A2(new_n1311), .ZN(new_n1312));
  AND2_X1   g1112(.A1(new_n1264), .A2(KEYINPUT60), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1264), .A2(KEYINPUT60), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1049), .B(new_n1134), .C1(new_n1313), .C2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n1287), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n879), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1315), .A2(G384), .A3(new_n1287), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1312), .A2(new_n1297), .A3(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(KEYINPUT62), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1312), .A2(new_n1297), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1298), .A2(G2897), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1319), .A2(new_n1324), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1317), .A2(G2897), .A3(new_n1298), .A4(new_n1318), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1323), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT61), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1298), .B1(new_n1301), .B2(new_n1311), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT62), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1330), .A2(new_n1331), .A3(new_n1320), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1322), .A2(new_n1328), .A3(new_n1329), .A4(new_n1332), .ZN(new_n1333));
  NOR3_X1   g1133(.A1(new_n1087), .A2(new_n1088), .A3(G396), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n833), .B1(new_n1292), .B2(new_n1086), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1118), .B1(new_n1022), .B2(new_n1046), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1336), .B1(new_n1289), .B2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(G387), .A2(G390), .ZN(new_n1339));
  OAI21_X1  g1139(.A(G396), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(new_n1293), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1118), .A2(new_n1022), .A3(new_n1046), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1339), .A2(new_n1341), .A3(new_n1342), .ZN(new_n1343));
  AND3_X1   g1143(.A1(new_n1338), .A2(KEYINPUT127), .A3(new_n1343), .ZN(new_n1344));
  AOI21_X1  g1144(.A(KEYINPUT127), .B1(new_n1338), .B2(new_n1343), .ZN(new_n1345));
  NOR2_X1   g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1333), .A2(new_n1346), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1338), .A2(new_n1343), .A3(new_n1329), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT63), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1348), .B1(new_n1321), .B2(new_n1349), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1330), .A2(KEYINPUT63), .A3(new_n1320), .ZN(new_n1351));
  NOR2_X1   g1151(.A1(new_n1323), .A2(KEYINPUT126), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT126), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1327), .B1(new_n1330), .B2(new_n1353), .ZN(new_n1354));
  OAI211_X1 g1154(.A(new_n1350), .B(new_n1351), .C1(new_n1352), .C2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1347), .A2(new_n1355), .ZN(G405));
  OAI21_X1  g1156(.A(new_n1301), .B1(new_n1262), .B2(new_n1290), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1357), .A2(new_n1320), .ZN(new_n1358));
  OAI211_X1 g1158(.A(new_n1301), .B(new_n1319), .C1(new_n1262), .C2(new_n1290), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1358), .A2(new_n1359), .ZN(new_n1360));
  XNOR2_X1  g1160(.A(new_n1360), .B(new_n1346), .ZN(G402));
endmodule


