

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591;

  XNOR2_X1 U327 ( .A(n382), .B(n416), .ZN(n383) );
  INV_X1 U328 ( .A(n542), .ZN(n406) );
  AND2_X1 U329 ( .A1(n408), .A2(n407), .ZN(n409) );
  XNOR2_X1 U330 ( .A(n343), .B(KEYINPUT9), .ZN(n344) );
  XNOR2_X1 U331 ( .A(n345), .B(n344), .ZN(n350) );
  XNOR2_X1 U332 ( .A(n384), .B(n383), .ZN(n404) );
  XOR2_X1 U333 ( .A(KEYINPUT121), .B(n453), .Z(n572) );
  XNOR2_X1 U334 ( .A(n351), .B(n562), .ZN(n547) );
  XNOR2_X1 U335 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n454) );
  XOR2_X1 U336 ( .A(G43GAT), .B(G134GAT), .Z(n330) );
  XOR2_X1 U337 ( .A(G15GAT), .B(G127GAT), .Z(n363) );
  XNOR2_X1 U338 ( .A(n330), .B(n363), .ZN(n296) );
  XNOR2_X1 U339 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n295) );
  XNOR2_X1 U340 ( .A(n295), .B(KEYINPUT79), .ZN(n443) );
  XNOR2_X1 U341 ( .A(n296), .B(n443), .ZN(n297) );
  XOR2_X1 U342 ( .A(G120GAT), .B(G71GAT), .Z(n382) );
  XOR2_X1 U343 ( .A(n297), .B(n382), .Z(n299) );
  XNOR2_X1 U344 ( .A(G190GAT), .B(G99GAT), .ZN(n298) );
  XNOR2_X1 U345 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U346 ( .A(KEYINPUT20), .B(KEYINPUT81), .Z(n301) );
  NAND2_X1 U347 ( .A1(G227GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U348 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U349 ( .A(n303), .B(n302), .Z(n310) );
  XOR2_X1 U350 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n305) );
  XNOR2_X1 U351 ( .A(KEYINPUT82), .B(KEYINPUT17), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U353 ( .A(n306), .B(G183GAT), .Z(n308) );
  XNOR2_X1 U354 ( .A(G169GAT), .B(G176GAT), .ZN(n307) );
  XNOR2_X1 U355 ( .A(n308), .B(n307), .ZN(n426) );
  XNOR2_X1 U356 ( .A(n426), .B(KEYINPUT80), .ZN(n309) );
  XNOR2_X1 U357 ( .A(n310), .B(n309), .ZN(n534) );
  XNOR2_X1 U358 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n311) );
  XNOR2_X1 U359 ( .A(n311), .B(G211GAT), .ZN(n413) );
  XOR2_X1 U360 ( .A(G22GAT), .B(G155GAT), .Z(n353) );
  XOR2_X1 U361 ( .A(n413), .B(n353), .Z(n313) );
  XNOR2_X1 U362 ( .A(G106GAT), .B(KEYINPUT84), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n328) );
  XOR2_X1 U364 ( .A(G162GAT), .B(KEYINPUT70), .Z(n315) );
  XNOR2_X1 U365 ( .A(G50GAT), .B(G218GAT), .ZN(n314) );
  XNOR2_X1 U366 ( .A(n315), .B(n314), .ZN(n348) );
  XOR2_X1 U367 ( .A(n348), .B(G204GAT), .Z(n317) );
  NAND2_X1 U368 ( .A1(G228GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U369 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U370 ( .A(KEYINPUT86), .B(KEYINPUT23), .Z(n319) );
  XNOR2_X1 U371 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U373 ( .A(n321), .B(n320), .Z(n326) );
  XOR2_X1 U374 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n323) );
  XNOR2_X1 U375 ( .A(G141GAT), .B(KEYINPUT85), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n430) );
  XNOR2_X1 U377 ( .A(G78GAT), .B(KEYINPUT67), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n324), .B(G148GAT), .ZN(n373) );
  XNOR2_X1 U379 ( .A(n430), .B(n373), .ZN(n325) );
  XNOR2_X1 U380 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U381 ( .A(n328), .B(n327), .Z(n466) );
  INV_X1 U382 ( .A(KEYINPUT75), .ZN(n351) );
  XOR2_X1 U383 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n329) );
  XNOR2_X1 U384 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U385 ( .A(G36GAT), .B(G190GAT), .Z(n422) );
  XNOR2_X1 U386 ( .A(n331), .B(n422), .ZN(n337) );
  INV_X1 U387 ( .A(n337), .ZN(n335) );
  XOR2_X1 U388 ( .A(KEYINPUT73), .B(KEYINPUT10), .Z(n333) );
  XNOR2_X1 U389 ( .A(KEYINPUT65), .B(KEYINPUT71), .ZN(n332) );
  XOR2_X1 U390 ( .A(n333), .B(n332), .Z(n336) );
  INV_X1 U391 ( .A(n336), .ZN(n334) );
  NAND2_X1 U392 ( .A1(n335), .A2(n334), .ZN(n339) );
  NAND2_X1 U393 ( .A1(n337), .A2(n336), .ZN(n338) );
  NAND2_X1 U394 ( .A1(n339), .A2(n338), .ZN(n341) );
  NAND2_X1 U395 ( .A1(G232GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U396 ( .A(n341), .B(n340), .ZN(n345) );
  XNOR2_X1 U397 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n342) );
  XNOR2_X1 U398 ( .A(n342), .B(KEYINPUT8), .ZN(n391) );
  XOR2_X1 U399 ( .A(n391), .B(KEYINPUT74), .Z(n343) );
  XOR2_X1 U400 ( .A(G92GAT), .B(G85GAT), .Z(n347) );
  XNOR2_X1 U401 ( .A(G99GAT), .B(G106GAT), .ZN(n346) );
  XNOR2_X1 U402 ( .A(n347), .B(n346), .ZN(n374) );
  XOR2_X1 U403 ( .A(n348), .B(n374), .Z(n349) );
  XNOR2_X1 U404 ( .A(n350), .B(n349), .ZN(n562) );
  XNOR2_X1 U405 ( .A(KEYINPUT36), .B(n547), .ZN(n586) );
  XNOR2_X1 U406 ( .A(G183GAT), .B(G71GAT), .ZN(n352) );
  XNOR2_X1 U407 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n377) );
  XNOR2_X1 U408 ( .A(n352), .B(n377), .ZN(n367) );
  XOR2_X1 U409 ( .A(G8GAT), .B(KEYINPUT76), .Z(n421) );
  XOR2_X1 U410 ( .A(n421), .B(n353), .Z(n355) );
  NAND2_X1 U411 ( .A1(G231GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U412 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U413 ( .A(KEYINPUT77), .B(KEYINPUT15), .Z(n357) );
  XNOR2_X1 U414 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n356) );
  XNOR2_X1 U415 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U416 ( .A(n359), .B(n358), .Z(n365) );
  XOR2_X1 U417 ( .A(G64GAT), .B(G211GAT), .Z(n361) );
  XNOR2_X1 U418 ( .A(G1GAT), .B(G78GAT), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U420 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U422 ( .A(n367), .B(n366), .ZN(n542) );
  NAND2_X1 U423 ( .A1(n586), .A2(n406), .ZN(n369) );
  XOR2_X1 U424 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n368) );
  XNOR2_X1 U425 ( .A(n369), .B(n368), .ZN(n385) );
  XOR2_X1 U426 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n371) );
  NAND2_X1 U427 ( .A1(G230GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U428 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U429 ( .A(n372), .B(KEYINPUT32), .Z(n376) );
  XNOR2_X1 U430 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U431 ( .A(n376), .B(n375), .ZN(n379) );
  INV_X1 U432 ( .A(n377), .ZN(n378) );
  XNOR2_X1 U433 ( .A(n379), .B(n378), .ZN(n381) );
  XOR2_X1 U434 ( .A(G176GAT), .B(KEYINPUT68), .Z(n380) );
  XNOR2_X1 U435 ( .A(n381), .B(n380), .ZN(n384) );
  XNOR2_X1 U436 ( .A(G204GAT), .B(G64GAT), .ZN(n416) );
  NAND2_X1 U437 ( .A1(n385), .A2(n404), .ZN(n386) );
  XNOR2_X1 U438 ( .A(n386), .B(KEYINPUT113), .ZN(n403) );
  XOR2_X1 U439 ( .A(G113GAT), .B(G15GAT), .Z(n388) );
  XNOR2_X1 U440 ( .A(G169GAT), .B(G50GAT), .ZN(n387) );
  XNOR2_X1 U441 ( .A(n388), .B(n387), .ZN(n402) );
  XOR2_X1 U442 ( .A(G43GAT), .B(G36GAT), .Z(n390) );
  NAND2_X1 U443 ( .A1(G229GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U444 ( .A(n390), .B(n389), .ZN(n392) );
  XOR2_X1 U445 ( .A(n392), .B(n391), .Z(n400) );
  XOR2_X1 U446 ( .A(G1GAT), .B(G197GAT), .Z(n394) );
  XNOR2_X1 U447 ( .A(G141GAT), .B(G22GAT), .ZN(n393) );
  XNOR2_X1 U448 ( .A(n394), .B(n393), .ZN(n398) );
  XOR2_X1 U449 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n396) );
  XNOR2_X1 U450 ( .A(G8GAT), .B(KEYINPUT30), .ZN(n395) );
  XNOR2_X1 U451 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U452 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U453 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U454 ( .A(n402), .B(n401), .ZN(n578) );
  INV_X1 U455 ( .A(n578), .ZN(n536) );
  NAND2_X1 U456 ( .A1(n403), .A2(n536), .ZN(n411) );
  XOR2_X1 U457 ( .A(KEYINPUT41), .B(n404), .Z(n539) );
  INV_X1 U458 ( .A(n539), .ZN(n569) );
  NAND2_X1 U459 ( .A1(n569), .A2(n578), .ZN(n405) );
  XNOR2_X1 U460 ( .A(KEYINPUT46), .B(n405), .ZN(n408) );
  NOR2_X1 U461 ( .A1(n562), .A2(n406), .ZN(n407) );
  XNOR2_X1 U462 ( .A(KEYINPUT47), .B(n409), .ZN(n410) );
  NAND2_X1 U463 ( .A1(n411), .A2(n410), .ZN(n412) );
  XNOR2_X1 U464 ( .A(n412), .B(KEYINPUT48), .ZN(n552) );
  XOR2_X1 U465 ( .A(n413), .B(KEYINPUT89), .Z(n415) );
  NAND2_X1 U466 ( .A1(G226GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U467 ( .A(n415), .B(n414), .ZN(n420) );
  XNOR2_X1 U468 ( .A(G218GAT), .B(G92GAT), .ZN(n418) );
  INV_X1 U469 ( .A(n416), .ZN(n417) );
  XNOR2_X1 U470 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U471 ( .A(n420), .B(n419), .Z(n424) );
  XNOR2_X1 U472 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U473 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U474 ( .A(n426), .B(n425), .ZN(n459) );
  NAND2_X1 U475 ( .A1(n552), .A2(n459), .ZN(n429) );
  XNOR2_X1 U476 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n427) );
  XNOR2_X1 U477 ( .A(n427), .B(KEYINPUT119), .ZN(n428) );
  XNOR2_X1 U478 ( .A(n429), .B(n428), .ZN(n450) );
  XOR2_X1 U479 ( .A(n430), .B(G134GAT), .Z(n432) );
  NAND2_X1 U480 ( .A1(G225GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U481 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U482 ( .A(G29GAT), .B(n433), .ZN(n449) );
  XOR2_X1 U483 ( .A(KEYINPUT88), .B(G57GAT), .Z(n435) );
  XNOR2_X1 U484 ( .A(G148GAT), .B(G155GAT), .ZN(n434) );
  XNOR2_X1 U485 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U486 ( .A(G85GAT), .B(G162GAT), .Z(n437) );
  XNOR2_X1 U487 ( .A(G120GAT), .B(G127GAT), .ZN(n436) );
  XNOR2_X1 U488 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U489 ( .A(n439), .B(n438), .ZN(n447) );
  XOR2_X1 U490 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n441) );
  XNOR2_X1 U491 ( .A(KEYINPUT5), .B(KEYINPUT1), .ZN(n440) );
  XNOR2_X1 U492 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U493 ( .A(KEYINPUT87), .B(n442), .Z(n445) );
  XNOR2_X1 U494 ( .A(G1GAT), .B(n443), .ZN(n444) );
  XNOR2_X1 U495 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U496 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U497 ( .A(n449), .B(n448), .ZN(n523) );
  NAND2_X1 U498 ( .A1(n450), .A2(n523), .ZN(n576) );
  NOR2_X1 U499 ( .A1(n466), .A2(n576), .ZN(n451) );
  XNOR2_X1 U500 ( .A(n451), .B(KEYINPUT55), .ZN(n452) );
  NOR2_X1 U501 ( .A1(n534), .A2(n452), .ZN(n453) );
  NAND2_X1 U502 ( .A1(n572), .A2(n547), .ZN(n455) );
  XNOR2_X1 U503 ( .A(n455), .B(n454), .ZN(G1351GAT) );
  XOR2_X1 U504 ( .A(KEYINPUT34), .B(KEYINPUT96), .Z(n457) );
  XNOR2_X1 U505 ( .A(G1GAT), .B(KEYINPUT95), .ZN(n456) );
  XNOR2_X1 U506 ( .A(n457), .B(n456), .ZN(n479) );
  NAND2_X1 U507 ( .A1(n404), .A2(n578), .ZN(n458) );
  XNOR2_X1 U508 ( .A(n458), .B(KEYINPUT69), .ZN(n493) );
  XOR2_X1 U509 ( .A(n466), .B(KEYINPUT28), .Z(n530) );
  INV_X1 U510 ( .A(n459), .ZN(n525) );
  XNOR2_X1 U511 ( .A(KEYINPUT27), .B(n525), .ZN(n468) );
  NOR2_X1 U512 ( .A1(n468), .A2(n523), .ZN(n460) );
  XNOR2_X1 U513 ( .A(n460), .B(KEYINPUT90), .ZN(n551) );
  NAND2_X1 U514 ( .A1(n530), .A2(n551), .ZN(n533) );
  XNOR2_X1 U515 ( .A(KEYINPUT91), .B(n533), .ZN(n462) );
  XOR2_X1 U516 ( .A(n534), .B(KEYINPUT83), .Z(n461) );
  NAND2_X1 U517 ( .A1(n462), .A2(n461), .ZN(n463) );
  XNOR2_X1 U518 ( .A(n463), .B(KEYINPUT92), .ZN(n473) );
  NOR2_X1 U519 ( .A1(n534), .A2(n525), .ZN(n464) );
  NOR2_X1 U520 ( .A1(n466), .A2(n464), .ZN(n465) );
  XNOR2_X1 U521 ( .A(n465), .B(KEYINPUT25), .ZN(n470) );
  NAND2_X1 U522 ( .A1(n466), .A2(n534), .ZN(n467) );
  XNOR2_X1 U523 ( .A(KEYINPUT26), .B(n467), .ZN(n577) );
  OR2_X1 U524 ( .A1(n468), .A2(n577), .ZN(n469) );
  NAND2_X1 U525 ( .A1(n470), .A2(n469), .ZN(n471) );
  NAND2_X1 U526 ( .A1(n523), .A2(n471), .ZN(n472) );
  NAND2_X1 U527 ( .A1(n473), .A2(n472), .ZN(n488) );
  NOR2_X1 U528 ( .A1(n542), .A2(n547), .ZN(n475) );
  XNOR2_X1 U529 ( .A(KEYINPUT16), .B(KEYINPUT78), .ZN(n474) );
  XNOR2_X1 U530 ( .A(n475), .B(n474), .ZN(n476) );
  NAND2_X1 U531 ( .A1(n488), .A2(n476), .ZN(n477) );
  XNOR2_X1 U532 ( .A(n477), .B(KEYINPUT93), .ZN(n508) );
  NAND2_X1 U533 ( .A1(n493), .A2(n508), .ZN(n486) );
  NOR2_X1 U534 ( .A1(n523), .A2(n486), .ZN(n478) );
  XOR2_X1 U535 ( .A(n479), .B(n478), .Z(n480) );
  XNOR2_X1 U536 ( .A(KEYINPUT94), .B(n480), .ZN(G1324GAT) );
  NOR2_X1 U537 ( .A1(n525), .A2(n486), .ZN(n481) );
  XOR2_X1 U538 ( .A(G8GAT), .B(n481), .Z(G1325GAT) );
  NOR2_X1 U539 ( .A1(n486), .A2(n534), .ZN(n485) );
  XOR2_X1 U540 ( .A(KEYINPUT97), .B(KEYINPUT35), .Z(n483) );
  XNOR2_X1 U541 ( .A(G15GAT), .B(KEYINPUT98), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(G1326GAT) );
  NOR2_X1 U544 ( .A1(n530), .A2(n486), .ZN(n487) );
  XOR2_X1 U545 ( .A(G22GAT), .B(n487), .Z(G1327GAT) );
  NAND2_X1 U546 ( .A1(n542), .A2(n488), .ZN(n489) );
  XNOR2_X1 U547 ( .A(KEYINPUT99), .B(n489), .ZN(n490) );
  NAND2_X1 U548 ( .A1(n490), .A2(n586), .ZN(n492) );
  XNOR2_X1 U549 ( .A(KEYINPUT100), .B(KEYINPUT37), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n492), .B(n491), .ZN(n521) );
  NAND2_X1 U551 ( .A1(n521), .A2(n493), .ZN(n494) );
  XNOR2_X1 U552 ( .A(n494), .B(KEYINPUT38), .ZN(n504) );
  NOR2_X1 U553 ( .A1(n523), .A2(n504), .ZN(n497) );
  XOR2_X1 U554 ( .A(G29GAT), .B(KEYINPUT39), .Z(n495) );
  XNOR2_X1 U555 ( .A(KEYINPUT101), .B(n495), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n497), .B(n496), .ZN(G1328GAT) );
  NOR2_X1 U557 ( .A1(n525), .A2(n504), .ZN(n498) );
  XOR2_X1 U558 ( .A(KEYINPUT102), .B(n498), .Z(n499) );
  XNOR2_X1 U559 ( .A(G36GAT), .B(n499), .ZN(G1329GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n501) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(KEYINPUT104), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n501), .B(n500), .ZN(n503) );
  NOR2_X1 U563 ( .A1(n534), .A2(n504), .ZN(n502) );
  XOR2_X1 U564 ( .A(n503), .B(n502), .Z(G1330GAT) );
  XNOR2_X1 U565 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n506) );
  NOR2_X1 U566 ( .A1(n530), .A2(n504), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U568 ( .A(G50GAT), .B(n507), .ZN(G1331GAT) );
  NOR2_X1 U569 ( .A1(n578), .A2(n539), .ZN(n522) );
  NAND2_X1 U570 ( .A1(n522), .A2(n508), .ZN(n518) );
  NOR2_X1 U571 ( .A1(n523), .A2(n518), .ZN(n510) );
  XNOR2_X1 U572 ( .A(KEYINPUT107), .B(KEYINPUT42), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U574 ( .A(G57GAT), .B(n511), .ZN(G1332GAT) );
  NOR2_X1 U575 ( .A1(n525), .A2(n518), .ZN(n513) );
  XNOR2_X1 U576 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U578 ( .A(G64GAT), .B(n514), .ZN(G1333GAT) );
  NOR2_X1 U579 ( .A1(n534), .A2(n518), .ZN(n516) );
  XNOR2_X1 U580 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U582 ( .A(G71GAT), .B(n517), .ZN(G1334GAT) );
  NOR2_X1 U583 ( .A1(n530), .A2(n518), .ZN(n520) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  NAND2_X1 U586 ( .A1(n522), .A2(n521), .ZN(n529) );
  NOR2_X1 U587 ( .A1(n523), .A2(n529), .ZN(n524) );
  XOR2_X1 U588 ( .A(G85GAT), .B(n524), .Z(G1336GAT) );
  NOR2_X1 U589 ( .A1(n525), .A2(n529), .ZN(n526) );
  XOR2_X1 U590 ( .A(G92GAT), .B(n526), .Z(G1337GAT) );
  NOR2_X1 U591 ( .A1(n534), .A2(n529), .ZN(n527) );
  XOR2_X1 U592 ( .A(KEYINPUT112), .B(n527), .Z(n528) );
  XNOR2_X1 U593 ( .A(G99GAT), .B(n528), .ZN(G1338GAT) );
  NOR2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U595 ( .A(KEYINPUT44), .B(n531), .Z(n532) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n532), .ZN(G1339GAT) );
  NOR2_X1 U597 ( .A1(n534), .A2(n533), .ZN(n535) );
  NAND2_X1 U598 ( .A1(n552), .A2(n535), .ZN(n546) );
  NOR2_X1 U599 ( .A1(n536), .A2(n546), .ZN(n537) );
  XOR2_X1 U600 ( .A(KEYINPUT114), .B(n537), .Z(n538) );
  XNOR2_X1 U601 ( .A(G113GAT), .B(n538), .ZN(G1340GAT) );
  NOR2_X1 U602 ( .A1(n539), .A2(n546), .ZN(n541) );
  XNOR2_X1 U603 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n540) );
  XNOR2_X1 U604 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  NOR2_X1 U605 ( .A1(n542), .A2(n546), .ZN(n544) );
  XNOR2_X1 U606 ( .A(KEYINPUT50), .B(KEYINPUT115), .ZN(n543) );
  XNOR2_X1 U607 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(n545), .ZN(G1342GAT) );
  XOR2_X1 U609 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  INV_X1 U610 ( .A(n546), .ZN(n548) );
  NAND2_X1 U611 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U612 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  NAND2_X1 U613 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U614 ( .A1(n577), .A2(n553), .ZN(n561) );
  NAND2_X1 U615 ( .A1(n578), .A2(n561), .ZN(n554) );
  XNOR2_X1 U616 ( .A(n554), .B(KEYINPUT116), .ZN(n555) );
  XNOR2_X1 U617 ( .A(G141GAT), .B(n555), .ZN(G1344GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n557) );
  NAND2_X1 U619 ( .A1(n561), .A2(n569), .ZN(n556) );
  XNOR2_X1 U620 ( .A(n557), .B(n556), .ZN(n559) );
  XOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT53), .Z(n558) );
  XNOR2_X1 U622 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U623 ( .A1(n406), .A2(n561), .ZN(n560) );
  XNOR2_X1 U624 ( .A(n560), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U625 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U626 ( .A(n563), .B(KEYINPUT118), .ZN(n564) );
  XNOR2_X1 U627 ( .A(G162GAT), .B(n564), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n578), .A2(n572), .ZN(n565) );
  XNOR2_X1 U629 ( .A(n565), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n567) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  XOR2_X1 U633 ( .A(KEYINPUT56), .B(n568), .Z(n571) );
  NAND2_X1 U634 ( .A1(n572), .A2(n569), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n571), .B(n570), .ZN(G1349GAT) );
  NAND2_X1 U636 ( .A1(n406), .A2(n572), .ZN(n573) );
  XNOR2_X1 U637 ( .A(n573), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(KEYINPUT60), .ZN(n575) );
  XOR2_X1 U640 ( .A(KEYINPUT59), .B(n575), .Z(n580) );
  NOR2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n587) );
  NAND2_X1 U642 ( .A1(n587), .A2(n578), .ZN(n579) );
  XNOR2_X1 U643 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .Z(n583) );
  INV_X1 U645 ( .A(n404), .ZN(n581) );
  NAND2_X1 U646 ( .A1(n587), .A2(n581), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  XOR2_X1 U648 ( .A(G211GAT), .B(KEYINPUT125), .Z(n585) );
  NAND2_X1 U649 ( .A1(n587), .A2(n406), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1354GAT) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n591) );
  XOR2_X1 U652 ( .A(KEYINPUT127), .B(KEYINPUT126), .Z(n589) );
  NAND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(G1355GAT) );
endmodule

