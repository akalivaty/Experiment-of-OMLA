

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581;

  XOR2_X1 U324 ( .A(KEYINPUT2), .B(G162GAT), .Z(n293) );
  XNOR2_X1 U325 ( .A(G155GAT), .B(G148GAT), .ZN(n292) );
  XNOR2_X1 U326 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U327 ( .A(KEYINPUT3), .B(n294), .Z(n381) );
  XOR2_X1 U328 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n296) );
  XNOR2_X1 U329 ( .A(KEYINPUT93), .B(KEYINPUT5), .ZN(n295) );
  XNOR2_X1 U330 ( .A(n296), .B(n295), .ZN(n303) );
  XOR2_X1 U331 ( .A(KEYINPUT94), .B(KEYINPUT4), .Z(n298) );
  XNOR2_X1 U332 ( .A(KEYINPUT1), .B(KEYINPUT92), .ZN(n297) );
  XNOR2_X1 U333 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U334 ( .A(n299), .B(KEYINPUT84), .Z(n301) );
  XOR2_X1 U335 ( .A(G85GAT), .B(G57GAT), .Z(n316) );
  XNOR2_X1 U336 ( .A(G29GAT), .B(n316), .ZN(n300) );
  XNOR2_X1 U337 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U338 ( .A(n303), .B(n302), .Z(n312) );
  XOR2_X1 U339 ( .A(KEYINPUT86), .B(G134GAT), .Z(n305) );
  XNOR2_X1 U340 ( .A(G127GAT), .B(G120GAT), .ZN(n304) );
  XNOR2_X1 U341 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U342 ( .A(KEYINPUT0), .B(n306), .Z(n394) );
  XNOR2_X1 U343 ( .A(G113GAT), .B(G141GAT), .ZN(n307) );
  XNOR2_X1 U344 ( .A(n307), .B(G1GAT), .ZN(n339) );
  XOR2_X1 U345 ( .A(KEYINPUT6), .B(n339), .Z(n309) );
  NAND2_X1 U346 ( .A1(G225GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U347 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U348 ( .A(n394), .B(n310), .ZN(n311) );
  XNOR2_X1 U349 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U350 ( .A(n381), .B(n313), .ZN(n405) );
  XNOR2_X1 U351 ( .A(KEYINPUT97), .B(n405), .ZN(n544) );
  XOR2_X1 U352 ( .A(KEYINPUT13), .B(KEYINPUT77), .Z(n315) );
  XNOR2_X1 U353 ( .A(G148GAT), .B(G92GAT), .ZN(n314) );
  XNOR2_X1 U354 ( .A(n315), .B(n314), .ZN(n317) );
  XOR2_X1 U355 ( .A(n317), .B(n316), .Z(n319) );
  XNOR2_X1 U356 ( .A(G120GAT), .B(G176GAT), .ZN(n318) );
  XNOR2_X1 U357 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U358 ( .A(KEYINPUT79), .B(G64GAT), .Z(n361) );
  XOR2_X1 U359 ( .A(n320), .B(n361), .Z(n324) );
  XOR2_X1 U360 ( .A(G99GAT), .B(G71GAT), .Z(n383) );
  XOR2_X1 U361 ( .A(G78GAT), .B(G204GAT), .Z(n322) );
  XNOR2_X1 U362 ( .A(G106GAT), .B(KEYINPUT76), .ZN(n321) );
  XNOR2_X1 U363 ( .A(n322), .B(n321), .ZN(n372) );
  XNOR2_X1 U364 ( .A(n383), .B(n372), .ZN(n323) );
  XNOR2_X1 U365 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U366 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n326) );
  NAND2_X1 U367 ( .A1(G230GAT), .A2(G233GAT), .ZN(n325) );
  XNOR2_X1 U368 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U369 ( .A(n328), .B(n327), .Z(n333) );
  XOR2_X1 U370 ( .A(KEYINPUT78), .B(KEYINPUT32), .Z(n330) );
  XNOR2_X1 U371 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n329) );
  XNOR2_X1 U372 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U373 ( .A(n331), .B(KEYINPUT75), .ZN(n332) );
  XNOR2_X1 U374 ( .A(n333), .B(n332), .ZN(n569) );
  XOR2_X1 U375 ( .A(KEYINPUT73), .B(KEYINPUT70), .Z(n335) );
  XNOR2_X1 U376 ( .A(KEYINPUT67), .B(KEYINPUT29), .ZN(n334) );
  XNOR2_X1 U377 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U378 ( .A(n336), .B(G197GAT), .Z(n338) );
  XOR2_X1 U379 ( .A(G22GAT), .B(G8GAT), .Z(n443) );
  XNOR2_X1 U380 ( .A(n443), .B(G43GAT), .ZN(n337) );
  XNOR2_X1 U381 ( .A(n338), .B(n337), .ZN(n343) );
  XOR2_X1 U382 ( .A(G169GAT), .B(G15GAT), .Z(n390) );
  XOR2_X1 U383 ( .A(n390), .B(n339), .Z(n341) );
  NAND2_X1 U384 ( .A1(G229GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U385 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U386 ( .A(n343), .B(n342), .Z(n352) );
  XNOR2_X1 U387 ( .A(G36GAT), .B(KEYINPUT72), .ZN(n344) );
  XNOR2_X1 U388 ( .A(n344), .B(G29GAT), .ZN(n345) );
  XOR2_X1 U389 ( .A(n345), .B(KEYINPUT7), .Z(n347) );
  XNOR2_X1 U390 ( .A(G50GAT), .B(KEYINPUT8), .ZN(n346) );
  XNOR2_X1 U391 ( .A(n347), .B(n346), .ZN(n410) );
  XOR2_X1 U392 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n349) );
  XNOR2_X1 U393 ( .A(KEYINPUT71), .B(KEYINPUT30), .ZN(n348) );
  XNOR2_X1 U394 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U395 ( .A(n410), .B(n350), .ZN(n351) );
  XNOR2_X1 U396 ( .A(n352), .B(n351), .ZN(n564) );
  XOR2_X1 U397 ( .A(n564), .B(KEYINPUT74), .Z(n550) );
  INV_X1 U398 ( .A(n550), .ZN(n511) );
  NOR2_X1 U399 ( .A1(n569), .A2(n511), .ZN(n463) );
  XOR2_X1 U400 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n354) );
  XNOR2_X1 U401 ( .A(G183GAT), .B(G176GAT), .ZN(n353) );
  XNOR2_X1 U402 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U403 ( .A(KEYINPUT18), .B(n355), .Z(n395) );
  XOR2_X1 U404 ( .A(KEYINPUT90), .B(G218GAT), .Z(n357) );
  XNOR2_X1 U405 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n356) );
  XNOR2_X1 U406 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U407 ( .A(G197GAT), .B(n358), .Z(n380) );
  XNOR2_X1 U408 ( .A(n395), .B(n380), .ZN(n369) );
  XOR2_X1 U409 ( .A(KEYINPUT98), .B(G204GAT), .Z(n360) );
  XNOR2_X1 U410 ( .A(G169GAT), .B(G8GAT), .ZN(n359) );
  XNOR2_X1 U411 ( .A(n360), .B(n359), .ZN(n365) );
  XOR2_X1 U412 ( .A(KEYINPUT85), .B(G92GAT), .Z(n426) );
  XOR2_X1 U413 ( .A(n361), .B(n426), .Z(n363) );
  XNOR2_X1 U414 ( .A(G36GAT), .B(G190GAT), .ZN(n362) );
  XNOR2_X1 U415 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U416 ( .A(n365), .B(n364), .Z(n367) );
  NAND2_X1 U417 ( .A1(G226GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U418 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U419 ( .A(n369), .B(n368), .ZN(n542) );
  XNOR2_X1 U420 ( .A(n542), .B(KEYINPUT27), .ZN(n402) );
  NOR2_X1 U421 ( .A1(n544), .A2(n402), .ZN(n526) );
  XOR2_X1 U422 ( .A(KEYINPUT91), .B(KEYINPUT23), .Z(n371) );
  XNOR2_X1 U423 ( .A(G50GAT), .B(KEYINPUT22), .ZN(n370) );
  XNOR2_X1 U424 ( .A(n371), .B(n370), .ZN(n373) );
  XOR2_X1 U425 ( .A(n373), .B(n372), .Z(n378) );
  XOR2_X1 U426 ( .A(G22GAT), .B(KEYINPUT24), .Z(n375) );
  NAND2_X1 U427 ( .A1(G228GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U428 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U429 ( .A(G141GAT), .B(n376), .ZN(n377) );
  XNOR2_X1 U430 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U431 ( .A(n380), .B(n379), .ZN(n382) );
  XOR2_X1 U432 ( .A(n382), .B(n381), .Z(n546) );
  XOR2_X1 U433 ( .A(KEYINPUT28), .B(n546), .Z(n494) );
  NAND2_X1 U434 ( .A1(n526), .A2(n494), .ZN(n508) );
  XOR2_X1 U435 ( .A(KEYINPUT88), .B(n383), .Z(n385) );
  XOR2_X1 U436 ( .A(G43GAT), .B(G190GAT), .Z(n427) );
  XNOR2_X1 U437 ( .A(G113GAT), .B(n427), .ZN(n384) );
  XNOR2_X1 U438 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U439 ( .A(KEYINPUT64), .B(KEYINPUT87), .Z(n387) );
  NAND2_X1 U440 ( .A1(G227GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U441 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U442 ( .A(n389), .B(n388), .Z(n392) );
  XNOR2_X1 U443 ( .A(n390), .B(KEYINPUT20), .ZN(n391) );
  XNOR2_X1 U444 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U445 ( .A(n394), .B(n393), .ZN(n396) );
  XNOR2_X1 U446 ( .A(n396), .B(n395), .ZN(n510) );
  INV_X1 U447 ( .A(n510), .ZN(n549) );
  XNOR2_X1 U448 ( .A(KEYINPUT89), .B(n549), .ZN(n397) );
  NOR2_X1 U449 ( .A1(n508), .A2(n397), .ZN(n409) );
  NOR2_X1 U450 ( .A1(n542), .A2(n549), .ZN(n398) );
  XOR2_X1 U451 ( .A(KEYINPUT99), .B(n398), .Z(n399) );
  NOR2_X1 U452 ( .A1(n546), .A2(n399), .ZN(n400) );
  XOR2_X1 U453 ( .A(KEYINPUT25), .B(n400), .Z(n404) );
  NAND2_X1 U454 ( .A1(n546), .A2(n549), .ZN(n401) );
  XNOR2_X1 U455 ( .A(n401), .B(KEYINPUT26), .ZN(n563) );
  NOR2_X1 U456 ( .A1(n563), .A2(n402), .ZN(n403) );
  NOR2_X1 U457 ( .A1(n404), .A2(n403), .ZN(n406) );
  NOR2_X1 U458 ( .A1(n406), .A2(n405), .ZN(n407) );
  XNOR2_X1 U459 ( .A(n407), .B(KEYINPUT100), .ZN(n408) );
  NOR2_X1 U460 ( .A1(n409), .A2(n408), .ZN(n459) );
  INV_X1 U461 ( .A(n410), .ZN(n431) );
  XOR2_X1 U462 ( .A(KEYINPUT9), .B(KEYINPUT66), .Z(n412) );
  XNOR2_X1 U463 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(n411) );
  XNOR2_X1 U464 ( .A(n412), .B(n411), .ZN(n416) );
  XOR2_X1 U465 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n414) );
  XNOR2_X1 U466 ( .A(KEYINPUT84), .B(KEYINPUT77), .ZN(n413) );
  XNOR2_X1 U467 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U468 ( .A(n416), .B(n415), .Z(n421) );
  XOR2_X1 U469 ( .A(G85GAT), .B(G162GAT), .Z(n418) );
  NAND2_X1 U470 ( .A1(G232GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U471 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U472 ( .A(G134GAT), .B(n419), .ZN(n420) );
  XNOR2_X1 U473 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U474 ( .A(KEYINPUT65), .B(G106GAT), .Z(n423) );
  XNOR2_X1 U475 ( .A(G99GAT), .B(G218GAT), .ZN(n422) );
  XNOR2_X1 U476 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U477 ( .A(n425), .B(n424), .Z(n429) );
  XNOR2_X1 U478 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U479 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U480 ( .A(n431), .B(n430), .Z(n538) );
  INV_X1 U481 ( .A(n538), .ZN(n557) );
  XOR2_X1 U482 ( .A(G71GAT), .B(G183GAT), .Z(n433) );
  XNOR2_X1 U483 ( .A(G15GAT), .B(G127GAT), .ZN(n432) );
  XNOR2_X1 U484 ( .A(n433), .B(n432), .ZN(n447) );
  XOR2_X1 U485 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n435) );
  NAND2_X1 U486 ( .A1(G231GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U487 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U488 ( .A(KEYINPUT15), .B(KEYINPUT13), .Z(n437) );
  XNOR2_X1 U489 ( .A(G1GAT), .B(G57GAT), .ZN(n436) );
  XNOR2_X1 U490 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U491 ( .A(n439), .B(n438), .Z(n445) );
  XOR2_X1 U492 ( .A(G64GAT), .B(G78GAT), .Z(n441) );
  XNOR2_X1 U493 ( .A(G211GAT), .B(G155GAT), .ZN(n440) );
  XNOR2_X1 U494 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U495 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U496 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U497 ( .A(n447), .B(n446), .Z(n572) );
  INV_X1 U498 ( .A(n572), .ZN(n535) );
  NOR2_X1 U499 ( .A1(n557), .A2(n535), .ZN(n448) );
  XOR2_X1 U500 ( .A(KEYINPUT16), .B(n448), .Z(n449) );
  NOR2_X1 U501 ( .A1(n459), .A2(n449), .ZN(n450) );
  XOR2_X1 U502 ( .A(KEYINPUT101), .B(n450), .Z(n475) );
  NAND2_X1 U503 ( .A1(n463), .A2(n475), .ZN(n457) );
  NOR2_X1 U504 ( .A1(n544), .A2(n457), .ZN(n451) );
  XOR2_X1 U505 ( .A(G1GAT), .B(n451), .Z(n452) );
  XNOR2_X1 U506 ( .A(KEYINPUT34), .B(n452), .ZN(G1324GAT) );
  NOR2_X1 U507 ( .A1(n542), .A2(n457), .ZN(n453) );
  XOR2_X1 U508 ( .A(KEYINPUT102), .B(n453), .Z(n454) );
  XNOR2_X1 U509 ( .A(G8GAT), .B(n454), .ZN(G1325GAT) );
  NOR2_X1 U510 ( .A1(n549), .A2(n457), .ZN(n456) );
  XNOR2_X1 U511 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n455) );
  XNOR2_X1 U512 ( .A(n456), .B(n455), .ZN(G1326GAT) );
  NOR2_X1 U513 ( .A1(n494), .A2(n457), .ZN(n458) );
  XOR2_X1 U514 ( .A(G22GAT), .B(n458), .Z(G1327GAT) );
  XNOR2_X1 U515 ( .A(KEYINPUT39), .B(KEYINPUT104), .ZN(n466) );
  XOR2_X1 U516 ( .A(KEYINPUT37), .B(KEYINPUT103), .Z(n462) );
  XNOR2_X1 U517 ( .A(KEYINPUT36), .B(n538), .ZN(n579) );
  NOR2_X1 U518 ( .A1(n579), .A2(n459), .ZN(n460) );
  NAND2_X1 U519 ( .A1(n460), .A2(n535), .ZN(n461) );
  XNOR2_X1 U520 ( .A(n462), .B(n461), .ZN(n486) );
  NAND2_X1 U521 ( .A1(n486), .A2(n463), .ZN(n464) );
  XNOR2_X1 U522 ( .A(KEYINPUT38), .B(n464), .ZN(n473) );
  NOR2_X1 U523 ( .A1(n544), .A2(n473), .ZN(n465) );
  XNOR2_X1 U524 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U525 ( .A(G29GAT), .B(n467), .ZN(G1328GAT) );
  XNOR2_X1 U526 ( .A(G36GAT), .B(KEYINPUT105), .ZN(n469) );
  NOR2_X1 U527 ( .A1(n542), .A2(n473), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n469), .B(n468), .ZN(G1329GAT) );
  NOR2_X1 U529 ( .A1(n473), .A2(n549), .ZN(n471) );
  XNOR2_X1 U530 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n470) );
  XNOR2_X1 U531 ( .A(n471), .B(n470), .ZN(n472) );
  XOR2_X1 U532 ( .A(G43GAT), .B(n472), .Z(G1330GAT) );
  NOR2_X1 U533 ( .A1(n473), .A2(n494), .ZN(n474) );
  XOR2_X1 U534 ( .A(G50GAT), .B(n474), .Z(G1331GAT) );
  XNOR2_X1 U535 ( .A(n569), .B(KEYINPUT41), .ZN(n529) );
  INV_X1 U536 ( .A(n529), .ZN(n552) );
  AND2_X1 U537 ( .A1(n564), .A2(n552), .ZN(n485) );
  NAND2_X1 U538 ( .A1(n475), .A2(n485), .ZN(n480) );
  NOR2_X1 U539 ( .A1(n544), .A2(n480), .ZN(n476) );
  XOR2_X1 U540 ( .A(G57GAT), .B(n476), .Z(n477) );
  XNOR2_X1 U541 ( .A(KEYINPUT42), .B(n477), .ZN(G1332GAT) );
  NOR2_X1 U542 ( .A1(n542), .A2(n480), .ZN(n478) );
  XOR2_X1 U543 ( .A(G64GAT), .B(n478), .Z(G1333GAT) );
  NOR2_X1 U544 ( .A1(n549), .A2(n480), .ZN(n479) );
  XOR2_X1 U545 ( .A(G71GAT), .B(n479), .Z(G1334GAT) );
  NOR2_X1 U546 ( .A1(n480), .A2(n494), .ZN(n484) );
  XOR2_X1 U547 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n482) );
  XNOR2_X1 U548 ( .A(G78GAT), .B(KEYINPUT108), .ZN(n481) );
  XNOR2_X1 U549 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U550 ( .A(n484), .B(n483), .ZN(G1335GAT) );
  NAND2_X1 U551 ( .A1(n486), .A2(n485), .ZN(n493) );
  NOR2_X1 U552 ( .A1(n544), .A2(n493), .ZN(n488) );
  XNOR2_X1 U553 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n487) );
  XNOR2_X1 U554 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U555 ( .A(G85GAT), .B(n489), .ZN(G1336GAT) );
  NOR2_X1 U556 ( .A1(n542), .A2(n493), .ZN(n491) );
  XNOR2_X1 U557 ( .A(G92GAT), .B(KEYINPUT111), .ZN(n490) );
  XNOR2_X1 U558 ( .A(n491), .B(n490), .ZN(G1337GAT) );
  NOR2_X1 U559 ( .A1(n549), .A2(n493), .ZN(n492) );
  XOR2_X1 U560 ( .A(G99GAT), .B(n492), .Z(G1338GAT) );
  NOR2_X1 U561 ( .A1(n494), .A2(n493), .ZN(n495) );
  XOR2_X1 U562 ( .A(KEYINPUT44), .B(n495), .Z(n496) );
  XNOR2_X1 U563 ( .A(G106GAT), .B(n496), .ZN(G1339GAT) );
  NOR2_X1 U564 ( .A1(n557), .A2(n572), .ZN(n500) );
  NOR2_X1 U565 ( .A1(n564), .A2(n529), .ZN(n498) );
  XOR2_X1 U566 ( .A(KEYINPUT112), .B(KEYINPUT46), .Z(n497) );
  XNOR2_X1 U567 ( .A(n498), .B(n497), .ZN(n499) );
  NAND2_X1 U568 ( .A1(n500), .A2(n499), .ZN(n501) );
  XNOR2_X1 U569 ( .A(n501), .B(KEYINPUT47), .ZN(n506) );
  NOR2_X1 U570 ( .A1(n579), .A2(n535), .ZN(n502) );
  XNOR2_X1 U571 ( .A(n502), .B(KEYINPUT45), .ZN(n503) );
  NAND2_X1 U572 ( .A1(n503), .A2(n511), .ZN(n504) );
  NOR2_X1 U573 ( .A1(n504), .A2(n569), .ZN(n505) );
  NOR2_X1 U574 ( .A1(n506), .A2(n505), .ZN(n507) );
  XNOR2_X1 U575 ( .A(KEYINPUT48), .B(n507), .ZN(n541) );
  NOR2_X1 U576 ( .A1(n541), .A2(n508), .ZN(n509) );
  NAND2_X1 U577 ( .A1(n510), .A2(n509), .ZN(n521) );
  NOR2_X1 U578 ( .A1(n511), .A2(n521), .ZN(n513) );
  XNOR2_X1 U579 ( .A(G113GAT), .B(KEYINPUT113), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n513), .B(n512), .ZN(G1340GAT) );
  NOR2_X1 U581 ( .A1(n521), .A2(n529), .ZN(n517) );
  XOR2_X1 U582 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n515) );
  XNOR2_X1 U583 ( .A(G120GAT), .B(KEYINPUT114), .ZN(n514) );
  XNOR2_X1 U584 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n517), .B(n516), .ZN(G1341GAT) );
  NOR2_X1 U586 ( .A1(n535), .A2(n521), .ZN(n519) );
  XNOR2_X1 U587 ( .A(KEYINPUT116), .B(KEYINPUT50), .ZN(n518) );
  XNOR2_X1 U588 ( .A(n519), .B(n518), .ZN(n520) );
  XOR2_X1 U589 ( .A(G127GAT), .B(n520), .Z(G1342GAT) );
  NOR2_X1 U590 ( .A1(n538), .A2(n521), .ZN(n523) );
  XNOR2_X1 U591 ( .A(KEYINPUT51), .B(KEYINPUT117), .ZN(n522) );
  XNOR2_X1 U592 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U593 ( .A(G134GAT), .B(n524), .Z(G1343GAT) );
  NOR2_X1 U594 ( .A1(n563), .A2(n541), .ZN(n525) );
  NAND2_X1 U595 ( .A1(n526), .A2(n525), .ZN(n537) );
  NOR2_X1 U596 ( .A1(n564), .A2(n537), .ZN(n527) );
  XOR2_X1 U597 ( .A(KEYINPUT118), .B(n527), .Z(n528) );
  XNOR2_X1 U598 ( .A(G141GAT), .B(n528), .ZN(G1344GAT) );
  NOR2_X1 U599 ( .A1(n529), .A2(n537), .ZN(n534) );
  XOR2_X1 U600 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n531) );
  XNOR2_X1 U601 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n530) );
  XNOR2_X1 U602 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U603 ( .A(KEYINPUT119), .B(n532), .ZN(n533) );
  XNOR2_X1 U604 ( .A(n534), .B(n533), .ZN(G1345GAT) );
  NOR2_X1 U605 ( .A1(n535), .A2(n537), .ZN(n536) );
  XOR2_X1 U606 ( .A(G155GAT), .B(n536), .Z(G1346GAT) );
  NOR2_X1 U607 ( .A1(n538), .A2(n537), .ZN(n540) );
  XNOR2_X1 U608 ( .A(G162GAT), .B(KEYINPUT121), .ZN(n539) );
  XNOR2_X1 U609 ( .A(n540), .B(n539), .ZN(G1347GAT) );
  NOR2_X1 U610 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U611 ( .A(KEYINPUT54), .B(n543), .ZN(n545) );
  NAND2_X1 U612 ( .A1(n545), .A2(n544), .ZN(n562) );
  NOR2_X1 U613 ( .A1(n546), .A2(n562), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n547), .B(KEYINPUT55), .ZN(n548) );
  NOR2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n558) );
  NAND2_X1 U616 ( .A1(n558), .A2(n550), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n551), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n554) );
  NAND2_X1 U619 ( .A1(n558), .A2(n552), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U621 ( .A(G176GAT), .B(n555), .ZN(G1349GAT) );
  NAND2_X1 U622 ( .A1(n558), .A2(n572), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT58), .B(KEYINPUT122), .Z(n560) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U627 ( .A(G190GAT), .B(n561), .Z(G1351GAT) );
  NOR2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n573) );
  INV_X1 U629 ( .A(n573), .ZN(n578) );
  NOR2_X1 U630 ( .A1(n578), .A2(n564), .ZN(n568) );
  XOR2_X1 U631 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n566) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .Z(n571) );
  NAND2_X1 U636 ( .A1(n573), .A2(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1353GAT) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(KEYINPUT124), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G211GAT), .B(n575), .ZN(G1354GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n577) );
  XNOR2_X1 U642 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n581) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U645 ( .A(n581), .B(n580), .Z(G1355GAT) );
endmodule

