//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 0 0 1 0 1 1 1 1 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n830, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950;
  XOR2_X1   g000(.A(G57gat), .B(G85gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G1gat), .B(G29gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G225gat), .A2(G233gat), .ZN(new_n207));
  XOR2_X1   g006(.A(G141gat), .B(G148gat), .Z(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT77), .ZN(new_n209));
  INV_X1    g008(.A(G155gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT78), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT78), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G155gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n213), .A3(G162gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT2), .ZN(new_n215));
  XNOR2_X1  g014(.A(G155gat), .B(G162gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(G141gat), .B(G148gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT77), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n209), .A2(new_n215), .A3(new_n216), .A4(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n216), .B1(new_n208), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(G127gat), .B(G134gat), .Z(new_n225));
  XNOR2_X1  g024(.A(G113gat), .B(G120gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n226), .ZN(new_n227));
  XOR2_X1   g026(.A(G113gat), .B(G120gat), .Z(new_n228));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n229));
  XNOR2_X1  g028(.A(G127gat), .B(G134gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n224), .A2(new_n232), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n227), .A2(new_n231), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(new_n223), .A3(new_n220), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n207), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NOR3_X1   g036(.A1(new_n224), .A2(new_n232), .A3(KEYINPUT4), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT4), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n217), .B(KEYINPUT77), .ZN(new_n240));
  XOR2_X1   g039(.A(G155gat), .B(G162gat), .Z(new_n241));
  AOI21_X1  g040(.A(new_n241), .B1(KEYINPUT2), .B2(new_n214), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n222), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n239), .B1(new_n243), .B2(new_n234), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n232), .B1(new_n224), .B2(KEYINPUT3), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  OAI22_X1  g046(.A1(new_n238), .A2(new_n244), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n207), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n237), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(KEYINPUT5), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n235), .A2(KEYINPUT4), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n243), .A2(new_n239), .A3(new_n234), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n234), .B1(new_n243), .B2(new_n246), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n224), .A2(KEYINPUT3), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n254), .A2(new_n257), .A3(new_n207), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT5), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT85), .B1(new_n251), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n259), .B1(new_n258), .B2(new_n237), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n252), .A2(new_n253), .B1(new_n255), .B2(new_n256), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT5), .B1(new_n263), .B2(new_n207), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT85), .ZN(new_n265));
  NOR3_X1   g064(.A1(new_n262), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n206), .B1(new_n261), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT86), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n260), .ZN(new_n269));
  INV_X1    g068(.A(new_n206), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT6), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n267), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n269), .A2(new_n270), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT6), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n265), .B1(new_n262), .B2(new_n264), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n236), .B1(new_n263), .B2(new_n207), .ZN(new_n276));
  OAI211_X1 g075(.A(KEYINPUT85), .B(new_n260), .C1(new_n276), .C2(new_n259), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n270), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n262), .A2(new_n264), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n279), .B1(new_n280), .B2(new_n206), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT86), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  AND3_X1   g081(.A1(new_n272), .A2(new_n274), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G226gat), .A2(G233gat), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT69), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n286), .A2(G190gat), .ZN(new_n287));
  INV_X1    g086(.A(G190gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n288), .A2(KEYINPUT69), .ZN(new_n289));
  OR2_X1    g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT27), .B(G183gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT71), .B(KEYINPUT28), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G183gat), .A2(G190gat), .ZN(new_n295));
  INV_X1    g094(.A(G169gat), .ZN(new_n296));
  INV_X1    g095(.A(G176gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(new_n298), .B(KEYINPUT26), .Z(new_n299));
  AOI21_X1  g098(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n300));
  AND3_X1   g099(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n294), .A2(new_n295), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT24), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n295), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(G183gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(new_n288), .ZN(new_n307));
  NAND3_X1  g106(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT65), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n300), .ZN(new_n312));
  NAND3_X1  g111(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT23), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n312), .A2(new_n313), .B1(new_n298), .B2(new_n314), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n296), .A2(KEYINPUT66), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n296), .A2(KEYINPUT66), .ZN(new_n317));
  OAI211_X1 g116(.A(KEYINPUT23), .B(new_n297), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n305), .A2(new_n307), .A3(KEYINPUT65), .A4(new_n308), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n311), .A2(new_n315), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT25), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n306), .B1(new_n287), .B2(new_n289), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT68), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n305), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n295), .A2(KEYINPUT68), .A3(new_n304), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n323), .A2(new_n308), .A3(new_n325), .A4(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n296), .A2(new_n297), .A3(KEYINPUT23), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n314), .B1(G169gat), .B2(G176gat), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n328), .B(new_n329), .C1(new_n301), .C2(new_n300), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n330), .A2(new_n321), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n322), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n303), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT29), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n285), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G197gat), .B(G204gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT22), .ZN(new_n338));
  NAND2_X1  g137(.A1(G211gat), .A2(G218gat), .ZN(new_n339));
  INV_X1    g138(.A(G211gat), .ZN(new_n340));
  INV_X1    g139(.A(G218gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n338), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT22), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n339), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(new_n337), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n336), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT70), .ZN(new_n350));
  AOI221_X4 g149(.A(new_n350), .B1(new_n327), .B2(new_n331), .C1(new_n320), .C2(new_n321), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT70), .B1(new_n322), .B2(new_n332), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n303), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT74), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n303), .B(KEYINPUT74), .C1(new_n351), .C2(new_n352), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n349), .B1(new_n357), .B2(new_n285), .ZN(new_n358));
  AOI211_X1 g157(.A(KEYINPUT75), .B(new_n284), .C1(new_n355), .C2(new_n356), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n348), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n333), .A2(new_n350), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n322), .A2(new_n332), .A3(KEYINPUT70), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT74), .B1(new_n363), .B2(new_n303), .ZN(new_n364));
  INV_X1    g163(.A(new_n356), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n335), .B(new_n284), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n334), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(new_n285), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n366), .A2(new_n347), .A3(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G8gat), .B(G36gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(G64gat), .B(G92gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n360), .A2(new_n369), .A3(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT76), .B(KEYINPUT30), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n348), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n285), .B1(new_n364), .B2(new_n365), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT75), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n357), .A2(new_n349), .A3(new_n285), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n377), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n369), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n372), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n360), .A2(KEYINPUT30), .A3(new_n369), .A4(new_n373), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n376), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n283), .A2(new_n385), .A3(KEYINPUT35), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n353), .A2(new_n232), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n303), .B(new_n234), .C1(new_n351), .C2(new_n352), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(G227gat), .ZN(new_n390));
  INV_X1    g189(.A(G233gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT34), .B1(new_n389), .B2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(KEYINPUT64), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n395), .A2(KEYINPUT34), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n387), .A2(new_n388), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G15gat), .B(G43gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(G71gat), .B(G99gat), .ZN(new_n400));
  XOR2_X1   g199(.A(new_n399), .B(new_n400), .Z(new_n401));
  NAND2_X1  g200(.A1(new_n389), .A2(new_n395), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT72), .B(KEYINPUT33), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n398), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n394), .B1(new_n387), .B2(new_n388), .ZN(new_n406));
  INV_X1    g205(.A(new_n403), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n401), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n408), .A2(new_n393), .A3(new_n397), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT73), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n402), .A2(new_n411), .A3(KEYINPUT32), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT32), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT73), .B1(new_n406), .B2(new_n413), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n410), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n415), .A2(new_n405), .A3(new_n409), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(G228gat), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n246), .B1(new_n347), .B2(KEYINPUT29), .ZN(new_n421));
  AOI211_X1 g220(.A(new_n420), .B(new_n391), .C1(new_n421), .C2(new_n224), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n335), .B1(new_n224), .B2(KEYINPUT3), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n347), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT81), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n423), .A2(KEYINPUT81), .A3(new_n347), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n422), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n424), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT80), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n346), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n345), .A2(KEYINPUT80), .A3(new_n337), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n343), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n335), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n243), .B1(new_n434), .B2(new_n246), .ZN(new_n435));
  OAI22_X1  g234(.A1(new_n429), .A2(new_n435), .B1(new_n420), .B2(new_n391), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n428), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(G22gat), .ZN(new_n438));
  INV_X1    g237(.A(G22gat), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n428), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(KEYINPUT82), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(G78gat), .B(G106gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(KEYINPUT31), .B(G50gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n441), .B(new_n445), .C1(KEYINPUT82), .C2(new_n438), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n438), .A2(new_n444), .A3(new_n440), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT83), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n438), .A2(KEYINPUT83), .A3(new_n444), .A4(new_n440), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n446), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n419), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n386), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n274), .B1(new_n273), .B2(new_n281), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n376), .A2(new_n455), .A3(new_n383), .A4(new_n384), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT35), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n446), .A2(new_n449), .A3(new_n450), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT36), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n415), .A2(new_n405), .A3(new_n409), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n405), .A2(new_n409), .B1(new_n414), .B2(new_n412), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n417), .A2(KEYINPUT36), .A3(new_n418), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n460), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n233), .A2(new_n207), .A3(new_n235), .ZN(new_n468));
  OAI211_X1 g267(.A(KEYINPUT39), .B(new_n468), .C1(new_n263), .C2(new_n207), .ZN(new_n469));
  OR3_X1    g268(.A1(new_n263), .A2(KEYINPUT39), .A3(new_n207), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT84), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n470), .A2(new_n471), .A3(new_n270), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n471), .B1(new_n470), .B2(new_n270), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n469), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT40), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT40), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n476), .B(new_n469), .C1(new_n472), .C2(new_n473), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n278), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n459), .B1(new_n385), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT37), .B1(new_n360), .B2(new_n369), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n347), .B1(new_n366), .B2(new_n368), .ZN(new_n481));
  INV_X1    g280(.A(new_n336), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n482), .B1(new_n358), .B2(new_n359), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n481), .B1(new_n483), .B2(new_n347), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n480), .B1(KEYINPUT37), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT38), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n372), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n283), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT37), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n489), .B1(new_n381), .B2(new_n382), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n360), .A2(KEYINPUT37), .A3(new_n369), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n373), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n374), .B1(new_n492), .B2(new_n486), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n479), .B1(new_n488), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n467), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n458), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G15gat), .B(G22gat), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT16), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n498), .B1(new_n499), .B2(G1gat), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(G1gat), .B2(new_n498), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(G8gat), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NOR3_X1   g302(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n504), .B(KEYINPUT88), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n505), .A2(new_n506), .B1(G29gat), .B2(G36gat), .ZN(new_n507));
  INV_X1    g306(.A(G50gat), .ZN(new_n508));
  OR2_X1    g307(.A1(new_n508), .A2(G43gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(G43gat), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n509), .A2(KEYINPUT15), .A3(new_n510), .ZN(new_n511));
  XOR2_X1   g310(.A(KEYINPUT87), .B(G43gat), .Z(new_n512));
  OAI21_X1  g311(.A(new_n509), .B1(new_n512), .B2(G50gat), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT15), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n506), .ZN(new_n516));
  INV_X1    g315(.A(G29gat), .ZN(new_n517));
  INV_X1    g316(.A(G36gat), .ZN(new_n518));
  OAI22_X1  g317(.A1(new_n516), .A2(new_n504), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n507), .A2(new_n515), .B1(new_n519), .B2(new_n511), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n503), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT89), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n515), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n511), .A2(new_n519), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT17), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n522), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n520), .A2(KEYINPUT89), .A3(KEYINPUT17), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n502), .B1(new_n525), .B2(new_n526), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n521), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G229gat), .A2(G233gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT18), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT90), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n536), .B1(new_n525), .B2(new_n502), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n521), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n532), .B(KEYINPUT13), .ZN(new_n539));
  NOR3_X1   g338(.A1(new_n503), .A2(new_n520), .A3(new_n536), .ZN(new_n540));
  OR3_X1    g339(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n531), .A2(KEYINPUT18), .A3(new_n532), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n535), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G113gat), .B(G141gat), .ZN(new_n544));
  INV_X1    g343(.A(G197gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT11), .B(G169gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n548), .B(KEYINPUT12), .Z(new_n549));
  NAND2_X1  g348(.A1(new_n543), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n549), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n535), .A2(new_n541), .A3(new_n542), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G85gat), .A2(G92gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n555), .B(new_n556), .Z(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT94), .B(G92gat), .ZN(new_n558));
  INV_X1    g357(.A(G85gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(G99gat), .ZN(new_n561));
  INV_X1    g360(.A(G106gat), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT8), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n557), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G99gat), .B(G106gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G71gat), .B(G78gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(G57gat), .B(G64gat), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n567), .B1(new_n569), .B2(KEYINPUT9), .ZN(new_n570));
  XOR2_X1   g369(.A(G71gat), .B(G78gat), .Z(new_n571));
  INV_X1    g370(.A(KEYINPUT91), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n567), .A2(KEYINPUT91), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n568), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT9), .ZN(new_n576));
  INV_X1    g375(.A(G71gat), .ZN(new_n577));
  INV_X1    g376(.A(G78gat), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n570), .B1(new_n575), .B2(new_n579), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n566), .B(new_n580), .C1(KEYINPUT98), .C2(new_n565), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT10), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n580), .B1(KEYINPUT98), .B2(new_n565), .ZN(new_n583));
  INV_X1    g382(.A(new_n565), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n564), .B(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n581), .A2(new_n582), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n566), .A2(KEYINPUT10), .A3(new_n580), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G230gat), .A2(G233gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n581), .A2(new_n586), .ZN(new_n592));
  INV_X1    g391(.A(new_n590), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G120gat), .B(G148gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(G176gat), .B(G204gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n598), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n591), .A2(new_n594), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n554), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT97), .ZN(new_n605));
  XOR2_X1   g404(.A(G190gat), .B(G218gat), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT95), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n607), .A2(KEYINPUT96), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n525), .A2(new_n526), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n529), .A2(new_n609), .A3(new_n585), .ZN(new_n610));
  NAND2_X1  g409(.A1(G232gat), .A2(G233gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT92), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT41), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n614), .B1(new_n525), .B2(new_n566), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n608), .B1(new_n610), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n607), .A2(KEYINPUT96), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n605), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n616), .A2(new_n617), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n616), .A2(new_n617), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n621), .A2(KEYINPUT97), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n612), .A2(new_n613), .ZN(new_n624));
  XOR2_X1   g423(.A(G134gat), .B(G162gat), .Z(new_n625));
  XOR2_X1   g424(.A(new_n624), .B(new_n625), .Z(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n620), .A2(new_n623), .A3(new_n627), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n605), .B(new_n626), .C1(new_n618), .C2(new_n619), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n580), .A2(KEYINPUT21), .ZN(new_n631));
  OAI21_X1  g430(.A(G183gat), .B1(new_n631), .B2(new_n502), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n580), .A2(KEYINPUT21), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n503), .A2(new_n633), .A3(new_n306), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n632), .A2(new_n634), .A3(new_n636), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n580), .A2(KEYINPUT21), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G211gat), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n639), .A2(new_n641), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G127gat), .B(G155gat), .ZN(new_n646));
  NAND2_X1  g445(.A1(G231gat), .A2(G233gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n643), .B1(new_n638), .B2(new_n640), .ZN(new_n650));
  OR3_X1    g449(.A1(new_n645), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n649), .B1(new_n645), .B2(new_n650), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n630), .A2(new_n653), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n497), .A2(new_n604), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n455), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT99), .B(G1gat), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(G1324gat));
  XOR2_X1   g458(.A(KEYINPUT16), .B(G8gat), .Z(new_n660));
  NAND3_X1  g459(.A1(new_n655), .A2(new_n385), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n663), .A2(KEYINPUT100), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  INV_X1    g464(.A(new_n655), .ZN(new_n666));
  INV_X1    g465(.A(new_n385), .ZN(new_n667));
  OAI21_X1  g466(.A(G8gat), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n663), .A2(KEYINPUT100), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n664), .A2(new_n665), .A3(new_n668), .A4(new_n669), .ZN(G1325gat));
  AOI21_X1  g469(.A(G15gat), .B1(new_n655), .B2(new_n419), .ZN(new_n671));
  INV_X1    g470(.A(new_n466), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n671), .B1(new_n673), .B2(G15gat), .ZN(G1326gat));
  NAND2_X1  g473(.A1(new_n655), .A2(new_n459), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G22gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT101), .B(KEYINPUT43), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1327gat));
  INV_X1    g477(.A(new_n630), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n496), .A2(KEYINPUT44), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n467), .A2(new_n494), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n683), .B1(new_n467), .B2(new_n494), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n458), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n679), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n681), .B1(new_n682), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n604), .A2(new_n653), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(G29gat), .B1(new_n690), .B2(new_n455), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n496), .A2(new_n679), .A3(new_n689), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n692), .A2(new_n517), .A3(new_n656), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT45), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n691), .A2(new_n694), .ZN(G1328gat));
  OAI21_X1  g494(.A(G36gat), .B1(new_n690), .B2(new_n667), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n692), .A2(new_n518), .A3(new_n385), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n697), .B(KEYINPUT46), .Z(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(G1329gat));
  AND2_X1   g498(.A1(new_n454), .A2(new_n457), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n495), .A2(KEYINPUT102), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n467), .A2(new_n494), .A3(new_n683), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n682), .B1(new_n703), .B2(new_n630), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n704), .A2(new_n466), .A3(new_n689), .A4(new_n680), .ZN(new_n705));
  INV_X1    g504(.A(new_n512), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n512), .A3(new_n419), .ZN(new_n708));
  AOI21_X1  g507(.A(KEYINPUT103), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n709), .B(new_n711), .ZN(G1330gat));
  NAND4_X1  g511(.A1(new_n704), .A2(new_n459), .A3(new_n689), .A4(new_n680), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT48), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n713), .A2(new_n714), .A3(G50gat), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n692), .A2(new_n508), .A3(new_n459), .ZN(new_n716));
  NAND2_X1  g515(.A1(KEYINPUT105), .A2(KEYINPUT48), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n713), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n688), .A2(KEYINPUT106), .A3(new_n459), .A4(new_n689), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(new_n721), .A3(G50gat), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n692), .A2(KEYINPUT105), .A3(new_n508), .A4(new_n459), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n718), .B1(new_n724), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g524(.A1(new_n703), .A2(new_n553), .ZN(new_n726));
  INV_X1    g525(.A(new_n602), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n654), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n656), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g531(.A1(new_n729), .A2(new_n667), .ZN(new_n733));
  NOR2_X1   g532(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n734));
  AND2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(new_n733), .B2(new_n734), .ZN(G1333gat));
  NAND3_X1  g536(.A1(new_n730), .A2(new_n577), .A3(new_n419), .ZN(new_n738));
  OAI21_X1  g537(.A(G71gat), .B1(new_n729), .B2(new_n672), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT50), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(G1334gat));
  NOR2_X1   g541(.A1(new_n729), .A2(new_n451), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(new_n578), .ZN(G1335gat));
  NOR2_X1   g543(.A1(new_n653), .A2(new_n553), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n704), .A2(new_n602), .A3(new_n680), .A4(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(G85gat), .B1(new_n746), .B2(new_n455), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n686), .A2(new_n679), .A3(new_n745), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT51), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n686), .A2(KEYINPUT51), .A3(new_n679), .A4(new_n745), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n656), .A2(new_n559), .A3(new_n602), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT107), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n747), .B1(new_n753), .B2(new_n755), .ZN(G1336gat));
  NOR2_X1   g555(.A1(new_n667), .A2(G92gat), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n752), .A2(KEYINPUT108), .A3(new_n602), .A4(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n558), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(new_n746), .B2(new_n667), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n727), .B1(new_n750), .B2(new_n751), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT108), .B1(new_n762), .B2(new_n757), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT52), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n752), .A2(new_n602), .A3(new_n757), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n762), .A2(KEYINPUT109), .A3(new_n757), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n767), .A2(new_n768), .A3(new_n760), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n764), .A2(new_n770), .ZN(G1337gat));
  AOI21_X1  g570(.A(G99gat), .B1(new_n762), .B2(new_n419), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n746), .A2(new_n561), .A3(new_n672), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(G1338gat));
  NAND4_X1  g573(.A1(new_n752), .A2(new_n562), .A3(new_n602), .A4(new_n459), .ZN(new_n775));
  OAI21_X1  g574(.A(G106gat), .B1(new_n746), .B2(new_n451), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n777), .A2(new_n779), .A3(KEYINPUT53), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n775), .B(new_n776), .C1(new_n778), .C2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(G1339gat));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n784));
  INV_X1    g583(.A(new_n532), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n529), .A2(new_n530), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n784), .B(new_n785), .C1(new_n786), .C2(new_n521), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT112), .B1(new_n531), .B2(new_n532), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n539), .B1(new_n538), .B2(new_n540), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n548), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n791), .A2(new_n552), .A3(new_n602), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n587), .A2(new_n593), .A3(new_n588), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n591), .A2(KEYINPUT54), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n593), .B1(new_n587), .B2(new_n588), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n600), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n794), .A2(KEYINPUT55), .A3(new_n797), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n798), .A2(new_n601), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n793), .A2(KEYINPUT54), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(new_n795), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n589), .A2(new_n796), .A3(new_n590), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n598), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n800), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT111), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g606(.A(KEYINPUT111), .B(new_n800), .C1(new_n802), .C2(new_n804), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n799), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n792), .B1(new_n809), .B2(new_n554), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n630), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n791), .A2(new_n552), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n628), .A2(new_n812), .A3(new_n629), .ZN(new_n813));
  INV_X1    g612(.A(new_n809), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n653), .B1(new_n811), .B2(new_n815), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n630), .A2(new_n554), .A3(new_n727), .A4(new_n653), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT113), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n385), .A2(new_n455), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n821));
  AOI22_X1  g620(.A1(new_n630), .A2(new_n810), .B1(new_n813), .B2(new_n814), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n821), .B(new_n817), .C1(new_n822), .C2(new_n653), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n819), .A2(new_n453), .A3(new_n820), .A4(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n553), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n602), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g628(.A1(new_n825), .A2(new_n653), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g630(.A1(new_n825), .A2(new_n679), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n832), .A2(KEYINPUT56), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n833), .A2(G134gat), .ZN(new_n834));
  OR3_X1    g633(.A1(new_n832), .A2(KEYINPUT114), .A3(KEYINPUT56), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT114), .B1(new_n832), .B2(KEYINPUT56), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n834), .B(new_n837), .ZN(G1343gat));
  NAND2_X1  g637(.A1(new_n672), .A2(new_n820), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n819), .A2(new_n841), .A3(new_n459), .A4(new_n823), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n553), .A2(new_n799), .A3(new_n805), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n792), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n791), .A2(KEYINPUT115), .A3(new_n602), .A4(new_n552), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n843), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n630), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n815), .ZN(new_n849));
  INV_X1    g648(.A(new_n653), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT116), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n653), .B1(new_n848), .B2(new_n815), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n818), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n451), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n840), .B(new_n842), .C1(new_n856), .C2(new_n841), .ZN(new_n857));
  OAI21_X1  g656(.A(G141gat), .B1(new_n857), .B2(new_n554), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n819), .A2(new_n459), .A3(new_n823), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(new_n839), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n554), .A2(G141gat), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n863), .A2(KEYINPUT118), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(KEYINPUT118), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n862), .A2(KEYINPUT119), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  OAI211_X1 g665(.A(KEYINPUT117), .B(G141gat), .C1(new_n857), .C2(new_n554), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n860), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT58), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n862), .A2(new_n864), .A3(new_n865), .ZN(new_n870));
  NAND2_X1  g669(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n870), .B(new_n871), .C1(new_n858), .C2(KEYINPUT58), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n869), .A2(new_n872), .ZN(G1344gat));
  INV_X1    g672(.A(KEYINPUT59), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n874), .B(G148gat), .C1(new_n857), .C2(new_n727), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n817), .B(KEYINPUT120), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT57), .B1(new_n851), .B2(new_n877), .ZN(new_n878));
  AOI22_X1  g677(.A1(new_n861), .A2(KEYINPUT57), .B1(new_n459), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(new_n602), .A3(new_n840), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(G148gat), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n876), .B1(new_n881), .B2(KEYINPUT59), .ZN(new_n882));
  AOI211_X1 g681(.A(KEYINPUT121), .B(new_n874), .C1(new_n880), .C2(G148gat), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n875), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(G148gat), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n862), .A2(new_n885), .A3(new_n602), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(G1345gat));
  AND2_X1   g686(.A1(new_n211), .A2(new_n213), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n888), .B1(new_n862), .B2(new_n653), .ZN(new_n889));
  INV_X1    g688(.A(new_n857), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n653), .A2(new_n888), .ZN(new_n891));
  XOR2_X1   g690(.A(new_n891), .B(KEYINPUT122), .Z(new_n892));
  AOI21_X1  g691(.A(new_n889), .B1(new_n890), .B2(new_n892), .ZN(G1346gat));
  AOI21_X1  g692(.A(G162gat), .B1(new_n862), .B2(new_n679), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n890), .A2(G162gat), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n894), .B1(new_n895), .B2(new_n679), .ZN(G1347gat));
  AND2_X1   g695(.A1(new_n819), .A2(new_n823), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n667), .A2(new_n656), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n897), .A2(new_n453), .A3(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n553), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(G169gat), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n316), .A2(new_n317), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(new_n901), .B2(new_n903), .ZN(G1348gat));
  NOR2_X1   g703(.A1(new_n899), .A2(new_n727), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(new_n297), .ZN(G1349gat));
  AOI21_X1  g705(.A(new_n306), .B1(new_n900), .B2(new_n653), .ZN(new_n907));
  INV_X1    g706(.A(new_n291), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n899), .A2(new_n908), .A3(new_n850), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g709(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n910), .B(new_n911), .ZN(G1350gat));
  OAI21_X1  g711(.A(G190gat), .B1(new_n899), .B2(new_n630), .ZN(new_n913));
  XOR2_X1   g712(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n290), .A3(new_n679), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n913), .A2(new_n915), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(G1351gat));
  INV_X1    g718(.A(new_n861), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n672), .A2(new_n898), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n924), .A2(new_n545), .A3(new_n553), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n879), .A2(new_n553), .A3(new_n922), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n926), .B2(new_n545), .ZN(G1352gat));
  INV_X1    g726(.A(G204gat), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n924), .A2(new_n928), .A3(new_n602), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n929), .A2(KEYINPUT62), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(KEYINPUT62), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n879), .A2(new_n602), .A3(new_n922), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n930), .B(new_n931), .C1(new_n928), .C2(new_n932), .ZN(G1353gat));
  NAND3_X1  g732(.A1(new_n924), .A2(new_n340), .A3(new_n653), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n861), .A2(KEYINPUT57), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n878), .A2(new_n459), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n935), .A2(new_n653), .A3(new_n936), .A4(new_n922), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT125), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n879), .A2(KEYINPUT125), .A3(new_n653), .A4(new_n922), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n939), .A2(G211gat), .A3(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT63), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n934), .B1(new_n943), .B2(new_n944), .ZN(G1354gat));
  OAI21_X1  g744(.A(new_n341), .B1(new_n923), .B2(new_n630), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n679), .A2(G218gat), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT126), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n879), .A2(new_n922), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


