//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 1 0 0 0 1 0 1 1 1 0 1 0 0 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 1 1 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n231, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1262, new_n1263, new_n1264, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1316, new_n1317,
    new_n1318, new_n1319;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT0), .ZN(new_n206));
  OAI21_X1  g0006(.A(G50), .B1(G58), .B2(G68), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT64), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n217));
  NAND3_X1  g0017(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n203), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n206), .B(new_n212), .C1(new_n219), .C2(KEYINPUT1), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n220), .B1(KEYINPUT1), .B2(new_n219), .ZN(G361));
  XOR2_X1   g0021(.A(G238), .B(G244), .Z(new_n222));
  XNOR2_X1  g0022(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n222), .B(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(G226), .B(G232), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(G250), .B(G257), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G264), .B(G270), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n226), .B(new_n229), .ZN(G358));
  XNOR2_X1  g0030(.A(G50), .B(G58), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT66), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G68), .B(G77), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XOR2_X1   g0035(.A(G107), .B(G116), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G351));
  INV_X1    g0038(.A(KEYINPUT13), .ZN(new_n239));
  NAND2_X1  g0039(.A1(G33), .A2(G41), .ZN(new_n240));
  NAND3_X1  g0040(.A1(new_n240), .A2(G1), .A3(G13), .ZN(new_n241));
  INV_X1    g0041(.A(new_n241), .ZN(new_n242));
  AND2_X1   g0042(.A1(KEYINPUT3), .A2(G33), .ZN(new_n243));
  NOR2_X1   g0043(.A1(KEYINPUT3), .A2(G33), .ZN(new_n244));
  NOR2_X1   g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G1698), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(KEYINPUT68), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT68), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G1698), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n247), .A2(new_n249), .A3(G226), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G232), .A2(G1698), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n245), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G97), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n242), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n241), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G274), .ZN(new_n260));
  INV_X1    g0060(.A(new_n209), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n260), .B1(new_n261), .B2(new_n240), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  INV_X1    g0063(.A(G45), .ZN(new_n264));
  AOI21_X1  g0064(.A(G1), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n259), .A2(G238), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n239), .B1(new_n255), .B2(new_n266), .ZN(new_n267));
  AND3_X1   g0067(.A1(new_n255), .A2(new_n239), .A3(new_n266), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT74), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n255), .A2(new_n239), .A3(new_n266), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT74), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n270), .A2(G190), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n255), .A2(new_n266), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT13), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n271), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G200), .ZN(new_n277));
  INV_X1    g0077(.A(G13), .ZN(new_n278));
  NOR3_X1   g0078(.A1(new_n278), .A2(new_n210), .A3(G1), .ZN(new_n279));
  INV_X1    g0079(.A(G68), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(new_n281), .B(KEYINPUT12), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G20), .A2(G33), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n283), .A2(G50), .B1(G20), .B2(new_n280), .ZN(new_n284));
  INV_X1    g0084(.A(G77), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n210), .A2(G33), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n209), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n287), .A2(KEYINPUT11), .A3(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n279), .A2(new_n289), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n256), .A2(G20), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(G68), .A3(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n282), .A2(new_n290), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(KEYINPUT11), .B1(new_n287), .B2(new_n289), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n273), .A2(new_n277), .A3(new_n296), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n270), .A2(KEYINPUT75), .A3(G179), .A4(new_n272), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n255), .A2(new_n269), .A3(new_n239), .A4(new_n266), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n272), .A2(new_n275), .A3(G179), .A4(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT75), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT14), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n304), .B1(new_n276), .B2(G169), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n304), .B(G169), .C1(new_n268), .C2(new_n267), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n296), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n297), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT16), .ZN(new_n312));
  OR2_X1    g0112(.A1(KEYINPUT3), .A2(G33), .ZN(new_n313));
  NAND2_X1  g0113(.A1(KEYINPUT3), .A2(G33), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n313), .A2(new_n210), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT7), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n313), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n314), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n280), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G58), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(new_n280), .ZN(new_n321));
  NOR2_X1   g0121(.A1(G58), .A2(G68), .ZN(new_n322));
  OAI21_X1  g0122(.A(G20), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n283), .A2(G159), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n312), .B1(new_n319), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(KEYINPUT7), .B1(new_n245), .B2(new_n210), .ZN(new_n327));
  NOR4_X1   g0127(.A1(new_n243), .A2(new_n244), .A3(new_n316), .A4(G20), .ZN(new_n328));
  OAI21_X1  g0128(.A(G68), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n325), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n329), .A2(KEYINPUT16), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n326), .A2(new_n331), .A3(new_n289), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT76), .ZN(new_n333));
  XNOR2_X1  g0133(.A(KEYINPUT8), .B(G58), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n279), .ZN(new_n335));
  INV_X1    g0135(.A(new_n334), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n292), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n288), .A2(new_n209), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n278), .A2(G1), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G20), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n333), .B(new_n335), .C1(new_n337), .C2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n291), .A2(new_n292), .A3(new_n336), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n333), .B1(new_n344), .B2(new_n335), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n332), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n265), .A2(new_n241), .A3(G274), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n241), .A2(G232), .A3(new_n257), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI211_X1 g0150(.A(G226), .B(G1698), .C1(new_n243), .C2(new_n244), .ZN(new_n351));
  NAND2_X1  g0151(.A1(G33), .A2(G87), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n247), .B(new_n249), .C1(new_n243), .C2(new_n244), .ZN(new_n353));
  INV_X1    g0153(.A(G223), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n351), .B(new_n352), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n350), .B1(new_n355), .B2(new_n242), .ZN(new_n356));
  INV_X1    g0156(.A(G190), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(G200), .B2(new_n356), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n347), .A2(KEYINPUT17), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(new_n332), .A3(new_n346), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT17), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT78), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n332), .A2(new_n346), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT77), .ZN(new_n367));
  INV_X1    g0167(.A(G179), .ZN(new_n368));
  AOI211_X1 g0168(.A(new_n368), .B(new_n350), .C1(new_n355), .C2(new_n242), .ZN(new_n369));
  INV_X1    g0169(.A(G169), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n355), .A2(new_n242), .ZN(new_n371));
  INV_X1    g0171(.A(new_n350), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n367), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n356), .A2(G179), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n375), .B(KEYINPUT77), .C1(new_n370), .C2(new_n356), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT18), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n366), .A2(new_n374), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n366), .A2(new_n374), .A3(new_n376), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT18), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n364), .A2(new_n365), .A3(new_n378), .A4(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n380), .A2(new_n378), .A3(new_n363), .A4(new_n360), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT78), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT73), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n384), .A2(KEYINPUT10), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n241), .A2(G226), .A3(new_n257), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n348), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT67), .ZN(new_n388));
  XNOR2_X1  g0188(.A(new_n387), .B(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n313), .A2(new_n314), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G1698), .ZN(new_n391));
  OAI22_X1  g0191(.A1(new_n391), .A2(new_n354), .B1(new_n285), .B2(new_n390), .ZN(new_n392));
  XNOR2_X1  g0192(.A(KEYINPUT68), .B(G1698), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT69), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n390), .A2(new_n393), .A3(new_n394), .A4(G222), .ZN(new_n395));
  INV_X1    g0195(.A(G222), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT69), .B1(new_n353), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n392), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n389), .B(G190), .C1(new_n398), .C2(new_n241), .ZN(new_n399));
  INV_X1    g0199(.A(G50), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n400), .B1(new_n256), .B2(G20), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n291), .A2(new_n401), .B1(new_n400), .B2(new_n279), .ZN(new_n402));
  INV_X1    g0202(.A(G150), .ZN(new_n403));
  INV_X1    g0203(.A(new_n283), .ZN(new_n404));
  OAI22_X1  g0204(.A1(new_n334), .A2(new_n286), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(G50), .A2(G58), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n210), .B1(new_n406), .B2(new_n280), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n402), .B1(new_n408), .B2(new_n338), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT9), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n409), .A2(new_n410), .B1(new_n384), .B2(KEYINPUT10), .ZN(new_n411));
  OAI211_X1 g0211(.A(KEYINPUT9), .B(new_n402), .C1(new_n408), .C2(new_n338), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n399), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  XNOR2_X1  g0213(.A(KEYINPUT72), .B(G200), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n397), .A2(new_n395), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n246), .B1(new_n313), .B2(new_n314), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n416), .A2(G223), .B1(new_n245), .B2(G77), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n242), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n414), .B1(new_n419), .B2(new_n389), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n385), .B1(new_n413), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n409), .A2(new_n410), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n384), .A2(KEYINPUT10), .ZN(new_n423));
  AND3_X1   g0223(.A1(new_n422), .A2(new_n412), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n419), .A2(new_n389), .ZN(new_n425));
  INV_X1    g0225(.A(new_n414), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n385), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n424), .A2(new_n427), .A3(new_n428), .A4(new_n399), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n425), .A2(new_n370), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n430), .B(new_n409), .C1(G179), .C2(new_n425), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n421), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n291), .A2(G77), .A3(new_n292), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(G77), .B2(new_n340), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n334), .A2(new_n404), .B1(new_n210), .B2(new_n285), .ZN(new_n435));
  XNOR2_X1  g0235(.A(KEYINPUT15), .B(G87), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n436), .A2(new_n286), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n289), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT70), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g0240(.A(KEYINPUT70), .B(new_n289), .C1(new_n435), .C2(new_n437), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n434), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n442), .A2(KEYINPUT71), .ZN(new_n443));
  INV_X1    g0243(.A(G244), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n348), .B1(new_n444), .B2(new_n258), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n245), .A2(G107), .ZN(new_n446));
  OAI211_X1 g0246(.A(G238), .B(G1698), .C1(new_n243), .C2(new_n244), .ZN(new_n447));
  INV_X1    g0247(.A(G232), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n446), .B(new_n447), .C1(new_n448), .C2(new_n353), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n445), .B1(new_n449), .B2(new_n242), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(G190), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(new_n414), .B2(new_n450), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n443), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n442), .A2(KEYINPUT71), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n450), .A2(G169), .ZN(new_n456));
  AOI211_X1 g0256(.A(G179), .B(new_n445), .C1(new_n449), .C2(new_n242), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n442), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n432), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n311), .A2(new_n381), .A3(new_n383), .A4(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT79), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n458), .B1(new_n453), .B2(new_n454), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n464), .A2(new_n421), .A3(new_n429), .A4(new_n431), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n465), .B1(KEYINPUT78), .B2(new_n382), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT79), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n466), .A2(new_n467), .A3(new_n311), .A4(new_n381), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT4), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n470), .B1(new_n353), .B2(new_n444), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n390), .A2(new_n393), .A3(KEYINPUT4), .A4(G244), .ZN(new_n472));
  NAND2_X1  g0272(.A1(G33), .A2(G283), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(KEYINPUT83), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT83), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n475), .A2(G33), .A3(G283), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g0277(.A(G250), .B(G1698), .C1(new_n243), .C2(new_n244), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n471), .A2(new_n472), .A3(new_n477), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n242), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n264), .A2(G1), .ZN(new_n481));
  NOR2_X1   g0281(.A1(KEYINPUT5), .A2(G41), .ZN(new_n482));
  AND2_X1   g0282(.A1(KEYINPUT5), .A2(G41), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n262), .B(new_n481), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n481), .B1(new_n483), .B2(new_n482), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(G257), .A3(new_n241), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n480), .A2(G190), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT84), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n256), .A2(G33), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n338), .A2(new_n340), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT82), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT82), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n291), .A2(new_n494), .A3(new_n491), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n493), .A2(new_n495), .A3(G97), .ZN(new_n496));
  INV_X1    g0296(.A(G97), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n279), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g0298(.A(new_n498), .B(KEYINPUT81), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(G107), .B1(new_n327), .B2(new_n328), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT80), .ZN(new_n502));
  INV_X1    g0302(.A(G107), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(new_n317), .B2(new_n318), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT80), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT6), .ZN(new_n507));
  AND2_X1   g0307(.A1(G97), .A2(G107), .ZN(new_n508));
  NOR2_X1   g0308(.A1(G97), .A2(G107), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n503), .A2(KEYINPUT6), .A3(G97), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n512), .A2(G20), .B1(G77), .B2(new_n283), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n502), .A2(new_n506), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n500), .B1(new_n514), .B2(new_n289), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n480), .A2(new_n488), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(G200), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n487), .B1(new_n479), .B2(new_n242), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT84), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(new_n519), .A3(G190), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n490), .A2(new_n515), .A3(new_n517), .A4(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n478), .A2(new_n477), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n390), .A2(new_n393), .A3(G244), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n522), .B1(new_n470), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n241), .B1(new_n524), .B2(new_n472), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n370), .B1(new_n525), .B2(new_n487), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n518), .A2(new_n368), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n283), .A2(G77), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n503), .A2(KEYINPUT6), .A3(G97), .ZN(new_n529));
  XNOR2_X1  g0329(.A(G97), .B(G107), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n529), .B1(new_n530), .B2(new_n507), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n528), .B1(new_n531), .B2(new_n210), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(KEYINPUT80), .B2(new_n501), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n338), .B1(new_n533), .B2(new_n506), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n526), .B(new_n527), .C1(new_n534), .C2(new_n500), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n521), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT85), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT19), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n210), .B1(new_n253), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(G87), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n509), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n210), .B(G68), .C1(new_n243), .C2(new_n244), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n539), .B1(new_n286), .B2(new_n497), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT86), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n338), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n543), .A2(new_n544), .A3(KEYINPUT86), .A4(new_n545), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n548), .A2(new_n549), .B1(new_n279), .B2(new_n436), .ZN(new_n550));
  INV_X1    g0350(.A(new_n436), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n493), .A2(new_n495), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(G33), .ZN(new_n554));
  INV_X1    g0354(.A(G116), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n556), .B1(new_n416), .B2(G244), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n390), .A2(new_n393), .A3(G238), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n241), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n241), .A2(G274), .A3(new_n481), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n256), .A2(G45), .ZN(new_n561));
  AND2_X1   g0361(.A1(G33), .A2(G41), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n561), .B(G250), .C1(new_n562), .C2(new_n209), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(G169), .B1(new_n559), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(G244), .B(G1698), .C1(new_n243), .C2(new_n244), .ZN(new_n566));
  INV_X1    g0366(.A(new_n556), .ZN(new_n567));
  INV_X1    g0367(.A(G238), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n566), .B(new_n567), .C1(new_n353), .C2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n564), .B1(new_n569), .B2(new_n242), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G179), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n553), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(G257), .B(G1698), .C1(new_n243), .C2(new_n244), .ZN(new_n574));
  NAND2_X1  g0374(.A1(G33), .A2(G294), .ZN(new_n575));
  OAI21_X1  g0375(.A(G250), .B1(new_n243), .B2(new_n244), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n247), .A2(new_n249), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n574), .B(new_n575), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n242), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n485), .A2(G264), .A3(new_n241), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n579), .A2(new_n484), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n581), .A2(KEYINPUT90), .A3(G169), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT91), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n485), .A2(KEYINPUT91), .A3(G264), .A4(new_n241), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n584), .A2(new_n585), .B1(new_n578), .B2(new_n242), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n586), .A2(G179), .A3(new_n484), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT90), .B1(new_n581), .B2(G169), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n210), .B(G87), .C1(new_n243), .C2(new_n244), .ZN(new_n590));
  XNOR2_X1  g0390(.A(KEYINPUT89), .B(KEYINPUT22), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT22), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n593), .A2(KEYINPUT89), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n390), .A2(new_n210), .A3(G87), .A4(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT23), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n210), .B2(G107), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n503), .A2(KEYINPUT23), .A3(G20), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n597), .A2(new_n598), .B1(new_n556), .B2(new_n210), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n592), .A2(new_n595), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT24), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT24), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n592), .A2(new_n595), .A3(new_n599), .A4(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n338), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n340), .A2(G107), .ZN(new_n605));
  XNOR2_X1  g0405(.A(new_n605), .B(KEYINPUT25), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n493), .A2(new_n495), .A3(G107), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI22_X1  g0408(.A1(new_n588), .A2(new_n589), .B1(new_n604), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n426), .B1(new_n559), .B2(new_n564), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n493), .A2(new_n495), .A3(G87), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n569), .A2(new_n242), .ZN(new_n612));
  INV_X1    g0412(.A(new_n564), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(G190), .A3(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n550), .A2(new_n610), .A3(new_n611), .A4(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n604), .ZN(new_n616));
  INV_X1    g0416(.A(new_n608), .ZN(new_n617));
  AOI21_X1  g0417(.A(G200), .B1(new_n586), .B2(new_n484), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n581), .A2(G190), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n616), .B(new_n617), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  AND4_X1   g0420(.A1(new_n573), .A2(new_n609), .A3(new_n615), .A4(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n279), .A2(new_n555), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n492), .B2(new_n555), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n210), .B1(new_n497), .B2(G33), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n477), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(KEYINPUT87), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT87), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n477), .A2(new_n628), .A3(new_n625), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n338), .B1(G20), .B2(new_n555), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n627), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g0431(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n632));
  AOI21_X1  g0432(.A(new_n623), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(KEYINPUT88), .A2(KEYINPUT20), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n627), .A2(new_n634), .A3(new_n630), .A4(new_n629), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n242), .B1(new_n390), .B2(G303), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n245), .B1(G264), .B2(G1698), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n393), .A2(G257), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n485), .A2(G270), .A3(new_n241), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n484), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n643), .A2(new_n370), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n636), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT21), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n640), .A2(new_n642), .A3(new_n368), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n636), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n636), .A2(new_n644), .A3(KEYINPUT21), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n643), .A2(G190), .ZN(new_n651));
  OAI21_X1  g0451(.A(G200), .B1(new_n640), .B2(new_n642), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n651), .A2(new_n633), .A3(new_n635), .A4(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n647), .A2(new_n649), .A3(new_n650), .A4(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n521), .A2(new_n535), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n654), .B1(KEYINPUT85), .B2(new_n655), .ZN(new_n656));
  AND4_X1   g0456(.A1(new_n469), .A2(new_n538), .A3(new_n621), .A4(new_n656), .ZN(G372));
  AND4_X1   g0457(.A1(new_n550), .A2(new_n610), .A3(new_n611), .A4(new_n614), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT92), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n570), .A2(new_n370), .ZN(new_n660));
  AOI211_X1 g0460(.A(new_n368), .B(new_n564), .C1(new_n569), .C2(new_n242), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n565), .A2(new_n571), .A3(KEYINPUT92), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n658), .B1(new_n664), .B2(new_n553), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  INV_X1    g0466(.A(new_n535), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n660), .A2(new_n661), .A3(new_n659), .ZN(new_n669));
  AOI21_X1  g0469(.A(KEYINPUT92), .B1(new_n565), .B2(new_n571), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n553), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n518), .A2(G169), .ZN(new_n672));
  AOI211_X1 g0472(.A(G179), .B(new_n487), .C1(new_n479), .C2(new_n242), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n513), .B1(new_n504), .B2(new_n505), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n501), .A2(KEYINPUT80), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n289), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n500), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n674), .A2(new_n679), .A3(new_n573), .A4(new_n615), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(KEYINPUT26), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n668), .A2(new_n671), .A3(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n609), .A2(new_n647), .A3(new_n649), .A4(new_n650), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n665), .A2(new_n535), .A3(new_n521), .A4(new_n620), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT93), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n521), .A2(new_n535), .A3(new_n620), .ZN(new_n687));
  AOI21_X1  g0487(.A(KEYINPUT93), .B1(new_n687), .B2(new_n665), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n682), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n469), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT94), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n375), .B1(new_n370), .B2(new_n356), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n366), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT18), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n366), .A2(new_n377), .A3(new_n692), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n309), .A2(new_n310), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n297), .B2(new_n459), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n696), .B1(new_n698), .B2(new_n364), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n421), .A2(new_n429), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n431), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n691), .A2(new_n702), .ZN(G369));
  AND3_X1   g0503(.A1(new_n647), .A2(new_n649), .A3(new_n650), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n339), .A2(new_n210), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n705), .A2(KEYINPUT27), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(KEYINPUT27), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(new_n707), .A3(G213), .ZN(new_n708));
  INV_X1    g0508(.A(G343), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n636), .A2(new_n710), .ZN(new_n711));
  MUX2_X1   g0511(.A(new_n704), .B(new_n654), .S(new_n711), .Z(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT95), .ZN(new_n713));
  INV_X1    g0513(.A(new_n609), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n710), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n710), .B1(new_n604), .B2(new_n608), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n609), .A2(new_n620), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n713), .A2(G330), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n647), .A2(new_n649), .A3(new_n650), .ZN(new_n720));
  INV_X1    g0520(.A(new_n710), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n609), .A2(new_n620), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n724), .B1(new_n714), .B2(new_n721), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n719), .A2(new_n725), .ZN(G399));
  NOR2_X1   g0526(.A1(new_n542), .A2(G116), .ZN(new_n727));
  XOR2_X1   g0527(.A(new_n727), .B(KEYINPUT96), .Z(new_n728));
  INV_X1    g0528(.A(new_n204), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G41), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n728), .A2(new_n256), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n731), .B1(new_n208), .B2(new_n730), .ZN(new_n732));
  XOR2_X1   g0532(.A(new_n732), .B(KEYINPUT28), .Z(new_n733));
  INV_X1    g0533(.A(new_n671), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n490), .A2(new_n520), .ZN(new_n735));
  INV_X1    g0535(.A(G200), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n677), .B(new_n678), .C1(new_n736), .C2(new_n518), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n535), .B(new_n620), .C1(new_n735), .C2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n671), .A2(new_n615), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n734), .B1(new_n740), .B2(new_n683), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n665), .A2(KEYINPUT97), .A3(new_n667), .A4(KEYINPUT26), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n665), .A2(KEYINPUT26), .A3(new_n667), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT97), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n744), .B1(new_n680), .B2(new_n666), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n742), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n741), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n747), .A2(KEYINPUT29), .A3(new_n721), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n684), .A2(new_n685), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n687), .A2(KEYINPUT93), .A3(new_n665), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n749), .A2(new_n750), .A3(new_n683), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n710), .B1(new_n751), .B2(new_n682), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n748), .B1(new_n752), .B2(KEYINPUT29), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(G330), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n656), .A2(new_n538), .A3(new_n621), .A4(new_n721), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n586), .A2(new_n570), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(new_n518), .A3(new_n648), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT30), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n757), .A2(new_n648), .A3(KEYINPUT30), .A4(new_n518), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n643), .A2(G179), .A3(new_n570), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n586), .A2(new_n484), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n762), .A2(new_n516), .A3(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n760), .A2(new_n761), .A3(new_n764), .ZN(new_n765));
  AND3_X1   g0565(.A1(new_n765), .A2(KEYINPUT31), .A3(new_n710), .ZN(new_n766));
  AOI21_X1  g0566(.A(KEYINPUT31), .B1(new_n765), .B2(new_n710), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n755), .B1(new_n756), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n754), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n733), .B1(new_n770), .B2(G1), .ZN(G364));
  NAND2_X1  g0571(.A1(new_n713), .A2(G330), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n278), .A2(G20), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n256), .B1(new_n773), .B2(G45), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n730), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n772), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n713), .A2(G330), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G13), .A2(G33), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(G20), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n712), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n729), .A2(new_n245), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT98), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G355), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(G116), .B2(new_n204), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n234), .A2(G45), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n788), .B(KEYINPUT99), .Z(new_n789));
  NOR2_X1   g0589(.A1(new_n729), .A2(new_n390), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(new_n264), .B2(new_n208), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n787), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(G20), .B1(KEYINPUT100), .B2(G169), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(KEYINPUT100), .A2(G169), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n209), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n782), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n776), .B1(new_n793), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT101), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n797), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n210), .A2(new_n368), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n804), .A2(G190), .A3(new_n736), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n390), .B1(new_n805), .B2(new_n320), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n210), .A2(G190), .ZN(new_n807));
  NOR2_X1   g0607(.A1(G179), .A2(G200), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G159), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT32), .ZN(new_n812));
  INV_X1    g0612(.A(new_n807), .ZN(new_n813));
  NOR3_X1   g0613(.A1(new_n813), .A2(new_n368), .A3(G200), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n806), .B(new_n812), .C1(G77), .C2(new_n814), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n414), .A2(new_n813), .A3(G179), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT102), .Z(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(G107), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n804), .A2(G200), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(G190), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(new_n357), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n820), .A2(G68), .B1(new_n821), .B2(G50), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n210), .B1(new_n808), .B2(G190), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(G97), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  NOR4_X1   g0626(.A1(new_n414), .A2(new_n210), .A3(G179), .A4(new_n357), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(G87), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n815), .A2(new_n818), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n821), .ZN(new_n830));
  INV_X1    g0630(.A(G326), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n820), .ZN(new_n833));
  OR2_X1    g0633(.A1(KEYINPUT33), .A2(G317), .ZN(new_n834));
  NAND2_X1  g0634(.A1(KEYINPUT33), .A2(G317), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n832), .B(new_n836), .C1(G294), .C2(new_n824), .ZN(new_n837));
  INV_X1    g0637(.A(new_n805), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n838), .A2(G322), .B1(new_n810), .B2(G329), .ZN(new_n839));
  INV_X1    g0639(.A(G311), .ZN(new_n840));
  INV_X1    g0640(.A(new_n814), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n839), .B(new_n245), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(G303), .B2(new_n827), .ZN(new_n843));
  INV_X1    g0643(.A(G283), .ZN(new_n844));
  INV_X1    g0644(.A(new_n817), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n837), .B(new_n843), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n803), .B1(new_n829), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(new_n800), .B2(new_n801), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n802), .A2(new_n848), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n778), .A2(new_n779), .B1(new_n783), .B2(new_n849), .ZN(G396));
  NAND2_X1  g0650(.A1(new_n458), .A2(new_n721), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n455), .B1(new_n442), .B2(new_n721), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n852), .B1(new_n853), .B2(new_n459), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n668), .A2(new_n671), .A3(new_n681), .ZN(new_n855));
  INV_X1    g0655(.A(new_n683), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(new_n740), .B2(KEYINPUT93), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n855), .B1(new_n857), .B2(new_n749), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n460), .A2(new_n710), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n752), .A2(new_n854), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n769), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n776), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n862), .B2(new_n861), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n797), .A2(new_n780), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n777), .B1(new_n865), .B2(new_n285), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n814), .A2(G159), .B1(new_n838), .B2(G143), .ZN(new_n867));
  INV_X1    g0667(.A(G137), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n867), .B1(new_n868), .B2(new_n830), .C1(new_n403), .C2(new_n833), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n869), .B(KEYINPUT34), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n817), .A2(G68), .ZN(new_n871));
  INV_X1    g0671(.A(G132), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n390), .B1(new_n823), .B2(new_n320), .C1(new_n872), .C2(new_n809), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(G50), .B2(new_n827), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n870), .A2(new_n871), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n817), .A2(G87), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n840), .B2(new_n809), .ZN(new_n877));
  XOR2_X1   g0677(.A(new_n877), .B(KEYINPUT103), .Z(new_n878));
  INV_X1    g0678(.A(G294), .ZN(new_n879));
  OAI221_X1 g0679(.A(new_n245), .B1(new_n879), .B2(new_n805), .C1(new_n841), .C2(new_n555), .ZN(new_n880));
  INV_X1    g0680(.A(G303), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n825), .B1(new_n833), .B2(new_n844), .C1(new_n881), .C2(new_n830), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n880), .B(new_n882), .C1(G107), .C2(new_n827), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n875), .B1(new_n878), .B2(new_n883), .ZN(new_n884));
  OAI221_X1 g0684(.A(new_n866), .B1(new_n854), .B2(new_n781), .C1(new_n803), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n864), .A2(new_n885), .ZN(G384));
  OR2_X1    g0686(.A1(new_n512), .A2(KEYINPUT35), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n512), .A2(KEYINPUT35), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n887), .A2(new_n888), .A3(G116), .A4(new_n211), .ZN(new_n889));
  XOR2_X1   g0689(.A(new_n889), .B(KEYINPUT36), .Z(new_n890));
  OAI211_X1 g0690(.A(new_n208), .B(G77), .C1(new_n320), .C2(new_n280), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n400), .A2(G68), .ZN(new_n892));
  AOI211_X1 g0692(.A(new_n256), .B(G13), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT105), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT37), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n379), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n361), .B1(new_n347), .B2(new_n708), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n895), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n708), .B1(new_n332), .B2(new_n346), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n347), .B2(new_n359), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n901), .A2(KEYINPUT105), .A3(new_n896), .A4(new_n379), .ZN(new_n902));
  INV_X1    g0702(.A(new_n693), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT37), .B1(new_n898), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n899), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n694), .A2(new_n360), .A3(new_n363), .A4(new_n695), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n900), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT38), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT39), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT38), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n382), .B2(new_n900), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n905), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n909), .A2(new_n910), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n382), .A2(new_n900), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT38), .B1(new_n905), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n913), .A2(KEYINPUT106), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT106), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n912), .A2(new_n905), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n916), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n914), .B1(new_n920), .B2(new_n910), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n697), .A2(new_n710), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT104), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n852), .B1(new_n689), .B2(new_n859), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n310), .A2(new_n710), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n311), .A2(new_n926), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n310), .B(new_n710), .C1(new_n309), .C2(new_n297), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n924), .B1(new_n925), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n860), .B1(new_n751), .B2(new_n682), .ZN(new_n932));
  OAI211_X1 g0732(.A(KEYINPUT104), .B(new_n929), .C1(new_n932), .C2(new_n852), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n912), .A2(new_n905), .A3(new_n918), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n918), .B1(new_n912), .B2(new_n905), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n905), .A2(new_n915), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n934), .A2(new_n935), .B1(new_n936), .B2(KEYINPUT38), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n931), .A2(new_n933), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n696), .A2(new_n708), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n923), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n463), .A2(new_n468), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n702), .B1(new_n753), .B2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n940), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n756), .A2(new_n768), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n944), .A2(new_n929), .A3(new_n854), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT40), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n945), .A2(new_n946), .A3(new_n937), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n909), .A2(new_n913), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n946), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n469), .A2(new_n944), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n951), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n952), .A2(G330), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n943), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n256), .B2(new_n773), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n943), .A2(new_n954), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n894), .B1(new_n956), .B2(new_n957), .ZN(G367));
  INV_X1    g0758(.A(new_n770), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n536), .B1(new_n515), .B2(new_n721), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n667), .A2(new_n710), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n725), .A2(new_n962), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n963), .A2(KEYINPUT44), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n963), .A2(KEYINPUT44), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n725), .A2(new_n962), .ZN(new_n968));
  XOR2_X1   g0768(.A(KEYINPUT111), .B(KEYINPUT45), .Z(new_n969));
  XNOR2_X1  g0769(.A(new_n968), .B(new_n969), .ZN(new_n970));
  AND3_X1   g0770(.A1(new_n967), .A2(new_n719), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n719), .B1(new_n967), .B2(new_n970), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n718), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n724), .B1(new_n974), .B2(new_n722), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n772), .B(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n959), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n730), .B(KEYINPUT41), .Z(new_n978));
  OAI21_X1  g0778(.A(new_n774), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n962), .ZN(new_n980));
  INV_X1    g0780(.A(new_n724), .ZN(new_n981));
  NOR3_X1   g0781(.A1(new_n980), .A2(KEYINPUT42), .A3(new_n981), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n982), .A2(KEYINPUT109), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(KEYINPUT109), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n962), .A2(new_n724), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n983), .A2(new_n984), .B1(KEYINPUT42), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n535), .B1(new_n960), .B2(new_n609), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n987), .A2(KEYINPUT108), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(KEYINPUT108), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n988), .A2(new_n721), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n721), .B1(new_n550), .B2(new_n611), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n739), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n734), .A2(new_n991), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n986), .A2(new_n990), .B1(KEYINPUT43), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n719), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n996), .A2(KEYINPUT110), .A3(new_n962), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT107), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT110), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n719), .B2(new_n980), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n997), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n998), .B1(new_n997), .B2(new_n1000), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n995), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  NOR3_X1   g0805(.A1(new_n1002), .A2(new_n995), .A3(new_n1003), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n1005), .A2(new_n1006), .B1(KEYINPUT43), .B2(new_n994), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1006), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1008), .A2(new_n1009), .A3(new_n1004), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n979), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(KEYINPUT112), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT112), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1007), .A2(new_n1013), .A3(new_n979), .A4(new_n1010), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n992), .A2(new_n782), .A3(new_n993), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n229), .A2(new_n790), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n798), .B1(new_n204), .B2(new_n436), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n776), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n823), .A2(new_n280), .ZN(new_n1019));
  INV_X1    g0819(.A(G143), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n830), .A2(new_n1020), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n1019), .B(new_n1021), .C1(G159), .C2(new_n820), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n245), .B1(new_n810), .B2(G137), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n403), .B2(new_n805), .C1(new_n841), .C2(new_n400), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G77), .B2(new_n816), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n827), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1022), .B(new_n1025), .C1(new_n320), .C2(new_n1026), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT113), .Z(new_n1028));
  AOI22_X1  g0828(.A1(new_n814), .A2(G283), .B1(G317), .B2(new_n810), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1029), .B(new_n245), .C1(new_n881), .C2(new_n805), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G97), .B2(new_n816), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n879), .A2(new_n833), .B1(new_n830), .B2(new_n840), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(G107), .B2(new_n824), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT46), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n1026), .B2(new_n555), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n827), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1031), .A2(new_n1033), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1028), .A2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT47), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1018), .B1(new_n1039), .B2(new_n797), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n1012), .A2(new_n1014), .B1(new_n1015), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(G387));
  INV_X1    g0842(.A(new_n782), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n718), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n791), .B1(new_n226), .B2(G45), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n728), .B2(new_n785), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n334), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1047));
  OAI21_X1  g0847(.A(KEYINPUT50), .B1(new_n334), .B2(G50), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1048), .B(new_n264), .C1(new_n280), .C2(new_n285), .ZN(new_n1049));
  NOR3_X1   g0849(.A1(new_n728), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1046), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n503), .B2(new_n729), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n776), .B1(new_n1052), .B2(new_n799), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n245), .B1(new_n810), .B2(G150), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1054), .B1(new_n400), .B2(new_n805), .C1(new_n841), .C2(new_n280), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(G77), .B2(new_n827), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n817), .A2(G97), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n824), .A2(new_n551), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G159), .A2(new_n821), .B1(new_n820), .B2(new_n336), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n1026), .A2(new_n879), .B1(new_n844), .B2(new_n823), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n814), .A2(G303), .B1(new_n838), .B2(G317), .ZN(new_n1062));
  INV_X1    g0862(.A(G322), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1062), .B1(new_n840), .B2(new_n833), .C1(new_n1063), .C2(new_n830), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT114), .Z(new_n1065));
  INV_X1    g0865(.A(KEYINPUT48), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1061), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n1066), .B2(new_n1065), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT49), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n245), .B1(new_n809), .B2(new_n831), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n816), .B2(G116), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT115), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1060), .B1(new_n1070), .B2(new_n1074), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1044), .B(new_n1053), .C1(new_n1075), .C2(new_n797), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n976), .B2(new_n775), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n976), .A2(new_n770), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1078), .A2(KEYINPUT116), .A3(new_n730), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n770), .B2(new_n976), .ZN(new_n1080));
  AOI21_X1  g0880(.A(KEYINPUT116), .B1(new_n1078), .B2(new_n730), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1077), .B1(new_n1080), .B2(new_n1081), .ZN(G393));
  INV_X1    g0882(.A(new_n973), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n774), .B1(new_n1083), .B2(KEYINPUT117), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(KEYINPUT117), .B2(new_n1083), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n237), .A2(new_n790), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n798), .B1(new_n497), .B2(new_n204), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n776), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G317), .A2(new_n821), .B1(new_n838), .B2(G311), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT119), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT52), .Z(new_n1091));
  OAI22_X1  g0891(.A1(new_n833), .A2(new_n881), .B1(new_n823), .B2(new_n555), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n245), .B1(new_n1063), .B2(new_n809), .C1(new_n841), .C2(new_n879), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1092), .B(new_n1093), .C1(G283), .C2(new_n827), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1091), .A2(new_n818), .A3(new_n1094), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n1095), .A2(KEYINPUT120), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(G150), .A2(new_n821), .B1(new_n838), .B2(G159), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT51), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n1026), .A2(new_n280), .B1(new_n1020), .B2(new_n809), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1099), .A2(KEYINPUT118), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n390), .B1(new_n833), .B2(new_n400), .C1(new_n334), .C2(new_n841), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G77), .B2(new_n824), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1099), .A2(KEYINPUT118), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1101), .A2(new_n1103), .A3(new_n876), .A4(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1095), .A2(KEYINPUT120), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1096), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1088), .B1(new_n1107), .B2(new_n797), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n1043), .B2(new_n962), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1085), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n730), .B1(new_n1083), .B2(new_n1078), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n1078), .B2(new_n1083), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(G390));
  AND2_X1   g0914(.A1(new_n912), .A2(new_n905), .ZN(new_n1115));
  NOR3_X1   g0915(.A1(new_n1115), .A2(new_n908), .A3(KEYINPUT39), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(KEYINPUT39), .B2(new_n937), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n780), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n865), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1119), .A2(new_n336), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n245), .B1(new_n809), .B2(new_n879), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n503), .A2(new_n833), .B1(new_n830), .B2(new_n844), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n1121), .B(new_n1122), .C1(G97), .C2(new_n814), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n805), .A2(new_n555), .B1(new_n823), .B2(new_n285), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT122), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1123), .A2(new_n828), .A3(new_n871), .A4(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(G128), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n1127), .A2(new_n830), .B1(new_n833), .B2(new_n868), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(G159), .B2(new_n824), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n816), .A2(G50), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(KEYINPUT54), .B(G143), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n245), .B1(new_n814), .B2(new_n1132), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n838), .A2(G132), .B1(new_n810), .B2(G125), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1129), .A2(new_n1130), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n827), .A2(G150), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT53), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1126), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n777), .B(new_n1120), .C1(new_n1138), .C2(new_n797), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1118), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n922), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n710), .B1(new_n741), .B2(new_n746), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n853), .A2(new_n459), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n852), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1141), .B(new_n948), .C1(new_n1144), .C2(new_n930), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n851), .B1(new_n858), .B2(new_n860), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n922), .B1(new_n1146), .B2(new_n929), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1145), .B1(new_n921), .B2(new_n1147), .ZN(new_n1148));
  AND4_X1   g0948(.A1(G330), .A2(new_n944), .A3(new_n929), .A4(new_n854), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1141), .B1(new_n925), .B2(new_n930), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n937), .A2(KEYINPUT39), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1151), .A2(new_n1152), .A3(new_n914), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n769), .A2(new_n854), .A3(new_n929), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1153), .A2(new_n1145), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1150), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1140), .B1(new_n1156), .B2(new_n774), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n730), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n469), .A2(new_n769), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1160), .B(new_n702), .C1(new_n753), .C2(new_n941), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n929), .B1(new_n769), .B2(new_n854), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1146), .B1(new_n1149), .B2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n944), .A2(G330), .A3(new_n854), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n930), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1166), .A2(new_n1144), .A3(new_n1154), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1162), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1159), .B1(new_n1156), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1161), .B1(new_n1164), .B2(new_n1167), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1171), .A2(new_n1150), .A3(new_n1155), .ZN(new_n1172));
  AOI21_X1  g0972(.A(KEYINPUT121), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n1153), .A2(new_n1145), .A3(new_n1154), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1154), .B1(new_n1153), .B2(new_n1145), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1169), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  AND4_X1   g0976(.A1(KEYINPUT121), .A2(new_n1176), .A3(new_n1172), .A4(new_n730), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1158), .B1(new_n1173), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(KEYINPUT123), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1176), .A2(new_n1172), .A3(new_n730), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT121), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1170), .A2(KEYINPUT121), .A3(new_n1172), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT123), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1184), .A2(new_n1185), .A3(new_n1158), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1179), .A2(new_n1186), .ZN(G378));
  INV_X1    g0987(.A(new_n708), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n409), .A2(new_n1188), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n432), .B(new_n1189), .Z(new_n1190));
  XNOR2_X1  g0990(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1190), .B(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n939), .B1(new_n1117), .B2(new_n1141), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n931), .A2(new_n933), .A3(new_n937), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1192), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n950), .A2(new_n755), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1192), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n923), .A2(new_n938), .A3(new_n939), .A4(new_n1197), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n1195), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1196), .B1(new_n1195), .B2(new_n1198), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n775), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n776), .B1(new_n1119), .B2(G50), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n263), .B(new_n245), .C1(new_n809), .C2(new_n844), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n841), .A2(new_n436), .B1(new_n503), .B2(new_n805), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(G77), .C2(new_n827), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n830), .A2(new_n555), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1019), .B(new_n1206), .C1(G97), .C2(new_n820), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n816), .A2(G58), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1205), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT58), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n245), .A2(new_n263), .ZN(new_n1211));
  AOI21_X1  g1011(.A(G50), .B1(new_n554), .B2(new_n263), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1209), .A2(new_n1210), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n814), .A2(G137), .B1(new_n838), .B2(G128), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n821), .A2(G125), .B1(G150), .B2(new_n824), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n827), .A2(new_n1132), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n820), .A2(G132), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n816), .A2(G159), .ZN(new_n1221));
  AOI211_X1 g1021(.A(G33), .B(G41), .C1(new_n810), .C2(G124), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1213), .B1(new_n1210), .B2(new_n1209), .C1(new_n1219), .C2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1202), .B1(new_n1224), .B2(new_n797), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n1197), .B2(new_n781), .ZN(new_n1226));
  XOR2_X1   g1026(.A(new_n1226), .B(KEYINPUT124), .Z(new_n1227));
  NAND2_X1  g1027(.A1(new_n1201), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1172), .A2(new_n1162), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT57), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1159), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1229), .B(KEYINPUT57), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1228), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(G375));
  NAND2_X1  g1035(.A1(new_n930), .A2(new_n780), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n776), .B1(new_n1119), .B2(G68), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n872), .A2(new_n830), .B1(new_n833), .B2(new_n1131), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(G50), .B2(new_n824), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n827), .A2(G159), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n805), .A2(new_n868), .B1(new_n809), .B2(new_n1127), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n245), .B(new_n1241), .C1(G150), .C2(new_n814), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1239), .A2(new_n1208), .A3(new_n1240), .A4(new_n1242), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n841), .A2(new_n503), .B1(new_n809), .B2(new_n881), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n390), .B(new_n1244), .C1(G283), .C2(new_n838), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n1058), .B1(new_n833), .B2(new_n555), .C1(new_n879), .C2(new_n830), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1245), .B(new_n1247), .C1(new_n497), .C2(new_n1026), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n845), .A2(new_n285), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1243), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1237), .B1(new_n1250), .B2(new_n797), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1168), .A2(new_n775), .B1(new_n1236), .B2(new_n1251), .ZN(new_n1252));
  OR2_X1    g1052(.A1(new_n1171), .A2(new_n978), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1162), .A2(new_n1168), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1252), .B1(new_n1253), .B2(new_n1254), .ZN(G381));
  INV_X1    g1055(.A(G384), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1113), .A2(new_n1256), .ZN(new_n1257));
  NOR4_X1   g1057(.A1(new_n1257), .A2(G396), .A3(G393), .A4(G381), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1158), .A2(new_n1180), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1258), .A2(new_n1041), .A3(new_n1234), .A4(new_n1260), .ZN(G407));
  NAND2_X1  g1061(.A1(new_n709), .A2(G213), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1234), .A2(new_n1260), .A3(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(G407), .A2(G213), .A3(new_n1264), .ZN(G409));
  NAND2_X1  g1065(.A1(G387), .A2(new_n1113), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1041), .A2(G390), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  XOR2_X1   g1068(.A(G393), .B(G396), .Z(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1266), .A2(new_n1269), .A3(new_n1267), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1169), .A2(KEYINPUT60), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1159), .B1(new_n1274), .B2(new_n1254), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1275), .B1(new_n1254), .B2(new_n1274), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1276), .A2(G384), .A3(new_n1252), .ZN(new_n1277));
  AOI21_X1  g1077(.A(G384), .B1(new_n1276), .B2(new_n1252), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1263), .A2(G2897), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G2897), .B(new_n1263), .C1(new_n1277), .C2(new_n1278), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1201), .B(new_n1226), .C1(new_n1230), .C2(new_n978), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1260), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT125), .ZN(new_n1286));
  AOI211_X1 g1086(.A(KEYINPUT123), .B(new_n1157), .C1(new_n1182), .C2(new_n1183), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1185), .B1(new_n1184), .B2(new_n1158), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1234), .B(new_n1286), .C1(new_n1287), .C2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1286), .B1(G378), .B2(new_n1234), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1285), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1283), .B1(new_n1292), .B2(new_n1262), .ZN(new_n1293));
  OAI21_X1  g1093(.A(KEYINPUT127), .B1(new_n1293), .B2(KEYINPUT61), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT127), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT61), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1288), .A2(new_n1287), .ZN(new_n1297));
  OAI21_X1  g1097(.A(KEYINPUT125), .B1(new_n1297), .B2(G375), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1289), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1263), .B1(new_n1299), .B2(new_n1285), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1295), .B(new_n1296), .C1(new_n1300), .C2(new_n1283), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1292), .A2(new_n1262), .A3(new_n1279), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(KEYINPUT62), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1294), .A2(new_n1301), .A3(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT126), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1300), .A2(new_n1305), .A3(new_n1279), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1302), .A2(KEYINPUT126), .ZN(new_n1307));
  AOI21_X1  g1107(.A(KEYINPUT62), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1273), .B1(new_n1304), .B2(new_n1308), .ZN(new_n1309));
  NOR3_X1   g1109(.A1(new_n1273), .A2(KEYINPUT61), .A3(new_n1293), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT63), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1306), .A2(new_n1307), .A3(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1300), .A2(KEYINPUT63), .A3(new_n1279), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1310), .A2(new_n1312), .A3(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1309), .A2(new_n1314), .ZN(G405));
  OAI21_X1  g1115(.A(new_n1299), .B1(new_n1234), .B2(new_n1259), .ZN(new_n1316));
  OR2_X1    g1116(.A1(new_n1316), .A2(new_n1279), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1279), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  XNOR2_X1  g1119(.A(new_n1319), .B(new_n1273), .ZN(G402));
endmodule


