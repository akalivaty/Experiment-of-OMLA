

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(G651), .A2(n673), .ZN(n668) );
  NAND2_X1 U553 ( .A1(n708), .A2(n812), .ZN(n713) );
  AND2_X1 U554 ( .A1(n550), .A2(G2104), .ZN(n913) );
  AND2_X1 U555 ( .A1(n784), .A2(KEYINPUT64), .ZN(n528) );
  NOR2_X1 U556 ( .A1(n824), .A2(n522), .ZN(n546) );
  NOR2_X1 U557 ( .A1(n713), .A2(n967), .ZN(n710) );
  AND2_X1 U558 ( .A1(n785), .A2(n770), .ZN(n769) );
  NOR2_X1 U559 ( .A1(n534), .A2(KEYINPUT33), .ZN(n533) );
  NOR2_X1 U560 ( .A1(n773), .A2(n535), .ZN(n534) );
  XNOR2_X1 U561 ( .A(n768), .B(n767), .ZN(n784) );
  NAND2_X1 U562 ( .A1(n520), .A2(n546), .ZN(n544) );
  XNOR2_X1 U563 ( .A(n543), .B(KEYINPUT68), .ZN(n542) );
  NAND2_X1 U564 ( .A1(n914), .A2(G137), .ZN(n543) );
  XNOR2_X1 U565 ( .A(n537), .B(n536), .ZN(n720) );
  INV_X1 U566 ( .A(KEYINPUT67), .ZN(n536) );
  NOR2_X1 U567 ( .A1(n711), .A2(n987), .ZN(n538) );
  INV_X1 U568 ( .A(n713), .ZN(n734) );
  XNOR2_X1 U569 ( .A(n525), .B(KEYINPUT31), .ZN(n760) );
  OR2_X1 U570 ( .A1(n744), .A2(n745), .ZN(n525) );
  NOR2_X1 U571 ( .A1(G1966), .A2(n791), .ZN(n764) );
  AND2_X1 U572 ( .A1(n531), .A2(n529), .ZN(n774) );
  NAND2_X1 U573 ( .A1(n530), .A2(n523), .ZN(n529) );
  AND2_X1 U574 ( .A1(n532), .A2(n533), .ZN(n531) );
  NAND2_X1 U575 ( .A1(G8), .A2(n713), .ZN(n791) );
  NOR2_X1 U576 ( .A1(n673), .A2(n567), .ZN(n662) );
  NOR2_X1 U577 ( .A1(G2104), .A2(G2105), .ZN(n548) );
  NOR2_X1 U578 ( .A1(G651), .A2(G543), .ZN(n659) );
  AND2_X1 U579 ( .A1(G2104), .A2(G2105), .ZN(n917) );
  NAND2_X1 U580 ( .A1(n545), .A2(n519), .ZN(n841) );
  NOR2_X1 U581 ( .A1(n541), .A2(n540), .ZN(G160) );
  XNOR2_X2 U582 ( .A(KEYINPUT70), .B(n564), .ZN(n604) );
  AND2_X1 U583 ( .A1(n554), .A2(G40), .ZN(n518) );
  AND2_X1 U584 ( .A1(n544), .A2(n840), .ZN(n519) );
  NAND2_X1 U585 ( .A1(n793), .A2(n792), .ZN(n520) );
  AND2_X1 U586 ( .A1(n760), .A2(n752), .ZN(n521) );
  NOR2_X2 U587 ( .A1(G2104), .A2(n550), .ZN(n627) );
  AND2_X1 U588 ( .A1(n994), .A2(n838), .ZN(n522) );
  AND2_X1 U589 ( .A1(n773), .A2(n535), .ZN(n523) );
  XNOR2_X1 U590 ( .A(KEYINPUT29), .B(KEYINPUT96), .ZN(n524) );
  INV_X1 U591 ( .A(KEYINPUT64), .ZN(n535) );
  NAND2_X1 U592 ( .A1(n761), .A2(n521), .ZN(n756) );
  NAND2_X1 U593 ( .A1(n526), .A2(n738), .ZN(n761) );
  XNOR2_X1 U594 ( .A(n527), .B(n524), .ZN(n526) );
  NAND2_X1 U595 ( .A1(n733), .A2(n732), .ZN(n527) );
  NAND2_X1 U596 ( .A1(n769), .A2(n528), .ZN(n532) );
  NAND2_X1 U597 ( .A1(n769), .A2(n784), .ZN(n530) );
  INV_X1 U598 ( .A(n720), .ZN(n712) );
  NAND2_X1 U599 ( .A1(n539), .A2(n538), .ZN(n537) );
  XNOR2_X1 U600 ( .A(n710), .B(n709), .ZN(n539) );
  INV_X1 U601 ( .A(n542), .ZN(n540) );
  INV_X1 U602 ( .A(n554), .ZN(n541) );
  NAND2_X1 U603 ( .A1(n518), .A2(n542), .ZN(n811) );
  NAND2_X1 U604 ( .A1(n794), .A2(n546), .ZN(n545) );
  AND2_X1 U605 ( .A1(n552), .A2(n551), .ZN(n547) );
  INV_X1 U606 ( .A(KEYINPUT95), .ZN(n718) );
  XNOR2_X1 U607 ( .A(n719), .B(n718), .ZN(n728) );
  INV_X1 U608 ( .A(KEYINPUT98), .ZN(n767) );
  INV_X1 U609 ( .A(KEYINPUT13), .ZN(n589) );
  NAND2_X1 U610 ( .A1(n596), .A2(n595), .ZN(n987) );
  AND2_X1 U611 ( .A1(n553), .A2(n547), .ZN(n554) );
  XOR2_X2 U612 ( .A(KEYINPUT17), .B(n548), .Z(n914) );
  INV_X1 U613 ( .A(G2105), .ZN(n550) );
  NAND2_X1 U614 ( .A1(G101), .A2(n913), .ZN(n549) );
  XOR2_X1 U615 ( .A(KEYINPUT23), .B(n549), .Z(n553) );
  NAND2_X1 U616 ( .A1(G125), .A2(n627), .ZN(n552) );
  NAND2_X1 U617 ( .A1(G113), .A2(n917), .ZN(n551) );
  AND2_X1 U618 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U619 ( .A1(G102), .A2(n913), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n555), .B(KEYINPUT88), .ZN(n558) );
  NAND2_X1 U621 ( .A1(G126), .A2(n627), .ZN(n556) );
  XOR2_X1 U622 ( .A(KEYINPUT87), .B(n556), .Z(n557) );
  NAND2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U624 ( .A1(n914), .A2(G138), .ZN(n560) );
  NAND2_X1 U625 ( .A1(n917), .A2(G114), .ZN(n559) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U627 ( .A1(n562), .A2(n561), .ZN(G164) );
  INV_X1 U628 ( .A(G57), .ZN(G237) );
  INV_X1 U629 ( .A(G132), .ZN(G219) );
  INV_X1 U630 ( .A(G82), .ZN(G220) );
  XOR2_X1 U631 ( .A(KEYINPUT0), .B(G543), .Z(n673) );
  NAND2_X1 U632 ( .A1(n668), .A2(G53), .ZN(n566) );
  INV_X1 U633 ( .A(G651), .ZN(n567) );
  NOR2_X1 U634 ( .A1(G543), .A2(n567), .ZN(n563) );
  XOR2_X1 U635 ( .A(KEYINPUT1), .B(n563), .Z(n564) );
  NAND2_X1 U636 ( .A1(G65), .A2(n604), .ZN(n565) );
  NAND2_X1 U637 ( .A1(n566), .A2(n565), .ZN(n571) );
  NAND2_X1 U638 ( .A1(G78), .A2(n662), .ZN(n569) );
  NAND2_X1 U639 ( .A1(G91), .A2(n659), .ZN(n568) );
  NAND2_X1 U640 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U641 ( .A1(n571), .A2(n570), .ZN(n988) );
  INV_X1 U642 ( .A(n988), .ZN(G299) );
  NAND2_X1 U643 ( .A1(n659), .A2(G89), .ZN(n572) );
  XNOR2_X1 U644 ( .A(n572), .B(KEYINPUT4), .ZN(n574) );
  NAND2_X1 U645 ( .A1(G76), .A2(n662), .ZN(n573) );
  NAND2_X1 U646 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U647 ( .A(n575), .B(KEYINPUT5), .ZN(n581) );
  NAND2_X1 U648 ( .A1(G63), .A2(n604), .ZN(n576) );
  XNOR2_X1 U649 ( .A(n576), .B(KEYINPUT76), .ZN(n578) );
  NAND2_X1 U650 ( .A1(G51), .A2(n668), .ZN(n577) );
  NAND2_X1 U651 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U652 ( .A(KEYINPUT6), .B(n579), .Z(n580) );
  NAND2_X1 U653 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U654 ( .A(n582), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U655 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U656 ( .A1(G7), .A2(G661), .ZN(n583) );
  XOR2_X1 U657 ( .A(n583), .B(KEYINPUT10), .Z(n842) );
  NAND2_X1 U658 ( .A1(n842), .A2(G567), .ZN(n584) );
  XOR2_X1 U659 ( .A(KEYINPUT11), .B(n584), .Z(G234) );
  NAND2_X1 U660 ( .A1(G68), .A2(n662), .ZN(n588) );
  NAND2_X1 U661 ( .A1(G81), .A2(n659), .ZN(n585) );
  XNOR2_X1 U662 ( .A(n585), .B(KEYINPUT72), .ZN(n586) );
  XNOR2_X1 U663 ( .A(n586), .B(KEYINPUT12), .ZN(n587) );
  NAND2_X1 U664 ( .A1(n588), .A2(n587), .ZN(n590) );
  XNOR2_X1 U665 ( .A(n590), .B(n589), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n604), .A2(G56), .ZN(n591) );
  XNOR2_X1 U667 ( .A(n591), .B(KEYINPUT14), .ZN(n592) );
  XNOR2_X1 U668 ( .A(n592), .B(KEYINPUT71), .ZN(n593) );
  NOR2_X1 U669 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U670 ( .A1(n668), .A2(G43), .ZN(n595) );
  INV_X1 U671 ( .A(G860), .ZN(n620) );
  OR2_X1 U672 ( .A1(n987), .A2(n620), .ZN(G153) );
  NAND2_X1 U673 ( .A1(n668), .A2(G52), .ZN(n598) );
  NAND2_X1 U674 ( .A1(G64), .A2(n604), .ZN(n597) );
  NAND2_X1 U675 ( .A1(n598), .A2(n597), .ZN(n603) );
  NAND2_X1 U676 ( .A1(G77), .A2(n662), .ZN(n600) );
  NAND2_X1 U677 ( .A1(G90), .A2(n659), .ZN(n599) );
  NAND2_X1 U678 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U679 ( .A(KEYINPUT9), .B(n601), .Z(n602) );
  NOR2_X1 U680 ( .A1(n603), .A2(n602), .ZN(G171) );
  INV_X1 U681 ( .A(G171), .ZN(G301) );
  NAND2_X1 U682 ( .A1(G868), .A2(G301), .ZN(n616) );
  NAND2_X1 U683 ( .A1(G92), .A2(n659), .ZN(n606) );
  NAND2_X1 U684 ( .A1(G66), .A2(n604), .ZN(n605) );
  NAND2_X1 U685 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U686 ( .A(n607), .B(KEYINPUT73), .ZN(n609) );
  NAND2_X1 U687 ( .A1(G79), .A2(n662), .ZN(n608) );
  NAND2_X1 U688 ( .A1(n609), .A2(n608), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n668), .A2(G54), .ZN(n610) );
  XOR2_X1 U690 ( .A(KEYINPUT74), .B(n610), .Z(n611) );
  NOR2_X1 U691 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U692 ( .A(n613), .B(KEYINPUT15), .ZN(n614) );
  XOR2_X1 U693 ( .A(n614), .B(KEYINPUT75), .Z(n986) );
  INV_X1 U694 ( .A(G868), .ZN(n687) );
  NAND2_X1 U695 ( .A1(n986), .A2(n687), .ZN(n615) );
  NAND2_X1 U696 ( .A1(n616), .A2(n615), .ZN(G284) );
  XOR2_X1 U697 ( .A(KEYINPUT77), .B(n687), .Z(n617) );
  NOR2_X1 U698 ( .A1(G286), .A2(n617), .ZN(n619) );
  NOR2_X1 U699 ( .A1(G868), .A2(G299), .ZN(n618) );
  NOR2_X1 U700 ( .A1(n619), .A2(n618), .ZN(G297) );
  NAND2_X1 U701 ( .A1(n620), .A2(G559), .ZN(n621) );
  INV_X1 U702 ( .A(n986), .ZN(n926) );
  NAND2_X1 U703 ( .A1(n621), .A2(n926), .ZN(n622) );
  XNOR2_X1 U704 ( .A(n622), .B(KEYINPUT16), .ZN(n623) );
  XNOR2_X1 U705 ( .A(KEYINPUT78), .B(n623), .ZN(G148) );
  NOR2_X1 U706 ( .A1(G868), .A2(n987), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n926), .A2(G868), .ZN(n624) );
  NOR2_X1 U708 ( .A1(G559), .A2(n624), .ZN(n625) );
  NOR2_X1 U709 ( .A1(n626), .A2(n625), .ZN(G282) );
  NAND2_X1 U710 ( .A1(G123), .A2(n627), .ZN(n628) );
  XNOR2_X1 U711 ( .A(n628), .B(KEYINPUT18), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n913), .A2(G99), .ZN(n629) );
  NAND2_X1 U713 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U714 ( .A1(G135), .A2(n914), .ZN(n632) );
  NAND2_X1 U715 ( .A1(G111), .A2(n917), .ZN(n631) );
  NAND2_X1 U716 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U717 ( .A1(n634), .A2(n633), .ZN(n942) );
  XNOR2_X1 U718 ( .A(n942), .B(G2096), .ZN(n635) );
  INV_X1 U719 ( .A(G2100), .ZN(n864) );
  NAND2_X1 U720 ( .A1(n635), .A2(n864), .ZN(G156) );
  NAND2_X1 U721 ( .A1(n662), .A2(G80), .ZN(n636) );
  XNOR2_X1 U722 ( .A(n636), .B(KEYINPUT80), .ZN(n638) );
  NAND2_X1 U723 ( .A1(G93), .A2(n659), .ZN(n637) );
  NAND2_X1 U724 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U725 ( .A1(n668), .A2(G55), .ZN(n640) );
  NAND2_X1 U726 ( .A1(G67), .A2(n604), .ZN(n639) );
  NAND2_X1 U727 ( .A1(n640), .A2(n639), .ZN(n641) );
  OR2_X1 U728 ( .A1(n642), .A2(n641), .ZN(n688) );
  NAND2_X1 U729 ( .A1(G559), .A2(n926), .ZN(n643) );
  XOR2_X1 U730 ( .A(n987), .B(n643), .Z(n684) );
  XNOR2_X1 U731 ( .A(KEYINPUT79), .B(n684), .ZN(n644) );
  NOR2_X1 U732 ( .A1(G860), .A2(n644), .ZN(n645) );
  XOR2_X1 U733 ( .A(n688), .B(n645), .Z(G145) );
  NAND2_X1 U734 ( .A1(G75), .A2(n662), .ZN(n647) );
  NAND2_X1 U735 ( .A1(G88), .A2(n659), .ZN(n646) );
  NAND2_X1 U736 ( .A1(n647), .A2(n646), .ZN(n651) );
  NAND2_X1 U737 ( .A1(n668), .A2(G50), .ZN(n649) );
  NAND2_X1 U738 ( .A1(G62), .A2(n604), .ZN(n648) );
  NAND2_X1 U739 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U740 ( .A1(n651), .A2(n650), .ZN(G166) );
  INV_X1 U741 ( .A(G166), .ZN(G303) );
  NAND2_X1 U742 ( .A1(G85), .A2(n659), .ZN(n653) );
  NAND2_X1 U743 ( .A1(G60), .A2(n604), .ZN(n652) );
  NAND2_X1 U744 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U745 ( .A1(G72), .A2(n662), .ZN(n654) );
  XNOR2_X1 U746 ( .A(KEYINPUT69), .B(n654), .ZN(n655) );
  NOR2_X1 U747 ( .A1(n656), .A2(n655), .ZN(n658) );
  NAND2_X1 U748 ( .A1(n668), .A2(G47), .ZN(n657) );
  NAND2_X1 U749 ( .A1(n658), .A2(n657), .ZN(G290) );
  NAND2_X1 U750 ( .A1(G86), .A2(n659), .ZN(n661) );
  NAND2_X1 U751 ( .A1(G61), .A2(n604), .ZN(n660) );
  NAND2_X1 U752 ( .A1(n661), .A2(n660), .ZN(n665) );
  NAND2_X1 U753 ( .A1(n662), .A2(G73), .ZN(n663) );
  XOR2_X1 U754 ( .A(KEYINPUT2), .B(n663), .Z(n664) );
  NOR2_X1 U755 ( .A1(n665), .A2(n664), .ZN(n667) );
  NAND2_X1 U756 ( .A1(n668), .A2(G48), .ZN(n666) );
  NAND2_X1 U757 ( .A1(n667), .A2(n666), .ZN(G305) );
  NAND2_X1 U758 ( .A1(G49), .A2(n668), .ZN(n669) );
  XNOR2_X1 U759 ( .A(n669), .B(KEYINPUT81), .ZN(n672) );
  NAND2_X1 U760 ( .A1(G74), .A2(G651), .ZN(n670) );
  XOR2_X1 U761 ( .A(KEYINPUT82), .B(n670), .Z(n671) );
  NOR2_X1 U762 ( .A1(n672), .A2(n671), .ZN(n677) );
  NAND2_X1 U763 ( .A1(G87), .A2(n673), .ZN(n674) );
  XNOR2_X1 U764 ( .A(KEYINPUT83), .B(n674), .ZN(n675) );
  NOR2_X1 U765 ( .A1(n604), .A2(n675), .ZN(n676) );
  NAND2_X1 U766 ( .A1(n677), .A2(n676), .ZN(G288) );
  XOR2_X1 U767 ( .A(n688), .B(G290), .Z(n678) );
  XNOR2_X1 U768 ( .A(n678), .B(G305), .ZN(n679) );
  XOR2_X1 U769 ( .A(n679), .B(KEYINPUT84), .Z(n681) );
  XOR2_X1 U770 ( .A(G299), .B(KEYINPUT19), .Z(n680) );
  XNOR2_X1 U771 ( .A(n681), .B(n680), .ZN(n682) );
  XOR2_X1 U772 ( .A(G303), .B(n682), .Z(n683) );
  XNOR2_X1 U773 ( .A(n683), .B(G288), .ZN(n929) );
  XOR2_X1 U774 ( .A(n684), .B(n929), .Z(n685) );
  XNOR2_X1 U775 ( .A(KEYINPUT85), .B(n685), .ZN(n686) );
  NOR2_X1 U776 ( .A1(n687), .A2(n686), .ZN(n690) );
  NOR2_X1 U777 ( .A1(G868), .A2(n688), .ZN(n689) );
  NOR2_X1 U778 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U779 ( .A(KEYINPUT86), .B(n691), .ZN(G295) );
  NAND2_X1 U780 ( .A1(G2078), .A2(G2084), .ZN(n692) );
  XOR2_X1 U781 ( .A(KEYINPUT20), .B(n692), .Z(n693) );
  NAND2_X1 U782 ( .A1(G2090), .A2(n693), .ZN(n694) );
  XNOR2_X1 U783 ( .A(KEYINPUT21), .B(n694), .ZN(n695) );
  NAND2_X1 U784 ( .A1(n695), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U785 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U786 ( .A1(G220), .A2(G219), .ZN(n696) );
  XOR2_X1 U787 ( .A(KEYINPUT22), .B(n696), .Z(n697) );
  NOR2_X1 U788 ( .A1(G218), .A2(n697), .ZN(n698) );
  NAND2_X1 U789 ( .A1(G96), .A2(n698), .ZN(n848) );
  NAND2_X1 U790 ( .A1(n848), .A2(G2106), .ZN(n702) );
  NAND2_X1 U791 ( .A1(G69), .A2(G120), .ZN(n699) );
  NOR2_X1 U792 ( .A1(G237), .A2(n699), .ZN(n700) );
  NAND2_X1 U793 ( .A1(G108), .A2(n700), .ZN(n847) );
  NAND2_X1 U794 ( .A1(n847), .A2(G567), .ZN(n701) );
  NAND2_X1 U795 ( .A1(n702), .A2(n701), .ZN(n863) );
  NAND2_X1 U796 ( .A1(G483), .A2(G661), .ZN(n703) );
  NOR2_X1 U797 ( .A1(n863), .A2(n703), .ZN(n845) );
  NAND2_X1 U798 ( .A1(n845), .A2(G36), .ZN(G176) );
  INV_X1 U799 ( .A(KEYINPUT92), .ZN(n704) );
  XNOR2_X1 U800 ( .A(n704), .B(n811), .ZN(n708) );
  NOR2_X1 U801 ( .A1(G164), .A2(G1384), .ZN(n707) );
  INV_X1 U802 ( .A(KEYINPUT65), .ZN(n706) );
  XNOR2_X1 U803 ( .A(n707), .B(n706), .ZN(n812) );
  XOR2_X1 U804 ( .A(G1996), .B(KEYINPUT94), .Z(n967) );
  XOR2_X1 U805 ( .A(KEYINPUT66), .B(KEYINPUT26), .Z(n709) );
  AND2_X1 U806 ( .A1(n713), .A2(G1341), .ZN(n711) );
  NAND2_X1 U807 ( .A1(n712), .A2(n926), .ZN(n717) );
  NOR2_X1 U808 ( .A1(n734), .A2(G1348), .ZN(n715) );
  NOR2_X1 U809 ( .A1(G2067), .A2(n713), .ZN(n714) );
  NOR2_X1 U810 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U811 ( .A1(n717), .A2(n716), .ZN(n719) );
  NAND2_X1 U812 ( .A1(n986), .A2(n720), .ZN(n726) );
  NAND2_X1 U813 ( .A1(n734), .A2(G2072), .ZN(n721) );
  XNOR2_X1 U814 ( .A(n721), .B(KEYINPUT27), .ZN(n723) );
  AND2_X1 U815 ( .A1(G1956), .A2(n713), .ZN(n722) );
  NOR2_X1 U816 ( .A1(n723), .A2(n722), .ZN(n729) );
  NOR2_X1 U817 ( .A1(n988), .A2(n729), .ZN(n724) );
  XNOR2_X1 U818 ( .A(n724), .B(KEYINPUT28), .ZN(n731) );
  INV_X1 U819 ( .A(n731), .ZN(n725) );
  AND2_X1 U820 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U821 ( .A1(n728), .A2(n727), .ZN(n733) );
  NAND2_X1 U822 ( .A1(n988), .A2(n729), .ZN(n730) );
  OR2_X1 U823 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U824 ( .A1(n734), .A2(G1961), .ZN(n735) );
  XOR2_X1 U825 ( .A(KEYINPUT93), .B(n735), .Z(n737) );
  XOR2_X1 U826 ( .A(KEYINPUT25), .B(G2078), .Z(n968) );
  NOR2_X1 U827 ( .A1(n713), .A2(n968), .ZN(n736) );
  NOR2_X1 U828 ( .A1(n737), .A2(n736), .ZN(n739) );
  OR2_X1 U829 ( .A1(n739), .A2(G301), .ZN(n738) );
  NAND2_X1 U830 ( .A1(n739), .A2(G301), .ZN(n740) );
  XNOR2_X1 U831 ( .A(n740), .B(KEYINPUT97), .ZN(n745) );
  NOR2_X1 U832 ( .A1(G2084), .A2(n713), .ZN(n762) );
  NOR2_X1 U833 ( .A1(n764), .A2(n762), .ZN(n741) );
  NAND2_X1 U834 ( .A1(G8), .A2(n741), .ZN(n742) );
  XNOR2_X1 U835 ( .A(KEYINPUT30), .B(n742), .ZN(n743) );
  NOR2_X1 U836 ( .A1(n743), .A2(G168), .ZN(n744) );
  INV_X1 U837 ( .A(G8), .ZN(n751) );
  NOR2_X1 U838 ( .A1(G1971), .A2(n791), .ZN(n747) );
  NOR2_X1 U839 ( .A1(G2090), .A2(n713), .ZN(n746) );
  NOR2_X1 U840 ( .A1(n747), .A2(n746), .ZN(n748) );
  XOR2_X1 U841 ( .A(KEYINPUT99), .B(n748), .Z(n749) );
  NAND2_X1 U842 ( .A1(n749), .A2(G303), .ZN(n750) );
  OR2_X1 U843 ( .A1(n751), .A2(n750), .ZN(n752) );
  INV_X1 U844 ( .A(n752), .ZN(n754) );
  AND2_X1 U845 ( .A1(G286), .A2(G8), .ZN(n753) );
  OR2_X1 U846 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U847 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U848 ( .A(KEYINPUT32), .B(n757), .ZN(n785) );
  INV_X1 U849 ( .A(n791), .ZN(n759) );
  NAND2_X1 U850 ( .A1(G288), .A2(G1976), .ZN(n758) );
  XNOR2_X1 U851 ( .A(n758), .B(KEYINPUT100), .ZN(n996) );
  AND2_X1 U852 ( .A1(n759), .A2(n996), .ZN(n770) );
  NAND2_X1 U853 ( .A1(n761), .A2(n760), .ZN(n766) );
  AND2_X1 U854 ( .A1(G8), .A2(n762), .ZN(n763) );
  NOR2_X1 U855 ( .A1(n764), .A2(n763), .ZN(n765) );
  AND2_X1 U856 ( .A1(n766), .A2(n765), .ZN(n768) );
  INV_X1 U857 ( .A(n770), .ZN(n772) );
  NOR2_X1 U858 ( .A1(G1976), .A2(G288), .ZN(n775) );
  NOR2_X1 U859 ( .A1(G1971), .A2(G303), .ZN(n771) );
  NOR2_X1 U860 ( .A1(n775), .A2(n771), .ZN(n995) );
  OR2_X1 U861 ( .A1(n772), .A2(n995), .ZN(n773) );
  XNOR2_X1 U862 ( .A(n774), .B(KEYINPUT101), .ZN(n779) );
  XOR2_X1 U863 ( .A(G1981), .B(G305), .Z(n1002) );
  NAND2_X1 U864 ( .A1(n775), .A2(KEYINPUT33), .ZN(n776) );
  OR2_X1 U865 ( .A1(n791), .A2(n776), .ZN(n777) );
  AND2_X1 U866 ( .A1(n1002), .A2(n777), .ZN(n778) );
  NAND2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n781) );
  INV_X1 U868 ( .A(KEYINPUT102), .ZN(n780) );
  XNOR2_X1 U869 ( .A(n781), .B(n780), .ZN(n794) );
  NOR2_X1 U870 ( .A1(G2090), .A2(G303), .ZN(n782) );
  XOR2_X1 U871 ( .A(KEYINPUT103), .B(n782), .Z(n783) );
  NAND2_X1 U872 ( .A1(G8), .A2(n783), .ZN(n787) );
  NAND2_X1 U873 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U874 ( .A1(n787), .A2(n786), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n788), .A2(n791), .ZN(n793) );
  NOR2_X1 U876 ( .A1(G1981), .A2(G305), .ZN(n789) );
  XOR2_X1 U877 ( .A(n789), .B(KEYINPUT24), .Z(n790) );
  OR2_X1 U878 ( .A1(n791), .A2(n790), .ZN(n792) );
  NAND2_X1 U879 ( .A1(G95), .A2(n913), .ZN(n796) );
  NAND2_X1 U880 ( .A1(G131), .A2(n914), .ZN(n795) );
  NAND2_X1 U881 ( .A1(n796), .A2(n795), .ZN(n800) );
  NAND2_X1 U882 ( .A1(G119), .A2(n627), .ZN(n798) );
  NAND2_X1 U883 ( .A1(G107), .A2(n917), .ZN(n797) );
  NAND2_X1 U884 ( .A1(n798), .A2(n797), .ZN(n799) );
  NOR2_X1 U885 ( .A1(n800), .A2(n799), .ZN(n905) );
  INV_X1 U886 ( .A(G1991), .ZN(n877) );
  NOR2_X1 U887 ( .A1(n905), .A2(n877), .ZN(n810) );
  NAND2_X1 U888 ( .A1(G105), .A2(n913), .ZN(n801) );
  XOR2_X1 U889 ( .A(KEYINPUT91), .B(n801), .Z(n802) );
  XNOR2_X1 U890 ( .A(n802), .B(KEYINPUT38), .ZN(n804) );
  NAND2_X1 U891 ( .A1(G129), .A2(n627), .ZN(n803) );
  NAND2_X1 U892 ( .A1(n804), .A2(n803), .ZN(n808) );
  NAND2_X1 U893 ( .A1(G141), .A2(n914), .ZN(n806) );
  NAND2_X1 U894 ( .A1(G117), .A2(n917), .ZN(n805) );
  NAND2_X1 U895 ( .A1(n806), .A2(n805), .ZN(n807) );
  OR2_X1 U896 ( .A1(n808), .A2(n807), .ZN(n901) );
  AND2_X1 U897 ( .A1(n901), .A2(G1996), .ZN(n809) );
  NOR2_X1 U898 ( .A1(n810), .A2(n809), .ZN(n945) );
  INV_X1 U899 ( .A(n945), .ZN(n813) );
  NOR2_X1 U900 ( .A1(n812), .A2(n811), .ZN(n838) );
  NAND2_X1 U901 ( .A1(n813), .A2(n838), .ZN(n827) );
  NAND2_X1 U902 ( .A1(G104), .A2(n913), .ZN(n815) );
  NAND2_X1 U903 ( .A1(G140), .A2(n914), .ZN(n814) );
  NAND2_X1 U904 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U905 ( .A(KEYINPUT34), .B(n816), .ZN(n821) );
  NAND2_X1 U906 ( .A1(G128), .A2(n627), .ZN(n818) );
  NAND2_X1 U907 ( .A1(G116), .A2(n917), .ZN(n817) );
  NAND2_X1 U908 ( .A1(n818), .A2(n817), .ZN(n819) );
  XOR2_X1 U909 ( .A(n819), .B(KEYINPUT35), .Z(n820) );
  NOR2_X1 U910 ( .A1(n821), .A2(n820), .ZN(n822) );
  XOR2_X1 U911 ( .A(KEYINPUT36), .B(n822), .Z(n823) );
  XOR2_X1 U912 ( .A(KEYINPUT90), .B(n823), .Z(n910) );
  XNOR2_X1 U913 ( .A(G2067), .B(KEYINPUT37), .ZN(n826) );
  NOR2_X1 U914 ( .A1(n910), .A2(n826), .ZN(n959) );
  NAND2_X1 U915 ( .A1(n838), .A2(n959), .ZN(n836) );
  NAND2_X1 U916 ( .A1(n827), .A2(n836), .ZN(n824) );
  XOR2_X1 U917 ( .A(G1986), .B(KEYINPUT89), .Z(n825) );
  XNOR2_X1 U918 ( .A(G290), .B(n825), .ZN(n994) );
  NAND2_X1 U919 ( .A1(n910), .A2(n826), .ZN(n948) );
  INV_X1 U920 ( .A(n827), .ZN(n831) );
  NOR2_X1 U921 ( .A1(G1986), .A2(G290), .ZN(n828) );
  AND2_X1 U922 ( .A1(n877), .A2(n905), .ZN(n943) );
  NOR2_X1 U923 ( .A1(n828), .A2(n943), .ZN(n829) );
  XNOR2_X1 U924 ( .A(n829), .B(KEYINPUT104), .ZN(n830) );
  NOR2_X1 U925 ( .A1(n831), .A2(n830), .ZN(n832) );
  NOR2_X1 U926 ( .A1(G1996), .A2(n901), .ZN(n940) );
  NOR2_X1 U927 ( .A1(n832), .A2(n940), .ZN(n834) );
  XOR2_X1 U928 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n833) );
  XNOR2_X1 U929 ( .A(n834), .B(n833), .ZN(n835) );
  NAND2_X1 U930 ( .A1(n836), .A2(n835), .ZN(n837) );
  NAND2_X1 U931 ( .A1(n948), .A2(n837), .ZN(n839) );
  NAND2_X1 U932 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U933 ( .A(n841), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n842), .ZN(G217) );
  INV_X1 U935 ( .A(n842), .ZN(G223) );
  AND2_X1 U936 ( .A1(G15), .A2(G2), .ZN(n843) );
  NAND2_X1 U937 ( .A1(G661), .A2(n843), .ZN(G259) );
  NAND2_X1 U938 ( .A1(G3), .A2(G1), .ZN(n844) );
  XNOR2_X1 U939 ( .A(KEYINPUT110), .B(n844), .ZN(n846) );
  NAND2_X1 U940 ( .A1(n846), .A2(n845), .ZN(G188) );
  INV_X1 U942 ( .A(G120), .ZN(G236) );
  INV_X1 U943 ( .A(G96), .ZN(G221) );
  INV_X1 U944 ( .A(G69), .ZN(G235) );
  NOR2_X1 U945 ( .A1(n848), .A2(n847), .ZN(n849) );
  XOR2_X1 U946 ( .A(n849), .B(KEYINPUT111), .Z(G325) );
  INV_X1 U947 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U948 ( .A(G1341), .B(G1348), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n850), .B(G2427), .ZN(n860) );
  XOR2_X1 U950 ( .A(G2438), .B(G2446), .Z(n852) );
  XNOR2_X1 U951 ( .A(G2451), .B(KEYINPUT107), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U953 ( .A(G2443), .B(KEYINPUT106), .Z(n854) );
  XNOR2_X1 U954 ( .A(G2430), .B(G2454), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U956 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U957 ( .A(KEYINPUT108), .B(G2435), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(n861) );
  NAND2_X1 U960 ( .A1(n861), .A2(G14), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n862), .B(KEYINPUT109), .ZN(G401) );
  INV_X1 U962 ( .A(n863), .ZN(G319) );
  XNOR2_X1 U963 ( .A(n864), .B(G2096), .ZN(n866) );
  XNOR2_X1 U964 ( .A(KEYINPUT42), .B(G2678), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n866), .B(n865), .ZN(n870) );
  XOR2_X1 U966 ( .A(KEYINPUT43), .B(G2090), .Z(n868) );
  XNOR2_X1 U967 ( .A(G2067), .B(G2072), .ZN(n867) );
  XNOR2_X1 U968 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U969 ( .A(n870), .B(n869), .Z(n872) );
  XNOR2_X1 U970 ( .A(G2078), .B(G2084), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(G227) );
  XOR2_X1 U972 ( .A(G1981), .B(G1961), .Z(n874) );
  XNOR2_X1 U973 ( .A(G1986), .B(G1966), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n874), .B(n873), .ZN(n885) );
  XOR2_X1 U975 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n876) );
  XNOR2_X1 U976 ( .A(G1996), .B(KEYINPUT41), .ZN(n875) );
  XNOR2_X1 U977 ( .A(n876), .B(n875), .ZN(n881) );
  XOR2_X1 U978 ( .A(G1976), .B(G1971), .Z(n879) );
  XOR2_X1 U979 ( .A(n877), .B(G1956), .Z(n878) );
  XNOR2_X1 U980 ( .A(n879), .B(n878), .ZN(n880) );
  XOR2_X1 U981 ( .A(n881), .B(n880), .Z(n883) );
  XNOR2_X1 U982 ( .A(KEYINPUT114), .B(G2474), .ZN(n882) );
  XNOR2_X1 U983 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U984 ( .A(n885), .B(n884), .ZN(G229) );
  NAND2_X1 U985 ( .A1(G124), .A2(n627), .ZN(n886) );
  XNOR2_X1 U986 ( .A(n886), .B(KEYINPUT44), .ZN(n888) );
  NAND2_X1 U987 ( .A1(n913), .A2(G100), .ZN(n887) );
  NAND2_X1 U988 ( .A1(n888), .A2(n887), .ZN(n892) );
  NAND2_X1 U989 ( .A1(G136), .A2(n914), .ZN(n890) );
  NAND2_X1 U990 ( .A1(G112), .A2(n917), .ZN(n889) );
  NAND2_X1 U991 ( .A1(n890), .A2(n889), .ZN(n891) );
  NOR2_X1 U992 ( .A1(n892), .A2(n891), .ZN(G162) );
  NAND2_X1 U993 ( .A1(G130), .A2(n627), .ZN(n894) );
  NAND2_X1 U994 ( .A1(G118), .A2(n917), .ZN(n893) );
  NAND2_X1 U995 ( .A1(n894), .A2(n893), .ZN(n900) );
  NAND2_X1 U996 ( .A1(n913), .A2(G106), .ZN(n895) );
  XOR2_X1 U997 ( .A(KEYINPUT115), .B(n895), .Z(n897) );
  NAND2_X1 U998 ( .A1(n914), .A2(G142), .ZN(n896) );
  NAND2_X1 U999 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U1000 ( .A(n898), .B(KEYINPUT45), .Z(n899) );
  NOR2_X1 U1001 ( .A1(n900), .A2(n899), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n902), .B(n901), .ZN(n909) );
  XNOR2_X1 U1003 ( .A(KEYINPUT48), .B(KEYINPUT116), .ZN(n903) );
  XNOR2_X1 U1004 ( .A(n903), .B(KEYINPUT46), .ZN(n904) );
  XOR2_X1 U1005 ( .A(n904), .B(n942), .Z(n907) );
  XNOR2_X1 U1006 ( .A(G164), .B(n905), .ZN(n906) );
  XNOR2_X1 U1007 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1008 ( .A(n909), .B(n908), .Z(n912) );
  XNOR2_X1 U1009 ( .A(n910), .B(G162), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(n912), .B(n911), .ZN(n924) );
  NAND2_X1 U1011 ( .A1(G103), .A2(n913), .ZN(n916) );
  NAND2_X1 U1012 ( .A1(G139), .A2(n914), .ZN(n915) );
  NAND2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(n922) );
  NAND2_X1 U1014 ( .A1(G127), .A2(n627), .ZN(n919) );
  NAND2_X1 U1015 ( .A1(G115), .A2(n917), .ZN(n918) );
  NAND2_X1 U1016 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1017 ( .A(KEYINPUT47), .B(n920), .Z(n921) );
  NOR2_X1 U1018 ( .A1(n922), .A2(n921), .ZN(n950) );
  XOR2_X1 U1019 ( .A(n950), .B(G160), .Z(n923) );
  XNOR2_X1 U1020 ( .A(n924), .B(n923), .ZN(n925) );
  NOR2_X1 U1021 ( .A1(G37), .A2(n925), .ZN(G395) );
  XNOR2_X1 U1022 ( .A(n987), .B(KEYINPUT117), .ZN(n928) );
  XOR2_X1 U1023 ( .A(G301), .B(n926), .Z(n927) );
  XNOR2_X1 U1024 ( .A(n928), .B(n927), .ZN(n931) );
  XOR2_X1 U1025 ( .A(n929), .B(G286), .Z(n930) );
  XNOR2_X1 U1026 ( .A(n931), .B(n930), .ZN(n932) );
  NOR2_X1 U1027 ( .A1(G37), .A2(n932), .ZN(G397) );
  NOR2_X1 U1028 ( .A1(G227), .A2(G229), .ZN(n933) );
  XOR2_X1 U1029 ( .A(KEYINPUT49), .B(n933), .Z(n934) );
  NAND2_X1 U1030 ( .A1(G319), .A2(n934), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(G401), .A2(n935), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(KEYINPUT118), .B(n936), .ZN(n938) );
  NOR2_X1 U1033 ( .A1(G395), .A2(G397), .ZN(n937) );
  NAND2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(G225) );
  INV_X1 U1035 ( .A(G225), .ZN(G308) );
  INV_X1 U1036 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1037 ( .A(G2090), .B(G162), .Z(n939) );
  NOR2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1039 ( .A(KEYINPUT51), .B(n941), .Z(n957) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n947) );
  XOR2_X1 U1042 ( .A(G160), .B(G2084), .Z(n946) );
  NOR2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n949) );
  NAND2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n955) );
  XOR2_X1 U1045 ( .A(G2072), .B(n950), .Z(n952) );
  XOR2_X1 U1046 ( .A(G164), .B(G2078), .Z(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1048 ( .A(KEYINPUT50), .B(n953), .Z(n954) );
  NOR2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1052 ( .A(KEYINPUT52), .B(n960), .ZN(n962) );
  INV_X1 U1053 ( .A(KEYINPUT55), .ZN(n961) );
  NAND2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1055 ( .A1(n963), .A2(G29), .ZN(n1044) );
  XNOR2_X1 U1056 ( .A(G2090), .B(G35), .ZN(n978) );
  XOR2_X1 U1057 ( .A(G25), .B(G1991), .Z(n964) );
  NAND2_X1 U1058 ( .A1(n964), .A2(G28), .ZN(n974) );
  XNOR2_X1 U1059 ( .A(G2067), .B(G26), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(G33), .B(G2072), .ZN(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n972) );
  XOR2_X1 U1062 ( .A(n967), .B(G32), .Z(n970) );
  XNOR2_X1 U1063 ( .A(G27), .B(n968), .ZN(n969) );
  NOR2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1067 ( .A(KEYINPUT119), .B(n975), .Z(n976) );
  XNOR2_X1 U1068 ( .A(n976), .B(KEYINPUT53), .ZN(n977) );
  NOR2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n981) );
  XOR2_X1 U1070 ( .A(G2084), .B(G34), .Z(n979) );
  XNOR2_X1 U1071 ( .A(KEYINPUT54), .B(n979), .ZN(n980) );
  NAND2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1073 ( .A(KEYINPUT55), .B(n982), .Z(n984) );
  INV_X1 U1074 ( .A(G29), .ZN(n983) );
  NAND2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1076 ( .A1(G11), .A2(n985), .ZN(n1042) );
  XNOR2_X1 U1077 ( .A(G16), .B(KEYINPUT56), .ZN(n1012) );
  XOR2_X1 U1078 ( .A(n986), .B(G1348), .Z(n1010) );
  XOR2_X1 U1079 ( .A(G301), .B(G1961), .Z(n992) );
  XNOR2_X1 U1080 ( .A(n987), .B(G1341), .ZN(n990) );
  XOR2_X1 U1081 ( .A(n988), .B(G1956), .Z(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n1001) );
  AND2_X1 U1085 ( .A1(G303), .A2(G1971), .ZN(n998) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1088 ( .A(n999), .B(KEYINPUT122), .ZN(n1000) );
  NAND2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1008) );
  XNOR2_X1 U1090 ( .A(G1966), .B(G168), .ZN(n1003) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(n1004), .B(KEYINPUT57), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(n1006), .B(n1005), .ZN(n1007) );
  NOR2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1040) );
  XNOR2_X1 U1098 ( .A(KEYINPUT59), .B(G1348), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(n1013), .B(G4), .ZN(n1020) );
  XNOR2_X1 U1100 ( .A(G1956), .B(G20), .ZN(n1018) );
  XNOR2_X1 U1101 ( .A(G1341), .B(G19), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(G6), .B(G1981), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1104 ( .A(KEYINPUT125), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1107 ( .A(KEYINPUT60), .B(n1021), .ZN(n1024) );
  XNOR2_X1 U1108 ( .A(KEYINPUT124), .B(G1961), .ZN(n1022) );
  XNOR2_X1 U1109 ( .A(G5), .B(n1022), .ZN(n1023) );
  NOR2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1027) );
  XOR2_X1 U1111 ( .A(G1966), .B(KEYINPUT126), .Z(n1025) );
  XNOR2_X1 U1112 ( .A(G21), .B(n1025), .ZN(n1026) );
  NAND2_X1 U1113 ( .A1(n1027), .A2(n1026), .ZN(n1035) );
  XNOR2_X1 U1114 ( .A(KEYINPUT127), .B(KEYINPUT58), .ZN(n1033) );
  XOR2_X1 U1115 ( .A(G1986), .B(G24), .Z(n1031) );
  XNOR2_X1 U1116 ( .A(G1971), .B(G22), .ZN(n1029) );
  XNOR2_X1 U1117 ( .A(G23), .B(G1976), .ZN(n1028) );
  NOR2_X1 U1118 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1119 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1120 ( .A(n1033), .B(n1032), .Z(n1034) );
  NOR2_X1 U1121 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1122 ( .A(n1036), .B(KEYINPUT61), .ZN(n1038) );
  XNOR2_X1 U1123 ( .A(G16), .B(KEYINPUT123), .ZN(n1037) );
  NAND2_X1 U1124 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NAND2_X1 U1125 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  NOR2_X1 U1126 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  NAND2_X1 U1127 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  XNOR2_X1 U1128 ( .A(KEYINPUT62), .B(n1045), .ZN(G150) );
  INV_X1 U1129 ( .A(G150), .ZN(G311) );
endmodule

