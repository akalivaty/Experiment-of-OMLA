//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 0 1 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n801,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  OAI22_X1  g003(.A1(KEYINPUT66), .A2(new_n188), .B1(new_n189), .B2(G137), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(KEYINPUT66), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G131), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT67), .ZN(new_n194));
  INV_X1    g008(.A(G137), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G134), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n189), .A2(KEYINPUT67), .A3(G137), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(G134), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(KEYINPUT66), .A3(new_n188), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n192), .A2(new_n193), .A3(new_n198), .A4(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT68), .ZN(new_n202));
  INV_X1    g016(.A(new_n191), .ZN(new_n203));
  AOI22_X1  g017(.A1(new_n203), .A2(new_n199), .B1(new_n196), .B2(new_n197), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT68), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n204), .A2(new_n205), .A3(new_n192), .A4(new_n193), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G143), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n210), .B1(new_n211), .B2(G146), .ZN(new_n212));
  NOR3_X1   g026(.A1(new_n208), .A2(KEYINPUT64), .A3(G143), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n209), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G128), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n215), .B1(new_n209), .B2(KEYINPUT1), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n211), .A2(G146), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n209), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT70), .B1(new_n195), .B2(G134), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n223), .B1(new_n189), .B2(G137), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT70), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n224), .B1(new_n225), .B2(new_n199), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G131), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n207), .A2(new_n222), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n193), .B1(new_n204), .B2(new_n192), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n229), .B1(new_n202), .B2(new_n206), .ZN(new_n230));
  AND2_X1   g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  NOR2_X1   g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n209), .A2(new_n220), .A3(new_n231), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT65), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n209), .A2(new_n220), .A3(new_n231), .A4(new_n236), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n214), .A2(new_n233), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n228), .B(KEYINPUT30), .C1(new_n230), .C2(new_n239), .ZN(new_n240));
  XOR2_X1   g054(.A(KEYINPUT2), .B(G113), .Z(new_n241));
  XNOR2_X1  g055(.A(G116), .B(G119), .ZN(new_n242));
  OR2_X1    g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n242), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n229), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n207), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT69), .B1(new_n248), .B2(new_n238), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n250));
  NOR3_X1   g064(.A1(new_n230), .A2(new_n250), .A3(new_n239), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n202), .A2(new_n206), .B1(G131), .B2(new_n226), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n222), .B1(new_n252), .B2(KEYINPUT71), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n207), .A2(KEYINPUT71), .A3(new_n227), .ZN(new_n254));
  OAI22_X1  g068(.A1(new_n249), .A2(new_n251), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT30), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n246), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AOI22_X1  g071(.A1(new_n248), .A2(new_n238), .B1(new_n252), .B2(new_n222), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n245), .B(KEYINPUT72), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  XOR2_X1   g074(.A(KEYINPUT73), .B(KEYINPUT27), .Z(new_n261));
  NOR2_X1   g075(.A1(G237), .A2(G953), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G210), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n261), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT26), .B(G101), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  NOR3_X1   g081(.A1(new_n257), .A2(KEYINPUT74), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT74), .ZN(new_n269));
  INV_X1    g083(.A(new_n245), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n270), .B1(new_n258), .B2(KEYINPUT30), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n252), .A2(KEYINPUT71), .ZN(new_n272));
  INV_X1    g086(.A(new_n222), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n207), .A2(new_n227), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT71), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n248), .A2(KEYINPUT69), .A3(new_n238), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n250), .B1(new_n230), .B2(new_n239), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n272), .A2(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n271), .B1(new_n279), .B2(KEYINPUT30), .ZN(new_n280));
  INV_X1    g094(.A(new_n267), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n269), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT31), .B1(new_n268), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT31), .B1(new_n280), .B2(new_n281), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n266), .ZN(new_n287));
  XNOR2_X1  g101(.A(KEYINPUT75), .B(KEYINPUT28), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n228), .B1(new_n230), .B2(new_n239), .ZN(new_n289));
  INV_X1    g103(.A(new_n259), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n274), .A2(new_n275), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n292), .A2(new_n222), .A3(new_n272), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n277), .A2(new_n278), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n270), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n291), .B1(new_n295), .B2(KEYINPUT76), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT76), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n297), .B1(new_n279), .B2(new_n270), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n288), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT77), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n290), .B1(new_n289), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n258), .A2(KEYINPUT77), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT28), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n287), .B1(new_n299), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT78), .B1(new_n286), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT74), .B1(new_n257), .B2(new_n267), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n280), .A2(new_n269), .A3(new_n281), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n284), .B1(new_n308), .B2(KEYINPUT31), .ZN(new_n309));
  INV_X1    g123(.A(new_n288), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n255), .A2(KEYINPUT76), .A3(new_n245), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n260), .ZN(new_n312));
  AOI21_X1  g126(.A(KEYINPUT76), .B1(new_n255), .B2(new_n245), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n310), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n303), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n266), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT78), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n309), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n187), .B1(new_n305), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT32), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT80), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT29), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n280), .A2(new_n260), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n287), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n315), .A2(new_n266), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n323), .B(new_n325), .C1(new_n299), .C2(new_n326), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n303), .A2(new_n323), .A3(new_n287), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n289), .A2(new_n290), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n260), .A2(new_n329), .A3(KEYINPUT79), .ZN(new_n330));
  OR3_X1    g144(.A1(new_n258), .A2(KEYINPUT79), .A3(new_n259), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n331), .A3(KEYINPUT28), .ZN(new_n332));
  AOI21_X1  g146(.A(G902), .B1(new_n328), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n327), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n322), .B1(new_n334), .B2(G472), .ZN(new_n335));
  INV_X1    g149(.A(G472), .ZN(new_n336));
  AOI211_X1 g150(.A(KEYINPUT80), .B(new_n336), .C1(new_n327), .C2(new_n333), .ZN(new_n337));
  OR2_X1    g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n187), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n317), .B1(new_n309), .B2(new_n316), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT31), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n341), .B1(new_n306), .B2(new_n307), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n304), .B(KEYINPUT78), .C1(new_n342), .C2(new_n284), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n339), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT32), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n321), .A2(new_n338), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n215), .A2(G119), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT82), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT23), .ZN(new_n350));
  INV_X1    g164(.A(G119), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n350), .B1(new_n351), .B2(G128), .ZN(new_n352));
  NOR2_X1   g166(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n353));
  OAI22_X1  g167(.A1(new_n349), .A2(new_n352), .B1(new_n347), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(G119), .B(G128), .ZN(new_n355));
  XOR2_X1   g169(.A(KEYINPUT24), .B(G110), .Z(new_n356));
  OAI22_X1  g170(.A1(new_n354), .A2(G110), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT16), .ZN(new_n358));
  INV_X1    g172(.A(G140), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n359), .A3(G125), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(G125), .ZN(new_n361));
  INV_X1    g175(.A(G125), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G140), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(G146), .B(new_n360), .C1(new_n364), .C2(new_n358), .ZN(new_n365));
  INV_X1    g179(.A(new_n364), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n208), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n357), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n360), .B1(new_n364), .B2(new_n358), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n208), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n370), .A2(new_n365), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n354), .A2(G110), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n356), .A2(new_n355), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n371), .A2(KEYINPUT83), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT83), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n372), .A2(new_n373), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n370), .A2(new_n365), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n368), .B1(new_n375), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G953), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(G221), .A3(G234), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(KEYINPUT84), .ZN(new_n383));
  XNOR2_X1  g197(.A(KEYINPUT22), .B(G137), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n383), .B(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G902), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT83), .B1(new_n371), .B2(new_n374), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n377), .A2(new_n376), .A3(new_n378), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(new_n368), .A3(new_n385), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n387), .A2(new_n388), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT85), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT25), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(KEYINPUT85), .A3(KEYINPUT25), .ZN(new_n397));
  XOR2_X1   g211(.A(KEYINPUT81), .B(G217), .Z(new_n398));
  AOI21_X1  g212(.A(new_n398), .B1(G234), .B2(new_n388), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n396), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n387), .A2(new_n392), .ZN(new_n401));
  NOR3_X1   g215(.A1(new_n401), .A2(G902), .A3(new_n399), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n400), .A2(KEYINPUT86), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(KEYINPUT86), .B1(new_n400), .B2(new_n403), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT9), .B(G234), .ZN(new_n407));
  OAI21_X1  g221(.A(G221), .B1(new_n407), .B2(G902), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  XOR2_X1   g223(.A(G110), .B(G140), .Z(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(KEYINPUT87), .ZN(new_n411));
  INV_X1    g225(.A(G227), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(G953), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n411), .B(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(G104), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT3), .B1(new_n415), .B2(G107), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT3), .ZN(new_n417));
  INV_X1    g231(.A(G107), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n418), .A3(G104), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n415), .A2(G107), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n416), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT88), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT88), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n416), .A2(new_n419), .A3(new_n423), .A4(new_n420), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n422), .A2(G101), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(G101), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n416), .A2(new_n419), .A3(new_n426), .A4(new_n420), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n427), .A2(KEYINPUT4), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT4), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n422), .A2(new_n430), .A3(G101), .A4(new_n424), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n429), .A2(new_n238), .A3(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n415), .A2(G107), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n418), .A2(G104), .ZN(new_n434));
  OAI21_X1  g248(.A(G101), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n427), .A2(new_n435), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n209), .A2(new_n220), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n221), .B1(new_n437), .B2(new_n216), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT10), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n222), .A2(KEYINPUT10), .A3(new_n436), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n432), .A2(new_n230), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT89), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n442), .A2(new_n441), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT89), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n445), .A2(new_n432), .A3(new_n446), .A4(new_n230), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n414), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT12), .ZN(new_n449));
  OR2_X1    g263(.A1(new_n449), .A2(KEYINPUT90), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(KEYINPUT90), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n439), .B1(new_n222), .B2(new_n436), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n450), .B(new_n451), .C1(new_n453), .C2(new_n230), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n248), .A2(KEYINPUT90), .A3(new_n449), .A4(new_n452), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n448), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n414), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n444), .A2(new_n447), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n445), .A2(new_n432), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n248), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n458), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  NOR3_X1   g277(.A1(new_n463), .A2(G469), .A3(G902), .ZN(new_n464));
  INV_X1    g278(.A(G469), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n458), .B1(new_n456), .B2(new_n459), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n448), .A2(KEYINPUT91), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n461), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n448), .A2(KEYINPUT91), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n467), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n465), .B1(new_n471), .B2(new_n388), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT92), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n464), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n470), .ZN(new_n475));
  AOI22_X1  g289(.A1(new_n448), .A2(KEYINPUT91), .B1(new_n248), .B2(new_n460), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n466), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n477), .A2(G902), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT92), .B1(new_n478), .B2(new_n465), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n409), .B1(new_n474), .B2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(G113), .B(G122), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(new_n415), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n262), .A2(G214), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT98), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n483), .B1(new_n484), .B2(new_n211), .ZN(new_n485));
  AND2_X1   g299(.A1(KEYINPUT98), .A2(G143), .ZN(new_n486));
  NOR2_X1   g300(.A1(KEYINPUT98), .A2(G143), .ZN(new_n487));
  OAI211_X1 g301(.A(G214), .B(new_n262), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(G131), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n485), .A2(new_n488), .A3(new_n193), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(KEYINPUT99), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT99), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n485), .A2(new_n493), .A3(new_n488), .A4(new_n193), .ZN(new_n494));
  NOR2_X1   g308(.A1(KEYINPUT100), .A2(KEYINPUT19), .ZN(new_n495));
  AND2_X1   g309(.A1(KEYINPUT100), .A2(KEYINPUT19), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n364), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n497), .B(new_n208), .C1(new_n364), .C2(new_n496), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n492), .A2(new_n365), .A3(new_n494), .A4(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT18), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n485), .B(new_n488), .C1(new_n500), .C2(new_n193), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n364), .B(G146), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n501), .B(new_n502), .C1(new_n490), .C2(new_n500), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n482), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n503), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT17), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n485), .A2(new_n488), .A3(new_n193), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n193), .B1(new_n485), .B2(new_n488), .ZN(new_n508));
  NOR3_X1   g322(.A1(new_n507), .A2(new_n508), .A3(new_n493), .ZN(new_n509));
  INV_X1    g323(.A(new_n494), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n378), .B1(KEYINPUT17), .B2(new_n508), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n505), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n504), .B1(new_n513), .B2(new_n482), .ZN(new_n514));
  NOR2_X1   g328(.A1(G475), .A2(G902), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT20), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n499), .A2(new_n503), .ZN(new_n518));
  INV_X1    g332(.A(new_n482), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT17), .B1(new_n492), .B2(new_n494), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n371), .B1(new_n506), .B2(new_n490), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n482), .B(new_n503), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT20), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n525), .A3(new_n515), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n517), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n503), .B1(new_n521), .B2(new_n522), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n519), .ZN(new_n529));
  AND2_X1   g343(.A1(new_n529), .A2(new_n523), .ZN(new_n530));
  OAI21_X1  g344(.A(G475), .B1(new_n530), .B2(G902), .ZN(new_n531));
  INV_X1    g345(.A(G116), .ZN(new_n532));
  OAI21_X1  g346(.A(KEYINPUT101), .B1(new_n532), .B2(G122), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT101), .ZN(new_n534));
  INV_X1    g348(.A(G122), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n535), .A3(G116), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n532), .A2(G122), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(G107), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n537), .A2(new_n418), .A3(new_n538), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT102), .ZN(new_n543));
  OAI22_X1  g357(.A1(new_n543), .A2(KEYINPUT13), .B1(new_n211), .B2(G128), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT13), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(KEYINPUT102), .ZN(new_n546));
  OAI21_X1  g360(.A(G134), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(G128), .B(G143), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n548), .B(G134), .C1(new_n544), .C2(new_n546), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n542), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n538), .A2(KEYINPUT14), .ZN(new_n554));
  OR3_X1    g368(.A1(new_n535), .A2(KEYINPUT14), .A3(G116), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n537), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G107), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n548), .B(new_n189), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n557), .A2(new_n558), .A3(new_n541), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n398), .A2(G953), .A3(new_n407), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n553), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT103), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n553), .A2(new_n559), .ZN(new_n564));
  INV_X1    g378(.A(new_n560), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n553), .A2(new_n559), .A3(KEYINPUT103), .A4(new_n560), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n563), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT15), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(G478), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n568), .A2(new_n388), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n570), .B1(new_n568), .B2(new_n388), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(G952), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(G953), .ZN(new_n575));
  INV_X1    g389(.A(G234), .ZN(new_n576));
  INV_X1    g390(.A(G237), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  AOI211_X1 g393(.A(new_n388), .B(new_n381), .C1(G234), .C2(G237), .ZN(new_n580));
  XNOR2_X1  g394(.A(KEYINPUT21), .B(G898), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n527), .A2(new_n531), .A3(new_n573), .A4(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(KEYINPUT104), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT97), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n429), .A2(new_n245), .A3(new_n431), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n242), .A2(KEYINPUT5), .ZN(new_n588));
  INV_X1    g402(.A(G113), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n532), .A2(G119), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT5), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n588), .A2(new_n592), .B1(new_n241), .B2(new_n242), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n436), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n587), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(G110), .B(G122), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT93), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n587), .A2(new_n598), .A3(new_n594), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(KEYINPUT6), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n214), .A2(new_n233), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n235), .A2(new_n237), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n362), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n211), .A2(G146), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n210), .A2(new_n211), .A3(G146), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n362), .B(new_n221), .C1(new_n609), .C2(new_n216), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n605), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(G224), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(G953), .ZN(new_n614));
  XOR2_X1   g428(.A(new_n612), .B(new_n614), .Z(new_n615));
  INV_X1    g429(.A(KEYINPUT6), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n595), .A2(new_n616), .A3(new_n599), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n602), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT95), .ZN(new_n619));
  OAI22_X1  g433(.A1(new_n605), .A2(new_n611), .B1(new_n619), .B2(new_n614), .ZN(new_n620));
  OAI21_X1  g434(.A(KEYINPUT7), .B1(new_n613), .B2(G953), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n598), .B(KEYINPUT8), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n593), .A2(new_n436), .A3(KEYINPUT94), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n351), .A2(G116), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n590), .A2(new_n626), .A3(new_n591), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n590), .A2(new_n591), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(G113), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n244), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n427), .A2(new_n435), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n625), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(KEYINPUT94), .B1(new_n593), .B2(new_n436), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n624), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI221_X1 g449(.A(new_n621), .B1(new_n619), .B2(new_n614), .C1(new_n605), .C2(new_n611), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n623), .A2(new_n601), .A3(new_n635), .A4(new_n636), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n637), .A2(new_n388), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n618), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(G210), .B1(G237), .B2(G902), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT96), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n618), .A2(new_n638), .A3(new_n640), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n618), .A2(new_n638), .A3(new_n640), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT96), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g462(.A(G214), .B1(G237), .B2(G902), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n586), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n645), .A2(KEYINPUT97), .A3(new_n649), .A4(new_n647), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n585), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n480), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n346), .A2(new_n406), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G101), .ZN(G3));
  OAI21_X1  g470(.A(new_n388), .B1(new_n305), .B2(new_n318), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(G472), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n473), .B(G469), .C1(new_n477), .C2(G902), .ZN(new_n659));
  OR2_X1    g473(.A1(new_n457), .A2(new_n462), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n660), .A2(new_n465), .A3(new_n388), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n472), .A2(new_n473), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n406), .B(new_n408), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n658), .A2(new_n665), .A3(new_n319), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n640), .B1(new_n618), .B2(new_n638), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n649), .B1(new_n646), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT105), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT105), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n671), .B(new_n649), .C1(new_n646), .C2(new_n668), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n553), .A2(new_n559), .ZN(new_n675));
  OR3_X1    g489(.A1(new_n675), .A2(KEYINPUT106), .A3(new_n560), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n560), .B1(new_n675), .B2(KEYINPUT106), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n676), .A2(KEYINPUT33), .A3(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT33), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n568), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n388), .A2(G478), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n568), .A2(new_n388), .ZN(new_n683));
  OAI22_X1  g497(.A1(new_n681), .A2(new_n682), .B1(G478), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n525), .B1(new_n524), .B2(new_n515), .ZN(new_n685));
  AOI211_X1 g499(.A(KEYINPUT20), .B(new_n516), .C1(new_n520), .C2(new_n523), .ZN(new_n686));
  INV_X1    g500(.A(G475), .ZN(new_n687));
  AOI21_X1  g501(.A(G902), .B1(new_n529), .B2(new_n523), .ZN(new_n688));
  OAI22_X1  g502(.A1(new_n685), .A2(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n684), .A2(new_n689), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n674), .A2(new_n583), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n667), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT34), .B(G104), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G6));
  NOR4_X1   g508(.A1(new_n673), .A2(new_n582), .A3(new_n573), .A4(new_n689), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n667), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT35), .B(G107), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G9));
  NOR2_X1   g512(.A1(new_n386), .A2(KEYINPUT36), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n380), .B(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n399), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(new_n388), .A3(new_n701), .ZN(new_n702));
  OR2_X1    g516(.A1(new_n702), .A2(KEYINPUT107), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(KEYINPUT107), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(new_n400), .A3(new_n704), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n480), .A2(new_n653), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n344), .B1(new_n657), .B2(G472), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT37), .B(G110), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G12));
  AND2_X1   g524(.A1(new_n346), .A2(new_n480), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n670), .A2(new_n705), .A3(new_n672), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n689), .A2(new_n573), .ZN(new_n713));
  INV_X1    g527(.A(new_n580), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n578), .B1(new_n714), .B2(G900), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n711), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G128), .ZN(G30));
  XNOR2_X1  g533(.A(new_n715), .B(KEYINPUT39), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n480), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(KEYINPUT40), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n648), .B(KEYINPUT38), .ZN(new_n723));
  INV_X1    g537(.A(new_n705), .ZN(new_n724));
  INV_X1    g538(.A(new_n689), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n573), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n724), .A2(new_n649), .A3(new_n726), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n722), .A2(new_n723), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n721), .A2(KEYINPUT40), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n330), .A2(new_n331), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n308), .B1(new_n287), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(G472), .B1(new_n731), .B2(G902), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n321), .A2(new_n345), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n728), .A2(new_n729), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G143), .ZN(G45));
  NAND3_X1  g549(.A1(new_n684), .A2(new_n689), .A3(new_n715), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n712), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n711), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G146), .ZN(G48));
  INV_X1    g553(.A(new_n406), .ZN(new_n740));
  OAI21_X1  g554(.A(G469), .B1(new_n463), .B2(G902), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n661), .A2(new_n408), .A3(new_n741), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n346), .A2(new_n691), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT41), .B(G113), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(KEYINPUT108), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n744), .B(new_n746), .ZN(G15));
  NAND3_X1  g561(.A1(new_n346), .A2(new_n695), .A3(new_n743), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G116), .ZN(G18));
  NOR3_X1   g563(.A1(new_n712), .A2(new_n585), .A3(new_n742), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n346), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G119), .ZN(G21));
  NAND3_X1  g566(.A1(new_n670), .A2(new_n672), .A3(new_n726), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n670), .A2(KEYINPUT109), .A3(new_n672), .A4(new_n726), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n742), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n583), .A3(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n400), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n402), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n266), .B1(new_n315), .B2(new_n332), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n187), .B1(new_n309), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(G902), .B1(new_n340), .B2(new_n343), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n761), .B(new_n763), .C1(new_n764), .C2(new_n336), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n759), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G122), .ZN(G24));
  INV_X1    g581(.A(KEYINPUT110), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n736), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n684), .A2(new_n689), .A3(KEYINPUT110), .A4(new_n715), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n712), .A2(new_n771), .A3(new_n742), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n772), .B(new_n763), .C1(new_n336), .C2(new_n764), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT111), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n658), .A2(new_n775), .A3(new_n763), .A4(new_n772), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G125), .ZN(G27));
  NOR2_X1   g592(.A1(new_n344), .A2(KEYINPUT32), .ZN(new_n779));
  AOI211_X1 g593(.A(new_n320), .B(new_n339), .C1(new_n340), .C2(new_n343), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n335), .A2(new_n337), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n740), .ZN(new_n783));
  NAND2_X1  g597(.A1(G469), .A2(G902), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n661), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT112), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n466), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n475), .A2(new_n476), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(G469), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT113), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n787), .A2(new_n791), .A3(G469), .A4(new_n788), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n785), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n650), .B1(new_n645), .B2(new_n647), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n408), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n793), .A2(KEYINPUT42), .A3(new_n795), .A4(new_n771), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n793), .A2(new_n795), .A3(new_n771), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n346), .A2(new_n761), .A3(new_n797), .ZN(new_n798));
  AOI22_X1  g612(.A1(new_n783), .A2(new_n796), .B1(new_n798), .B2(KEYINPUT42), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G131), .ZN(G33));
  NOR3_X1   g614(.A1(new_n793), .A2(new_n795), .A3(new_n716), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n346), .A2(new_n406), .A3(new_n801), .ZN(new_n802));
  XOR2_X1   g616(.A(KEYINPUT114), .B(G134), .Z(new_n803));
  XNOR2_X1  g617(.A(new_n802), .B(new_n803), .ZN(G36));
  INV_X1    g618(.A(KEYINPUT44), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n725), .A2(new_n684), .ZN(new_n806));
  XOR2_X1   g620(.A(new_n806), .B(KEYINPUT43), .Z(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n705), .ZN(new_n808));
  OR3_X1    g622(.A1(new_n707), .A2(new_n805), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n787), .A2(KEYINPUT45), .A3(new_n788), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT45), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n471), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n810), .A2(G469), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT46), .B1(new_n813), .B2(new_n784), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n464), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(KEYINPUT46), .A3(new_n784), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n817), .A2(new_n408), .A3(new_n720), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n805), .B1(new_n707), .B2(new_n808), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n809), .A2(new_n818), .A3(new_n794), .A4(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G137), .ZN(G39));
  INV_X1    g635(.A(new_n794), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n406), .A2(new_n822), .A3(new_n736), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n817), .A2(KEYINPUT47), .A3(new_n408), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT47), .B1(new_n817), .B2(new_n408), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n782), .B(new_n823), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G140), .ZN(G42));
  NAND2_X1  g642(.A1(new_n661), .A2(new_n741), .ZN(new_n829));
  XOR2_X1   g643(.A(new_n829), .B(KEYINPUT115), .Z(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT49), .ZN(new_n831));
  INV_X1    g645(.A(new_n733), .ZN(new_n832));
  INV_X1    g646(.A(new_n761), .ZN(new_n833));
  NOR4_X1   g647(.A1(new_n833), .A2(new_n409), .A3(new_n650), .A4(new_n806), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n831), .A2(new_n832), .A3(new_n723), .A4(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n836));
  INV_X1    g650(.A(new_n793), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n724), .A2(new_n408), .A3(new_n715), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n757), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n774), .A2(new_n776), .B1(new_n733), .B2(new_n840), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n346), .B(new_n480), .C1(new_n717), .C2(new_n737), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n841), .A2(KEYINPUT52), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT52), .B1(new_n841), .B2(new_n842), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n655), .A2(new_n744), .A3(new_n748), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n725), .A2(new_n573), .A3(new_n715), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n847), .B(KEYINPUT116), .Z(new_n848));
  NOR3_X1   g662(.A1(new_n848), .A2(new_n724), .A3(new_n822), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n346), .A2(new_n480), .A3(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n797), .A2(new_n658), .A3(new_n705), .A4(new_n763), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n802), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n750), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n708), .B1(new_n782), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n651), .A2(new_n652), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n855), .B(new_n583), .C1(new_n690), .C2(new_n713), .ZN(new_n856));
  OAI22_X1  g670(.A1(new_n666), .A2(new_n856), .B1(new_n765), .B2(new_n759), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n799), .A2(new_n846), .A3(new_n852), .A4(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n836), .B1(new_n845), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n841), .A2(new_n842), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT52), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n841), .A2(KEYINPUT52), .A3(new_n842), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n799), .A2(new_n852), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n655), .A2(new_n744), .A3(new_n748), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n867), .A2(new_n854), .A3(new_n857), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n865), .A2(new_n866), .A3(KEYINPUT53), .A4(new_n868), .ZN(new_n869));
  XNOR2_X1  g683(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n860), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n860), .B2(new_n869), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g688(.A(KEYINPUT118), .B(KEYINPUT51), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n876), .B1(new_n825), .B2(new_n826), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT47), .ZN(new_n878));
  INV_X1    g692(.A(new_n816), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n879), .A2(new_n814), .A3(new_n464), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n878), .B1(new_n880), .B2(new_n409), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n881), .A2(new_n824), .A3(KEYINPUT119), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n830), .A2(new_n409), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n883), .B(KEYINPUT120), .Z(new_n884));
  NAND3_X1  g698(.A1(new_n877), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n807), .A2(new_n579), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n765), .A2(new_n822), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n765), .A2(new_n886), .ZN(new_n889));
  INV_X1    g703(.A(new_n723), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n650), .B1(new_n891), .B2(KEYINPUT50), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n889), .A2(new_n758), .A3(new_n893), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n891), .A2(KEYINPUT50), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n743), .A2(new_n579), .A3(new_n794), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n733), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n684), .A2(new_n689), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n658), .A2(new_n705), .A3(new_n763), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n886), .A2(new_n742), .A3(new_n822), .ZN(new_n903));
  AOI22_X1  g717(.A1(new_n899), .A2(new_n900), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n896), .A2(new_n897), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n875), .B1(new_n888), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n899), .A2(new_n690), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n889), .A2(new_n674), .A3(new_n758), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n907), .A2(new_n575), .A3(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n782), .A2(new_n833), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n903), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n911), .A2(KEYINPUT48), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(KEYINPUT48), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n909), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT51), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n881), .A2(new_n824), .A3(new_n883), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n915), .B1(new_n916), .B2(new_n887), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n917), .A2(new_n897), .A3(new_n896), .A4(new_n904), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n914), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n906), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT122), .B1(new_n874), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n860), .A2(new_n869), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT54), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n860), .A2(new_n869), .A3(new_n870), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n923), .A2(KEYINPUT122), .A3(new_n924), .A4(new_n920), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n574), .A2(new_n381), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n835), .B1(new_n921), .B2(new_n927), .ZN(G75));
  NAND2_X1  g742(.A1(new_n602), .A2(new_n617), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(new_n615), .Z(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT55), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n388), .B1(new_n860), .B2(new_n869), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(G210), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT56), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AOI211_X1 g750(.A(KEYINPUT56), .B(new_n931), .C1(new_n933), .C2(G210), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n381), .A2(G952), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(G51));
  XOR2_X1   g753(.A(new_n784), .B(KEYINPUT57), .Z(new_n940));
  AOI21_X1  g754(.A(new_n870), .B1(new_n860), .B2(new_n869), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n940), .B1(new_n871), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n660), .ZN(new_n943));
  INV_X1    g757(.A(new_n813), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n933), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n938), .B1(new_n943), .B2(new_n945), .ZN(G54));
  NAND2_X1  g760(.A1(KEYINPUT58), .A2(G475), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT123), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n933), .A2(new_n524), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n524), .B1(new_n933), .B2(new_n948), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n949), .A2(new_n950), .A3(new_n938), .ZN(G60));
  INV_X1    g765(.A(new_n681), .ZN(new_n952));
  NAND2_X1  g766(.A1(G478), .A2(G902), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT59), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n952), .B(new_n954), .C1(new_n871), .C2(new_n941), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n955), .B1(G952), .B2(new_n381), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n923), .A2(new_n924), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n952), .B1(new_n957), .B2(new_n954), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n956), .A2(new_n958), .ZN(G63));
  AND2_X1   g773(.A1(new_n860), .A2(new_n869), .ZN(new_n960));
  NAND2_X1  g774(.A1(G217), .A2(G902), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT60), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n401), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n962), .B1(new_n860), .B2(new_n869), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n938), .B1(new_n964), .B2(new_n700), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n964), .A2(new_n700), .ZN(new_n967));
  AOI21_X1  g781(.A(KEYINPUT61), .B1(new_n967), .B2(KEYINPUT124), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT124), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(new_n964), .B2(new_n700), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n963), .B(new_n965), .C1(new_n971), .C2(KEYINPUT61), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n969), .A2(new_n972), .ZN(G66));
  OAI21_X1  g787(.A(G953), .B1(new_n581), .B2(new_n613), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n868), .B2(G953), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n929), .B1(G898), .B2(new_n381), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(G69));
  NAND3_X1  g791(.A1(new_n910), .A2(new_n818), .A3(new_n757), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT125), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n842), .A2(new_n777), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n827), .A2(new_n820), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n799), .A2(new_n802), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT126), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n982), .A2(new_n381), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n240), .B1(new_n279), .B2(KEYINPUT30), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n496), .A2(new_n495), .ZN(new_n987));
  MUX2_X1   g801(.A(new_n496), .B(new_n987), .S(new_n364), .Z(new_n988));
  XOR2_X1   g802(.A(new_n986), .B(new_n988), .Z(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n990), .B1(G900), .B2(G953), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n985), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n827), .A2(new_n820), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n794), .B1(new_n690), .B2(new_n713), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n721), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n993), .B1(new_n783), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n980), .A2(new_n734), .ZN(new_n997));
  OR2_X1    g811(.A1(new_n997), .A2(KEYINPUT62), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(KEYINPUT62), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n996), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n381), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n992), .B1(new_n1002), .B2(new_n989), .ZN(new_n1003));
  INV_X1    g817(.A(G900), .ZN(new_n1004));
  OAI21_X1  g818(.A(G953), .B1(new_n412), .B2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT127), .Z(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  OAI211_X1 g822(.A(new_n992), .B(new_n1006), .C1(new_n1002), .C2(new_n989), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(G72));
  NAND3_X1  g824(.A1(new_n280), .A2(new_n287), .A3(new_n260), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n982), .A2(new_n868), .A3(new_n984), .ZN(new_n1012));
  NAND2_X1  g826(.A1(G472), .A2(G902), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1013), .B(KEYINPUT63), .Z(new_n1014));
  AOI21_X1  g828(.A(new_n1011), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n325), .A2(new_n306), .A3(new_n307), .ZN(new_n1016));
  AND3_X1   g830(.A1(new_n922), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n324), .A2(new_n266), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n996), .A2(new_n998), .A3(new_n868), .A4(new_n999), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1018), .B1(new_n1019), .B2(new_n1014), .ZN(new_n1020));
  NOR4_X1   g834(.A1(new_n1015), .A2(new_n1017), .A3(new_n1020), .A4(new_n938), .ZN(G57));
endmodule


