

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806;

  BUF_X1 U376 ( .A(n750), .Z(n354) );
  AND2_X1 U377 ( .A1(n456), .A2(n454), .ZN(n453) );
  OR2_X1 U378 ( .A1(n687), .A2(n753), .ZN(n368) );
  AND2_X1 U379 ( .A1(n542), .A2(n541), .ZN(n618) );
  XNOR2_X1 U380 ( .A(n423), .B(n422), .ZN(n404) );
  XNOR2_X1 U381 ( .A(n547), .B(n499), .ZN(n405) );
  BUF_X1 U382 ( .A(G104), .Z(n359) );
  NOR2_X2 U383 ( .A1(G237), .A2(G953), .ZN(n489) );
  NOR2_X2 U384 ( .A1(n640), .A2(n639), .ZN(n715) );
  AND2_X2 U385 ( .A1(n467), .A2(n443), .ZN(n441) );
  XNOR2_X2 U386 ( .A(n577), .B(KEYINPUT111), .ZN(n682) );
  XNOR2_X2 U387 ( .A(G143), .B(G128), .ZN(n547) );
  INV_X4 U388 ( .A(G146), .ZN(n688) );
  XNOR2_X2 U389 ( .A(n473), .B(n472), .ZN(n609) );
  BUF_X1 U390 ( .A(n805), .Z(n355) );
  XOR2_X1 U391 ( .A(KEYINPUT95), .B(KEYINPUT81), .Z(n373) );
  NAND2_X2 U392 ( .A1(n465), .A2(n482), .ZN(n357) );
  AND2_X2 U393 ( .A1(n783), .A2(n664), .ZN(n665) );
  XNOR2_X2 U394 ( .A(G137), .B(G128), .ZN(n463) );
  NOR2_X2 U395 ( .A1(n702), .A2(G902), .ZN(n539) );
  NOR2_X2 U396 ( .A1(n576), .A2(n642), .ZN(n577) );
  XNOR2_X2 U397 ( .A(n636), .B(n635), .ZN(n645) );
  NAND2_X1 U398 ( .A1(n401), .A2(n611), .ZN(n707) );
  XNOR2_X1 U399 ( .A(G902), .B(KEYINPUT15), .ZN(n666) );
  INV_X4 U400 ( .A(G953), .ZN(n797) );
  NOR2_X1 U401 ( .A1(n731), .A2(n730), .ZN(n382) );
  NAND2_X1 U402 ( .A1(n413), .A2(n410), .ZN(n748) );
  XNOR2_X1 U403 ( .A(n496), .B(n495), .ZN(n612) );
  XNOR2_X1 U404 ( .A(n505), .B(n504), .ZN(n611) );
  XNOR2_X1 U405 ( .A(n515), .B(G101), .ZN(n549) );
  XOR2_X1 U406 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n490) );
  INV_X1 U407 ( .A(n660), .ZN(n356) );
  XNOR2_X1 U408 ( .A(n735), .B(n431), .ZN(n658) );
  NOR2_X1 U409 ( .A1(n696), .A2(G902), .ZN(n383) );
  XNOR2_X1 U410 ( .A(n491), .B(n490), .ZN(n358) );
  XNOR2_X1 U411 ( .A(n491), .B(n490), .ZN(n795) );
  XNOR2_X1 U412 ( .A(n551), .B(G140), .ZN(n491) );
  XNOR2_X2 U413 ( .A(n539), .B(n538), .ZN(n637) );
  BUF_X1 U414 ( .A(n672), .Z(n360) );
  XNOR2_X1 U415 ( .A(n451), .B(KEYINPUT45), .ZN(n361) );
  XNOR2_X1 U416 ( .A(n451), .B(KEYINPUT45), .ZN(n783) );
  NOR2_X2 U417 ( .A1(n805), .A2(n715), .ZN(n392) );
  XNOR2_X2 U418 ( .A(n646), .B(KEYINPUT32), .ZN(n805) );
  XNOR2_X1 U419 ( .A(n607), .B(KEYINPUT38), .ZN(n750) );
  INV_X1 U420 ( .A(KEYINPUT68), .ZN(n515) );
  XNOR2_X1 U421 ( .A(n405), .B(n508), .ZN(n564) );
  NAND2_X1 U422 ( .A1(n469), .A2(n374), .ZN(n466) );
  XNOR2_X1 U423 ( .A(n537), .B(n536), .ZN(n538) );
  INV_X1 U424 ( .A(KEYINPUT25), .ZN(n536) );
  XNOR2_X1 U425 ( .A(n487), .B(n398), .ZN(n397) );
  XNOR2_X1 U426 ( .A(G122), .B(KEYINPUT12), .ZN(n487) );
  XNOR2_X1 U427 ( .A(KEYINPUT103), .B(KEYINPUT11), .ZN(n398) );
  XOR2_X1 U428 ( .A(n359), .B(G113), .Z(n488) );
  XNOR2_X1 U429 ( .A(n393), .B(n448), .ZN(n447) );
  XNOR2_X1 U430 ( .A(n572), .B(n548), .ZN(n393) );
  AND2_X1 U431 ( .A1(n367), .A2(n419), .ZN(n418) );
  XNOR2_X1 U432 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U433 ( .A(n523), .B(n522), .ZN(n524) );
  INV_X1 U434 ( .A(KEYINPUT76), .ZN(n522) );
  NAND2_X1 U435 ( .A1(n417), .A2(n749), .ZN(n412) );
  NAND2_X1 U436 ( .A1(n612), .A2(n611), .ZN(n752) );
  OR2_X1 U437 ( .A1(n750), .A2(n417), .ZN(n416) );
  NAND2_X1 U438 ( .A1(n415), .A2(n375), .ZN(n414) );
  OR2_X1 U439 ( .A1(n752), .A2(n400), .ZN(n415) );
  XOR2_X1 U440 ( .A(G119), .B(G113), .Z(n514) );
  XNOR2_X1 U441 ( .A(KEYINPUT5), .B(G116), .ZN(n509) );
  INV_X1 U442 ( .A(G134), .ZN(n499) );
  XNOR2_X1 U443 ( .A(n497), .B(G122), .ZN(n556) );
  XNOR2_X1 U444 ( .A(G116), .B(G107), .ZN(n497) );
  NAND2_X1 U445 ( .A1(n707), .A2(n438), .ZN(n437) );
  NOR2_X1 U446 ( .A1(n707), .A2(n400), .ZN(n542) );
  BUF_X1 U447 ( .A(n735), .Z(n429) );
  INV_X1 U448 ( .A(KEYINPUT1), .ZN(n407) );
  NAND2_X1 U449 ( .A1(n434), .A2(n432), .ZN(n686) );
  NAND2_X1 U450 ( .A1(n433), .A2(n436), .ZN(n432) );
  AND2_X1 U451 ( .A1(n435), .A2(n437), .ZN(n434) );
  NOR2_X1 U452 ( .A1(n707), .A2(n438), .ZN(n436) );
  INV_X1 U453 ( .A(KEYINPUT86), .ZN(n455) );
  NOR2_X1 U454 ( .A1(n686), .A2(n806), .ZN(n615) );
  AND2_X1 U455 ( .A1(n680), .A2(n470), .ZN(n469) );
  NAND2_X1 U456 ( .A1(n723), .A2(KEYINPUT92), .ZN(n470) );
  XOR2_X1 U457 ( .A(KEYINPUT101), .B(KEYINPUT20), .Z(n520) );
  XNOR2_X1 U458 ( .A(n553), .B(KEYINPUT4), .ZN(n450) );
  INV_X1 U459 ( .A(KEYINPUT44), .ZN(n648) );
  INV_X1 U460 ( .A(G237), .ZN(n506) );
  AND2_X1 U461 ( .A1(n669), .A2(n670), .ZN(n477) );
  XNOR2_X1 U462 ( .A(n428), .B(n427), .ZN(n593) );
  INV_X1 U463 ( .A(KEYINPUT72), .ZN(n427) );
  XNOR2_X1 U464 ( .A(n527), .B(KEYINPUT99), .ZN(n624) );
  INV_X1 U465 ( .A(G902), .ZN(n574) );
  INV_X1 U466 ( .A(KEYINPUT6), .ZN(n431) );
  XNOR2_X1 U467 ( .A(n446), .B(n557), .ZN(n786) );
  XNOR2_X1 U468 ( .A(n555), .B(n556), .ZN(n446) );
  INV_X1 U469 ( .A(KEYINPUT77), .ZN(n543) );
  XNOR2_X1 U470 ( .A(n461), .B(G110), .ZN(n460) );
  INV_X1 U471 ( .A(KEYINPUT24), .ZN(n461) );
  XNOR2_X1 U472 ( .A(n488), .B(n369), .ZN(n395) );
  XNOR2_X1 U473 ( .A(n399), .B(n397), .ZN(n396) );
  XNOR2_X1 U474 ( .A(G140), .B(G107), .ZN(n567) );
  XNOR2_X1 U475 ( .A(n425), .B(KEYINPUT80), .ZN(n568) );
  NAND2_X1 U476 ( .A1(n797), .A2(G227), .ZN(n425) );
  NAND2_X1 U477 ( .A1(n362), .A2(n371), .ZN(n729) );
  AND2_X1 U478 ( .A1(n416), .A2(n414), .ZN(n413) );
  NOR2_X1 U479 ( .A1(n752), .A2(n412), .ZN(n411) );
  INV_X1 U480 ( .A(KEYINPUT40), .ZN(n438) );
  INV_X1 U481 ( .A(KEYINPUT79), .ZN(n472) );
  INV_X1 U482 ( .A(KEYINPUT19), .ZN(n422) );
  XNOR2_X1 U483 ( .A(KEYINPUT66), .B(KEYINPUT22), .ZN(n635) );
  XNOR2_X1 U484 ( .A(n517), .B(n516), .ZN(n696) );
  XNOR2_X1 U485 ( .A(n503), .B(n402), .ZN(n775) );
  XNOR2_X1 U486 ( .A(n403), .B(n556), .ZN(n402) );
  XNOR2_X1 U487 ( .A(n498), .B(KEYINPUT105), .ZN(n403) );
  INV_X1 U488 ( .A(n612), .ZN(n401) );
  INV_X1 U489 ( .A(n611), .ZN(n585) );
  NOR2_X1 U490 ( .A1(n429), .A2(n406), .ZN(n652) );
  NOR2_X1 U491 ( .A1(n767), .A2(n376), .ZN(n444) );
  AND2_X1 U492 ( .A1(n361), .A2(KEYINPUT2), .ZN(n362) );
  XOR2_X1 U493 ( .A(n381), .B(KEYINPUT109), .Z(n363) );
  AND2_X1 U494 ( .A1(n729), .A2(n377), .ZN(n364) );
  NOR2_X1 U495 ( .A1(n612), .A2(n611), .ZN(n365) );
  OR2_X1 U496 ( .A1(n765), .A2(n426), .ZN(n366) );
  NOR2_X1 U497 ( .A1(n452), .A2(n657), .ZN(n367) );
  XNOR2_X1 U498 ( .A(G143), .B(G131), .ZN(n369) );
  AND2_X1 U499 ( .A1(n804), .A2(KEYINPUT69), .ZN(n370) );
  INV_X1 U500 ( .A(n749), .ZN(n400) );
  AND2_X1 U501 ( .A1(n380), .A2(n379), .ZN(n371) );
  AND2_X1 U502 ( .A1(n445), .A2(n444), .ZN(n372) );
  NAND2_X1 U503 ( .A1(n621), .A2(n622), .ZN(n374) );
  XOR2_X1 U504 ( .A(KEYINPUT41), .B(KEYINPUT110), .Z(n375) );
  OR2_X1 U505 ( .A1(n426), .A2(n724), .ZN(n376) );
  OR2_X1 U506 ( .A1(n669), .A2(n670), .ZN(n377) );
  XOR2_X1 U507 ( .A(n691), .B(n690), .Z(n378) );
  INV_X1 U508 ( .A(KEYINPUT91), .ZN(n443) );
  AND2_X1 U509 ( .A1(n675), .A2(n426), .ZN(n779) );
  NAND2_X1 U510 ( .A1(n464), .A2(n482), .ZN(n379) );
  NAND2_X1 U511 ( .A1(n464), .A2(n482), .ZN(n467) );
  NAND2_X1 U512 ( .A1(n357), .A2(n466), .ZN(n380) );
  NAND2_X1 U513 ( .A1(n357), .A2(n466), .ZN(n468) );
  BUF_X1 U514 ( .A(n597), .Z(n394) );
  NAND2_X1 U515 ( .A1(n394), .A2(n409), .ZN(n381) );
  NAND2_X1 U516 ( .A1(n394), .A2(n409), .ZN(n408) );
  XNOR2_X1 U517 ( .A(n610), .B(KEYINPUT39), .ZN(n623) );
  AND2_X1 U518 ( .A1(n593), .A2(n658), .ZN(n541) );
  BUF_X1 U519 ( .A(G953), .Z(n426) );
  XNOR2_X1 U520 ( .A(n564), .B(n513), .ZN(n517) );
  XNOR2_X1 U521 ( .A(n596), .B(n595), .ZN(n409) );
  XNOR2_X1 U522 ( .A(n382), .B(KEYINPUT89), .ZN(n445) );
  XNOR2_X2 U523 ( .A(n383), .B(n518), .ZN(n735) );
  NOR2_X1 U524 ( .A1(n459), .A2(n458), .ZN(n384) );
  INV_X1 U525 ( .A(n650), .ZN(n385) );
  NOR2_X2 U526 ( .A1(n459), .A2(n458), .ZN(n774) );
  NOR2_X1 U527 ( .A1(n478), .A2(n670), .ZN(n458) );
  XNOR2_X1 U528 ( .A(n424), .B(KEYINPUT88), .ZN(n478) );
  INV_X1 U529 ( .A(n653), .ZN(n386) );
  XNOR2_X1 U530 ( .A(n565), .B(KEYINPUT100), .ZN(n387) );
  XNOR2_X1 U531 ( .A(n565), .B(KEYINPUT100), .ZN(n794) );
  XNOR2_X1 U532 ( .A(n408), .B(KEYINPUT109), .ZN(n598) );
  XOR2_X1 U533 ( .A(KEYINPUT62), .B(n696), .Z(n697) );
  NOR2_X2 U534 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U535 ( .A1(n447), .A2(n786), .ZN(n390) );
  NAND2_X1 U536 ( .A1(n388), .A2(n389), .ZN(n391) );
  NAND2_X1 U537 ( .A1(n391), .A2(n390), .ZN(n672) );
  INV_X1 U538 ( .A(n447), .ZN(n388) );
  INV_X1 U539 ( .A(n786), .ZN(n389) );
  NAND2_X1 U540 ( .A1(n370), .A2(n392), .ZN(n419) );
  NAND2_X1 U541 ( .A1(n392), .A2(n647), .ZN(n421) );
  NAND2_X1 U542 ( .A1(n453), .A2(n606), .ZN(n485) );
  AND2_X1 U543 ( .A1(n479), .A2(KEYINPUT92), .ZN(n464) );
  NAND2_X1 U544 ( .A1(n480), .A2(n481), .ZN(n479) );
  INV_X1 U545 ( .A(n645), .ZN(n640) );
  XNOR2_X1 U546 ( .A(n546), .B(n547), .ZN(n548) );
  XNOR2_X1 U547 ( .A(n572), .B(n571), .ZN(n573) );
  INV_X1 U548 ( .A(n564), .ZN(n565) );
  XNOR2_X1 U549 ( .A(n396), .B(n395), .ZN(n492) );
  NAND2_X1 U550 ( .A1(n510), .A2(G214), .ZN(n399) );
  XNOR2_X1 U551 ( .A(n489), .B(KEYINPUT78), .ZN(n510) );
  NAND2_X1 U552 ( .A1(n404), .A2(n626), .ZN(n627) );
  NAND2_X1 U553 ( .A1(n598), .A2(n404), .ZN(n600) );
  XNOR2_X1 U554 ( .A(n405), .B(n502), .ZN(n503) );
  INV_X1 U555 ( .A(n394), .ZN(n406) );
  XNOR2_X2 U556 ( .A(n597), .B(n407), .ZN(n738) );
  NAND2_X1 U557 ( .A1(n354), .A2(n749), .ZN(n754) );
  NAND2_X1 U558 ( .A1(n750), .A2(n411), .ZN(n410) );
  INV_X1 U559 ( .A(n375), .ZN(n417) );
  NAND2_X1 U560 ( .A1(n420), .A2(n418), .ZN(n451) );
  XNOR2_X1 U561 ( .A(n421), .B(n648), .ZN(n420) );
  NOR2_X2 U562 ( .A1(n607), .A2(n400), .ZN(n423) );
  XNOR2_X2 U563 ( .A(n562), .B(n561), .ZN(n607) );
  XNOR2_X2 U564 ( .A(n632), .B(KEYINPUT35), .ZN(n804) );
  NAND2_X1 U565 ( .A1(n665), .A2(n725), .ZN(n424) );
  XNOR2_X1 U566 ( .A(n463), .B(n486), .ZN(n462) );
  NOR2_X1 U567 ( .A1(n581), .A2(n739), .ZN(n474) );
  OR2_X2 U568 ( .A1(n687), .A2(n601), .ZN(n603) );
  XNOR2_X1 U569 ( .A(n462), .B(n460), .ZN(n533) );
  NAND2_X1 U570 ( .A1(n540), .A2(n637), .ZN(n428) );
  OR2_X1 U571 ( .A1(n386), .A2(n430), .ZN(n649) );
  INV_X1 U572 ( .A(n429), .ZN(n430) );
  INV_X1 U573 ( .A(n623), .ZN(n433) );
  NAND2_X1 U574 ( .A1(n623), .A2(n438), .ZN(n435) );
  NAND2_X1 U575 ( .A1(n439), .A2(KEYINPUT91), .ZN(n442) );
  NAND2_X1 U576 ( .A1(n468), .A2(n379), .ZN(n439) );
  NAND2_X1 U577 ( .A1(n442), .A2(n440), .ZN(n725) );
  NAND2_X1 U578 ( .A1(n441), .A2(n380), .ZN(n440) );
  XNOR2_X2 U579 ( .A(n688), .B(G125), .ZN(n551) );
  XNOR2_X1 U580 ( .A(n552), .B(n449), .ZN(n448) );
  XNOR2_X1 U581 ( .A(n551), .B(n450), .ZN(n449) );
  XNOR2_X2 U582 ( .A(n788), .B(KEYINPUT73), .ZN(n572) );
  INV_X1 U583 ( .A(n706), .ZN(n452) );
  NAND2_X1 U584 ( .A1(n605), .A2(n455), .ZN(n454) );
  NAND2_X1 U585 ( .A1(n457), .A2(n604), .ZN(n456) );
  AND2_X2 U586 ( .A1(n603), .A2(n605), .ZN(n457) );
  NAND2_X1 U587 ( .A1(n471), .A2(n364), .ZN(n459) );
  AND2_X2 U588 ( .A1(n479), .A2(n469), .ZN(n465) );
  NAND2_X1 U589 ( .A1(n478), .A2(n477), .ZN(n471) );
  NAND2_X1 U590 ( .A1(n475), .A2(n474), .ZN(n473) );
  XNOR2_X1 U591 ( .A(n582), .B(n476), .ZN(n475) );
  INV_X1 U592 ( .A(KEYINPUT30), .ZN(n476) );
  NOR2_X1 U593 ( .A1(n616), .A2(n617), .ZN(n480) );
  INV_X1 U594 ( .A(n485), .ZN(n481) );
  AND2_X2 U595 ( .A1(n484), .A2(n483), .ZN(n482) );
  NAND2_X1 U596 ( .A1(n616), .A2(n617), .ZN(n483) );
  NAND2_X1 U597 ( .A1(n485), .A2(n617), .ZN(n484) );
  NAND2_X1 U598 ( .A1(n693), .A2(n699), .ZN(n695) );
  XNOR2_X1 U599 ( .A(n692), .B(n378), .ZN(n693) );
  XNOR2_X1 U600 ( .A(n554), .B(KEYINPUT75), .ZN(n555) );
  BUF_X1 U601 ( .A(n637), .Z(n733) );
  XNOR2_X2 U602 ( .A(G119), .B(KEYINPUT23), .ZN(n486) );
  INV_X1 U603 ( .A(KEYINPUT18), .ZN(n553) );
  XNOR2_X1 U604 ( .A(n494), .B(n493), .ZN(n495) );
  BUF_X1 U605 ( .A(n725), .Z(n796) );
  XNOR2_X1 U606 ( .A(n492), .B(n358), .ZN(n691) );
  NOR2_X1 U607 ( .A1(G902), .A2(n691), .ZN(n496) );
  XNOR2_X1 U608 ( .A(KEYINPUT104), .B(KEYINPUT13), .ZN(n494) );
  INV_X1 U609 ( .A(G475), .ZN(n493) );
  XOR2_X1 U610 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n498) );
  NAND2_X1 U611 ( .A1(n797), .A2(G234), .ZN(n501) );
  XNOR2_X1 U612 ( .A(KEYINPUT87), .B(KEYINPUT8), .ZN(n500) );
  XNOR2_X1 U613 ( .A(n501), .B(n500), .ZN(n531) );
  NAND2_X1 U614 ( .A1(n531), .A2(G217), .ZN(n502) );
  NAND2_X1 U615 ( .A1(n775), .A2(n574), .ZN(n505) );
  INV_X1 U616 ( .A(G478), .ZN(n504) );
  NAND2_X1 U617 ( .A1(n574), .A2(n506), .ZN(n558) );
  NAND2_X1 U618 ( .A1(n558), .A2(G214), .ZN(n749) );
  XNOR2_X1 U619 ( .A(G137), .B(G131), .ZN(n507) );
  XNOR2_X1 U620 ( .A(n507), .B(KEYINPUT4), .ZN(n508) );
  XNOR2_X1 U621 ( .A(n509), .B(KEYINPUT102), .ZN(n512) );
  NAND2_X1 U622 ( .A1(n510), .A2(G210), .ZN(n511) );
  XNOR2_X1 U623 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U624 ( .A(n514), .B(KEYINPUT3), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n549), .B(n688), .ZN(n566) );
  XNOR2_X1 U626 ( .A(n566), .B(n557), .ZN(n516) );
  INV_X1 U627 ( .A(G472), .ZN(n518) );
  NAND2_X1 U628 ( .A1(G234), .A2(n666), .ZN(n519) );
  XNOR2_X1 U629 ( .A(n520), .B(n519), .ZN(n535) );
  NAND2_X1 U630 ( .A1(n535), .A2(G221), .ZN(n521) );
  XNOR2_X1 U631 ( .A(n521), .B(KEYINPUT21), .ZN(n732) );
  INV_X1 U632 ( .A(n732), .ZN(n530) );
  XOR2_X1 U633 ( .A(KEYINPUT98), .B(KEYINPUT14), .Z(n525) );
  NAND2_X1 U634 ( .A1(G234), .A2(G237), .ZN(n523) );
  NAND2_X1 U635 ( .A1(G952), .A2(n526), .ZN(n765) );
  NAND2_X1 U636 ( .A1(n526), .A2(G902), .ZN(n527) );
  NAND2_X1 U637 ( .A1(n426), .A2(n624), .ZN(n528) );
  OR2_X1 U638 ( .A1(n528), .A2(G900), .ZN(n529) );
  NAND2_X1 U639 ( .A1(n366), .A2(n529), .ZN(n580) );
  AND2_X1 U640 ( .A1(n530), .A2(n580), .ZN(n540) );
  NAND2_X1 U641 ( .A1(G221), .A2(n531), .ZN(n532) );
  XNOR2_X1 U642 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U643 ( .A(n534), .B(n795), .ZN(n702) );
  NAND2_X1 U644 ( .A1(n535), .A2(G217), .ZN(n537) );
  XNOR2_X2 U645 ( .A(G110), .B(G104), .ZN(n544) );
  XNOR2_X2 U646 ( .A(n544), .B(n543), .ZN(n788) );
  NAND2_X1 U647 ( .A1(G224), .A2(n797), .ZN(n545) );
  XNOR2_X1 U648 ( .A(n373), .B(n545), .ZN(n546) );
  XOR2_X1 U649 ( .A(KEYINPUT96), .B(KEYINPUT17), .Z(n550) );
  XNOR2_X1 U650 ( .A(n549), .B(n550), .ZN(n552) );
  XOR2_X1 U651 ( .A(KEYINPUT74), .B(KEYINPUT16), .Z(n554) );
  NAND2_X1 U652 ( .A1(n672), .A2(n666), .ZN(n562) );
  XOR2_X1 U653 ( .A(KEYINPUT84), .B(KEYINPUT97), .Z(n560) );
  NAND2_X1 U654 ( .A1(n558), .A2(G210), .ZN(n559) );
  XNOR2_X1 U655 ( .A(n560), .B(n559), .ZN(n561) );
  INV_X1 U656 ( .A(n607), .ZN(n583) );
  NAND2_X1 U657 ( .A1(n618), .A2(n583), .ZN(n563) );
  XNOR2_X1 U658 ( .A(n563), .B(KEYINPUT36), .ZN(n576) );
  INV_X1 U659 ( .A(n566), .ZN(n570) );
  XNOR2_X1 U660 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U661 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U662 ( .A(n794), .B(n573), .ZN(n770) );
  NAND2_X1 U663 ( .A1(n770), .A2(n574), .ZN(n575) );
  XNOR2_X2 U664 ( .A(n575), .B(G469), .ZN(n597) );
  XNOR2_X1 U665 ( .A(n738), .B(KEYINPUT94), .ZN(n642) );
  XNOR2_X1 U666 ( .A(n682), .B(KEYINPUT93), .ZN(n592) );
  NOR2_X1 U667 ( .A1(n637), .A2(n732), .ZN(n579) );
  INV_X1 U668 ( .A(KEYINPUT70), .ZN(n578) );
  XNOR2_X1 U669 ( .A(n579), .B(n578), .ZN(n739) );
  NAND2_X1 U670 ( .A1(n597), .A2(n580), .ZN(n581) );
  NAND2_X1 U671 ( .A1(n735), .A2(n749), .ZN(n582) );
  NAND2_X1 U672 ( .A1(n583), .A2(n365), .ZN(n584) );
  NOR2_X1 U673 ( .A1(n609), .A2(n584), .ZN(n716) );
  INV_X1 U674 ( .A(n716), .ZN(n590) );
  AND2_X1 U675 ( .A1(n612), .A2(n585), .ZN(n720) );
  INV_X1 U676 ( .A(n720), .ZN(n586) );
  NAND2_X1 U677 ( .A1(n586), .A2(n707), .ZN(n588) );
  INV_X1 U678 ( .A(KEYINPUT106), .ZN(n587) );
  XNOR2_X1 U679 ( .A(n588), .B(n587), .ZN(n753) );
  NAND2_X1 U680 ( .A1(n753), .A2(KEYINPUT47), .ZN(n589) );
  NAND2_X1 U681 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U682 ( .A1(n592), .A2(n591), .ZN(n606) );
  NAND2_X1 U683 ( .A1(n593), .A2(n735), .ZN(n596) );
  INV_X1 U684 ( .A(KEYINPUT108), .ZN(n594) );
  XNOR2_X1 U685 ( .A(n594), .B(KEYINPUT28), .ZN(n595) );
  INV_X1 U686 ( .A(KEYINPUT83), .ZN(n599) );
  XNOR2_X2 U687 ( .A(n600), .B(n599), .ZN(n687) );
  INV_X1 U688 ( .A(KEYINPUT47), .ZN(n601) );
  NAND2_X1 U689 ( .A1(n368), .A2(n601), .ZN(n604) );
  INV_X1 U690 ( .A(n687), .ZN(n683) );
  NOR2_X1 U691 ( .A1(n601), .A2(KEYINPUT86), .ZN(n602) );
  NAND2_X1 U692 ( .A1(n687), .A2(n602), .ZN(n605) );
  INV_X1 U693 ( .A(n750), .ZN(n608) );
  NOR2_X1 U694 ( .A1(n748), .A2(n363), .ZN(n613) );
  XNOR2_X1 U695 ( .A(n613), .B(KEYINPUT42), .ZN(n806) );
  XOR2_X1 U696 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n614) );
  XNOR2_X1 U697 ( .A(n615), .B(n614), .ZN(n616) );
  INV_X1 U698 ( .A(KEYINPUT48), .ZN(n617) );
  NAND2_X1 U699 ( .A1(n618), .A2(n738), .ZN(n619) );
  XNOR2_X1 U700 ( .A(n619), .B(KEYINPUT43), .ZN(n620) );
  AND2_X1 U701 ( .A1(n607), .A2(n620), .ZN(n723) );
  INV_X1 U702 ( .A(n723), .ZN(n621) );
  INV_X1 U703 ( .A(KEYINPUT92), .ZN(n622) );
  NAND2_X1 U704 ( .A1(n433), .A2(n720), .ZN(n680) );
  NOR2_X1 U705 ( .A1(G898), .A2(n797), .ZN(n790) );
  NAND2_X1 U706 ( .A1(n790), .A2(n624), .ZN(n625) );
  NAND2_X1 U707 ( .A1(n625), .A2(n366), .ZN(n626) );
  XNOR2_X2 U708 ( .A(n627), .B(KEYINPUT0), .ZN(n655) );
  INV_X1 U709 ( .A(n739), .ZN(n653) );
  NAND2_X1 U710 ( .A1(n653), .A2(n658), .ZN(n628) );
  NOR2_X1 U711 ( .A1(n628), .A2(n738), .ZN(n629) );
  XNOR2_X1 U712 ( .A(n629), .B(KEYINPUT33), .ZN(n757) );
  NOR2_X1 U713 ( .A1(n655), .A2(n757), .ZN(n630) );
  XNOR2_X1 U714 ( .A(n630), .B(KEYINPUT34), .ZN(n631) );
  NAND2_X1 U715 ( .A1(n631), .A2(n365), .ZN(n632) );
  NOR2_X1 U716 ( .A1(n804), .A2(KEYINPUT69), .ZN(n647) );
  NOR2_X1 U717 ( .A1(n732), .A2(n752), .ZN(n633) );
  XNOR2_X1 U718 ( .A(n633), .B(KEYINPUT107), .ZN(n634) );
  NOR2_X2 U719 ( .A1(n655), .A2(n634), .ZN(n636) );
  INV_X1 U720 ( .A(n733), .ZN(n659) );
  NOR2_X1 U721 ( .A1(n429), .A2(n659), .ZN(n638) );
  NAND2_X1 U722 ( .A1(n738), .A2(n638), .ZN(n639) );
  XNOR2_X1 U723 ( .A(n356), .B(KEYINPUT82), .ZN(n641) );
  OR2_X1 U724 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U725 ( .A1(n643), .A2(n659), .ZN(n644) );
  AND2_X2 U726 ( .A1(n645), .A2(n644), .ZN(n646) );
  INV_X1 U727 ( .A(n655), .ZN(n650) );
  NOR2_X1 U728 ( .A1(n649), .A2(n738), .ZN(n744) );
  NAND2_X1 U729 ( .A1(n650), .A2(n744), .ZN(n651) );
  XNOR2_X1 U730 ( .A(n651), .B(KEYINPUT31), .ZN(n721) );
  NAND2_X1 U731 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U732 ( .A1(n385), .A2(n654), .ZN(n710) );
  NOR2_X1 U733 ( .A1(n721), .A2(n710), .ZN(n656) );
  NOR2_X1 U734 ( .A1(n753), .A2(n656), .ZN(n657) );
  INV_X1 U735 ( .A(n738), .ZN(n662) );
  INV_X1 U736 ( .A(n658), .ZN(n660) );
  NAND2_X1 U737 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U738 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U739 ( .A1(n645), .A2(n663), .ZN(n706) );
  INV_X1 U740 ( .A(n666), .ZN(n664) );
  XOR2_X1 U741 ( .A(KEYINPUT90), .B(n666), .Z(n667) );
  NAND2_X1 U742 ( .A1(n667), .A2(KEYINPUT2), .ZN(n668) );
  XOR2_X1 U743 ( .A(KEYINPUT67), .B(n668), .Z(n669) );
  INV_X1 U744 ( .A(KEYINPUT65), .ZN(n670) );
  NAND2_X1 U745 ( .A1(n774), .A2(G210), .ZN(n674) );
  XOR2_X1 U746 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n671) );
  XNOR2_X1 U747 ( .A(n360), .B(n671), .ZN(n673) );
  XNOR2_X1 U748 ( .A(n674), .B(n673), .ZN(n676) );
  INV_X1 U749 ( .A(G952), .ZN(n675) );
  INV_X1 U750 ( .A(n779), .ZN(n699) );
  NAND2_X1 U751 ( .A1(n676), .A2(n699), .ZN(n678) );
  INV_X1 U752 ( .A(KEYINPUT56), .ZN(n677) );
  XNOR2_X1 U753 ( .A(n678), .B(n677), .ZN(G51) );
  XOR2_X1 U754 ( .A(G134), .B(KEYINPUT115), .Z(n679) );
  XNOR2_X1 U755 ( .A(n680), .B(n679), .ZN(G36) );
  XOR2_X1 U756 ( .A(G125), .B(KEYINPUT37), .Z(n681) );
  XNOR2_X1 U757 ( .A(n682), .B(n681), .ZN(G27) );
  NAND2_X1 U758 ( .A1(n683), .A2(n720), .ZN(n685) );
  XOR2_X1 U759 ( .A(G128), .B(KEYINPUT29), .Z(n684) );
  XNOR2_X1 U760 ( .A(n685), .B(n684), .ZN(G30) );
  XOR2_X1 U761 ( .A(n686), .B(G131), .Z(G33) );
  NOR2_X1 U762 ( .A1(n687), .A2(n707), .ZN(n689) );
  XNOR2_X1 U763 ( .A(n689), .B(n688), .ZN(G48) );
  NAND2_X1 U764 ( .A1(n774), .A2(G475), .ZN(n692) );
  XOR2_X1 U765 ( .A(KEYINPUT122), .B(KEYINPUT59), .Z(n690) );
  XNOR2_X1 U766 ( .A(KEYINPUT123), .B(KEYINPUT60), .ZN(n694) );
  XNOR2_X1 U767 ( .A(n695), .B(n694), .ZN(G60) );
  NAND2_X1 U768 ( .A1(n774), .A2(G472), .ZN(n698) );
  XNOR2_X1 U769 ( .A(n698), .B(n697), .ZN(n700) );
  NAND2_X1 U770 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U771 ( .A(n701), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U772 ( .A1(n384), .A2(G217), .ZN(n704) );
  XOR2_X1 U773 ( .A(n702), .B(KEYINPUT125), .Z(n703) );
  XNOR2_X1 U774 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U775 ( .A1(n705), .A2(n779), .ZN(G66) );
  XNOR2_X1 U776 ( .A(G101), .B(n706), .ZN(G3) );
  INV_X1 U777 ( .A(n707), .ZN(n717) );
  NAND2_X1 U778 ( .A1(n710), .A2(n717), .ZN(n708) );
  XNOR2_X1 U779 ( .A(n708), .B(KEYINPUT112), .ZN(n709) );
  XNOR2_X1 U780 ( .A(n359), .B(n709), .ZN(G6) );
  XOR2_X1 U781 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n712) );
  NAND2_X1 U782 ( .A1(n710), .A2(n720), .ZN(n711) );
  XNOR2_X1 U783 ( .A(n712), .B(n711), .ZN(n714) );
  XOR2_X1 U784 ( .A(G107), .B(KEYINPUT113), .Z(n713) );
  XNOR2_X1 U785 ( .A(n714), .B(n713), .ZN(G9) );
  XOR2_X1 U786 ( .A(n715), .B(G110), .Z(G12) );
  XOR2_X1 U787 ( .A(G143), .B(n716), .Z(G45) );
  NAND2_X1 U788 ( .A1(n721), .A2(n717), .ZN(n718) );
  XNOR2_X1 U789 ( .A(n718), .B(KEYINPUT114), .ZN(n719) );
  XNOR2_X1 U790 ( .A(G113), .B(n719), .ZN(G15) );
  NAND2_X1 U791 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U792 ( .A(n722), .B(G116), .ZN(G18) );
  XOR2_X1 U793 ( .A(G140), .B(n723), .Z(G42) );
  NOR2_X1 U794 ( .A1(n748), .A2(n757), .ZN(n724) );
  NAND2_X1 U795 ( .A1(n796), .A2(n361), .ZN(n727) );
  INV_X1 U796 ( .A(KEYINPUT2), .ZN(n726) );
  NAND2_X1 U797 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U798 ( .A(n728), .B(KEYINPUT85), .ZN(n731) );
  INV_X1 U799 ( .A(n729), .ZN(n730) );
  XOR2_X1 U800 ( .A(KEYINPUT52), .B(KEYINPUT120), .Z(n764) );
  NAND2_X1 U801 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U802 ( .A(KEYINPUT49), .B(n734), .ZN(n736) );
  NOR2_X1 U803 ( .A1(n736), .A2(n429), .ZN(n737) );
  XOR2_X1 U804 ( .A(KEYINPUT116), .B(n737), .Z(n742) );
  NAND2_X1 U805 ( .A1(n386), .A2(n738), .ZN(n740) );
  XOR2_X1 U806 ( .A(KEYINPUT50), .B(n740), .Z(n741) );
  NOR2_X1 U807 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U808 ( .A(KEYINPUT117), .B(n743), .Z(n745) );
  NOR2_X1 U809 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U810 ( .A(KEYINPUT51), .B(n746), .Z(n747) );
  NOR2_X1 U811 ( .A1(n748), .A2(n747), .ZN(n761) );
  NOR2_X1 U812 ( .A1(n354), .A2(n749), .ZN(n751) );
  NOR2_X1 U813 ( .A1(n752), .A2(n751), .ZN(n756) );
  NOR2_X1 U814 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U815 ( .A1(n756), .A2(n755), .ZN(n758) );
  NOR2_X1 U816 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U817 ( .A(n759), .B(KEYINPUT118), .ZN(n760) );
  NOR2_X1 U818 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U819 ( .A(n762), .B(KEYINPUT119), .ZN(n763) );
  XNOR2_X1 U820 ( .A(n764), .B(n763), .ZN(n766) );
  NOR2_X1 U821 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U822 ( .A(KEYINPUT53), .B(n372), .ZN(G75) );
  NAND2_X1 U823 ( .A1(n384), .A2(G469), .ZN(n772) );
  XNOR2_X1 U824 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n768) );
  XOR2_X1 U825 ( .A(n768), .B(KEYINPUT57), .Z(n769) );
  XNOR2_X1 U826 ( .A(n770), .B(n769), .ZN(n771) );
  XNOR2_X1 U827 ( .A(n772), .B(n771), .ZN(n773) );
  NOR2_X1 U828 ( .A1(n779), .A2(n773), .ZN(G54) );
  NAND2_X1 U829 ( .A1(n384), .A2(G478), .ZN(n777) );
  XOR2_X1 U830 ( .A(KEYINPUT124), .B(n775), .Z(n776) );
  XNOR2_X1 U831 ( .A(n777), .B(n776), .ZN(n778) );
  NOR2_X1 U832 ( .A1(n779), .A2(n778), .ZN(G63) );
  NAND2_X1 U833 ( .A1(G224), .A2(n426), .ZN(n780) );
  XNOR2_X1 U834 ( .A(n780), .B(KEYINPUT126), .ZN(n781) );
  XNOR2_X1 U835 ( .A(KEYINPUT61), .B(n781), .ZN(n782) );
  NAND2_X1 U836 ( .A1(G898), .A2(n782), .ZN(n785) );
  NAND2_X1 U837 ( .A1(n361), .A2(n797), .ZN(n784) );
  NAND2_X1 U838 ( .A1(n785), .A2(n784), .ZN(n792) );
  XOR2_X1 U839 ( .A(G101), .B(n786), .Z(n787) );
  XNOR2_X1 U840 ( .A(n788), .B(n787), .ZN(n789) );
  NOR2_X1 U841 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U842 ( .A(n792), .B(n791), .Z(n793) );
  XNOR2_X1 U843 ( .A(KEYINPUT127), .B(n793), .ZN(G69) );
  XOR2_X1 U844 ( .A(n387), .B(n358), .Z(n799) );
  XNOR2_X1 U845 ( .A(n796), .B(n799), .ZN(n798) );
  NAND2_X1 U846 ( .A1(n798), .A2(n797), .ZN(n803) );
  XOR2_X1 U847 ( .A(G227), .B(n799), .Z(n800) );
  NAND2_X1 U848 ( .A1(n800), .A2(G900), .ZN(n801) );
  NAND2_X1 U849 ( .A1(n801), .A2(n426), .ZN(n802) );
  NAND2_X1 U850 ( .A1(n803), .A2(n802), .ZN(G72) );
  XOR2_X1 U851 ( .A(n804), .B(G122), .Z(G24) );
  XOR2_X1 U852 ( .A(n355), .B(G119), .Z(G21) );
  XOR2_X1 U853 ( .A(G137), .B(n806), .Z(G39) );
endmodule

