

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595;

  XNOR2_X2 U324 ( .A(n311), .B(G64GAT), .ZN(n355) );
  XNOR2_X2 U325 ( .A(G176GAT), .B(G92GAT), .ZN(n311) );
  NOR2_X2 U326 ( .A1(n484), .A2(n483), .ZN(n570) );
  OR2_X1 U327 ( .A1(n575), .A2(n481), .ZN(n482) );
  INV_X1 U328 ( .A(KEYINPUT95), .ZN(n376) );
  NAND2_X1 U329 ( .A1(n412), .A2(n411), .ZN(n498) );
  XOR2_X1 U330 ( .A(n369), .B(n368), .Z(n292) );
  NOR2_X1 U331 ( .A1(n593), .A2(n496), .ZN(n463) );
  INV_X1 U332 ( .A(n426), .ZN(n427) );
  XNOR2_X1 U333 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U334 ( .A(n430), .B(n429), .ZN(n432) );
  XNOR2_X1 U335 ( .A(n370), .B(n292), .ZN(n371) );
  XNOR2_X1 U336 ( .A(n372), .B(n371), .ZN(n375) );
  XNOR2_X1 U337 ( .A(n558), .B(n435), .ZN(n593) );
  XNOR2_X1 U338 ( .A(n456), .B(KEYINPUT38), .ZN(n457) );
  XOR2_X1 U339 ( .A(n480), .B(KEYINPUT28), .Z(n537) );
  XNOR2_X1 U340 ( .A(n458), .B(n457), .ZN(n516) );
  XNOR2_X1 U341 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n485) );
  XNOR2_X1 U342 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U343 ( .A(n486), .B(n485), .ZN(G1351GAT) );
  XNOR2_X1 U344 ( .A(n462), .B(n461), .ZN(G1330GAT) );
  XOR2_X1 U345 ( .A(G8GAT), .B(G113GAT), .Z(n294) );
  XNOR2_X1 U346 ( .A(G169GAT), .B(G141GAT), .ZN(n293) );
  XNOR2_X1 U347 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U348 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n296) );
  XNOR2_X1 U349 ( .A(G1GAT), .B(KEYINPUT65), .ZN(n295) );
  XNOR2_X1 U350 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U351 ( .A(n298), .B(n297), .ZN(n310) );
  XNOR2_X1 U352 ( .A(G197GAT), .B(G29GAT), .ZN(n299) );
  XNOR2_X1 U353 ( .A(n299), .B(G50GAT), .ZN(n301) );
  XNOR2_X1 U354 ( .A(G22GAT), .B(G15GAT), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n300), .B(KEYINPUT68), .ZN(n442) );
  XOR2_X1 U356 ( .A(n301), .B(n442), .Z(n308) );
  XOR2_X1 U357 ( .A(G43GAT), .B(KEYINPUT8), .Z(n303) );
  XNOR2_X1 U358 ( .A(KEYINPUT7), .B(KEYINPUT67), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n303), .B(n302), .ZN(n425) );
  XOR2_X1 U360 ( .A(n425), .B(KEYINPUT66), .Z(n305) );
  NAND2_X1 U361 ( .A1(G229GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U362 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U363 ( .A(n306), .B(G36GAT), .ZN(n307) );
  XNOR2_X1 U364 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U365 ( .A(n310), .B(n309), .ZN(n579) );
  XOR2_X1 U366 ( .A(G120GAT), .B(G148GAT), .Z(n363) );
  XOR2_X1 U367 ( .A(n363), .B(n355), .Z(n313) );
  NAND2_X1 U368 ( .A1(G230GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n313), .B(n312), .ZN(n315) );
  INV_X1 U370 ( .A(KEYINPUT33), .ZN(n314) );
  XNOR2_X1 U371 ( .A(n315), .B(n314), .ZN(n318) );
  XNOR2_X1 U372 ( .A(G99GAT), .B(G85GAT), .ZN(n316) );
  XNOR2_X1 U373 ( .A(n316), .B(KEYINPUT72), .ZN(n417) );
  XNOR2_X1 U374 ( .A(n417), .B(KEYINPUT32), .ZN(n317) );
  XNOR2_X1 U375 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U376 ( .A(KEYINPUT70), .B(KEYINPUT69), .Z(n320) );
  XNOR2_X1 U377 ( .A(KEYINPUT31), .B(KEYINPUT73), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U379 ( .A(n322), .B(n321), .ZN(n327) );
  XOR2_X1 U380 ( .A(G78GAT), .B(G204GAT), .Z(n324) );
  XNOR2_X1 U381 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n323) );
  XNOR2_X1 U382 ( .A(n324), .B(n323), .ZN(n332) );
  XNOR2_X1 U383 ( .A(G71GAT), .B(G57GAT), .ZN(n325) );
  XNOR2_X1 U384 ( .A(n325), .B(KEYINPUT13), .ZN(n436) );
  XOR2_X1 U385 ( .A(n332), .B(n436), .Z(n326) );
  XNOR2_X1 U386 ( .A(n327), .B(n326), .ZN(n584) );
  NAND2_X1 U387 ( .A1(n579), .A2(n584), .ZN(n500) );
  XOR2_X1 U388 ( .A(G211GAT), .B(KEYINPUT21), .Z(n329) );
  XNOR2_X1 U389 ( .A(G197GAT), .B(KEYINPUT86), .ZN(n328) );
  XNOR2_X1 U390 ( .A(n329), .B(n328), .ZN(n346) );
  XOR2_X1 U391 ( .A(KEYINPUT24), .B(n346), .Z(n331) );
  XOR2_X1 U392 ( .A(G50GAT), .B(G218GAT), .Z(n424) );
  XNOR2_X1 U393 ( .A(G22GAT), .B(n424), .ZN(n330) );
  XNOR2_X1 U394 ( .A(n331), .B(n330), .ZN(n336) );
  XOR2_X1 U395 ( .A(n332), .B(KEYINPUT23), .Z(n334) );
  NAND2_X1 U396 ( .A1(G228GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U397 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U398 ( .A(n336), .B(n335), .Z(n345) );
  XNOR2_X1 U399 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n337) );
  XNOR2_X1 U400 ( .A(n337), .B(KEYINPUT87), .ZN(n338) );
  XOR2_X1 U401 ( .A(n338), .B(KEYINPUT2), .Z(n340) );
  XNOR2_X1 U402 ( .A(G141GAT), .B(G162GAT), .ZN(n339) );
  XNOR2_X1 U403 ( .A(n340), .B(n339), .ZN(n373) );
  XOR2_X1 U404 ( .A(KEYINPUT22), .B(KEYINPUT85), .Z(n342) );
  XNOR2_X1 U405 ( .A(G148GAT), .B(KEYINPUT84), .ZN(n341) );
  XNOR2_X1 U406 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U407 ( .A(n373), .B(n343), .ZN(n344) );
  XNOR2_X1 U408 ( .A(n345), .B(n344), .ZN(n480) );
  XOR2_X1 U409 ( .A(G36GAT), .B(G190GAT), .Z(n426) );
  XNOR2_X1 U410 ( .A(n346), .B(KEYINPUT92), .ZN(n348) );
  AND2_X1 U411 ( .A1(G226GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U412 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U413 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n350) );
  XNOR2_X1 U414 ( .A(G204GAT), .B(G218GAT), .ZN(n349) );
  XOR2_X1 U415 ( .A(n350), .B(n349), .Z(n351) );
  XNOR2_X1 U416 ( .A(n352), .B(n351), .ZN(n357) );
  XOR2_X1 U417 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n354) );
  XNOR2_X1 U418 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n353) );
  XNOR2_X1 U419 ( .A(n354), .B(n353), .ZN(n392) );
  XNOR2_X1 U420 ( .A(n392), .B(n355), .ZN(n356) );
  XNOR2_X1 U421 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U422 ( .A(n426), .B(n358), .ZN(n359) );
  XOR2_X1 U423 ( .A(G8GAT), .B(G183GAT), .Z(n440) );
  XNOR2_X1 U424 ( .A(n359), .B(n440), .ZN(n533) );
  INV_X1 U425 ( .A(n533), .ZN(n476) );
  XOR2_X1 U426 ( .A(KEYINPUT27), .B(n476), .Z(n402) );
  XNOR2_X1 U427 ( .A(KEYINPUT4), .B(KEYINPUT90), .ZN(n360) );
  XNOR2_X1 U428 ( .A(n360), .B(G57GAT), .ZN(n362) );
  XNOR2_X1 U429 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n361) );
  XNOR2_X1 U430 ( .A(n362), .B(n361), .ZN(n365) );
  XNOR2_X1 U431 ( .A(n363), .B(G85GAT), .ZN(n364) );
  XNOR2_X1 U432 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U433 ( .A(G1GAT), .B(G127GAT), .Z(n441) );
  XOR2_X1 U434 ( .A(n366), .B(n441), .Z(n372) );
  XNOR2_X1 U435 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n367) );
  XNOR2_X1 U436 ( .A(n367), .B(KEYINPUT76), .ZN(n393) );
  XOR2_X1 U437 ( .A(G29GAT), .B(G134GAT), .Z(n422) );
  XNOR2_X1 U438 ( .A(n393), .B(n422), .ZN(n370) );
  XOR2_X1 U439 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n369) );
  NAND2_X1 U440 ( .A1(G225GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U441 ( .A(n373), .B(KEYINPUT5), .ZN(n374) );
  XNOR2_X1 U442 ( .A(n375), .B(n374), .ZN(n409) );
  XNOR2_X1 U443 ( .A(KEYINPUT91), .B(n409), .ZN(n574) );
  NAND2_X1 U444 ( .A1(n402), .A2(n574), .ZN(n377) );
  XNOR2_X1 U445 ( .A(n377), .B(n376), .ZN(n487) );
  NOR2_X1 U446 ( .A1(n537), .A2(n487), .ZN(n400) );
  NAND2_X1 U447 ( .A1(G227GAT), .A2(G233GAT), .ZN(n383) );
  XOR2_X1 U448 ( .A(G176GAT), .B(G183GAT), .Z(n379) );
  XNOR2_X1 U449 ( .A(G43GAT), .B(G190GAT), .ZN(n378) );
  XNOR2_X1 U450 ( .A(n379), .B(n378), .ZN(n381) );
  XOR2_X1 U451 ( .A(G99GAT), .B(G134GAT), .Z(n380) );
  XNOR2_X1 U452 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U453 ( .A(n383), .B(n382), .ZN(n399) );
  XOR2_X1 U454 ( .A(KEYINPUT78), .B(KEYINPUT80), .Z(n385) );
  XNOR2_X1 U455 ( .A(KEYINPUT20), .B(KEYINPUT79), .ZN(n384) );
  XNOR2_X1 U456 ( .A(n385), .B(n384), .ZN(n397) );
  XOR2_X1 U457 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n387) );
  XNOR2_X1 U458 ( .A(KEYINPUT77), .B(G71GAT), .ZN(n386) );
  XNOR2_X1 U459 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U460 ( .A(G120GAT), .B(G127GAT), .Z(n389) );
  XNOR2_X1 U461 ( .A(G15GAT), .B(KEYINPUT83), .ZN(n388) );
  XNOR2_X1 U462 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U463 ( .A(n391), .B(n390), .Z(n395) );
  XNOR2_X1 U464 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U465 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U466 ( .A(n397), .B(n396), .Z(n398) );
  XNOR2_X1 U467 ( .A(n399), .B(n398), .ZN(n484) );
  NAND2_X1 U468 ( .A1(n400), .A2(n484), .ZN(n412) );
  INV_X1 U469 ( .A(n484), .ZN(n535) );
  NOR2_X1 U470 ( .A1(n535), .A2(n480), .ZN(n401) );
  XNOR2_X1 U471 ( .A(n401), .B(KEYINPUT26), .ZN(n576) );
  NAND2_X1 U472 ( .A1(n402), .A2(n576), .ZN(n403) );
  XNOR2_X1 U473 ( .A(KEYINPUT96), .B(n403), .ZN(n408) );
  NOR2_X1 U474 ( .A1(n484), .A2(n476), .ZN(n404) );
  XNOR2_X1 U475 ( .A(KEYINPUT97), .B(n404), .ZN(n405) );
  NAND2_X1 U476 ( .A1(n405), .A2(n480), .ZN(n406) );
  XOR2_X1 U477 ( .A(KEYINPUT25), .B(n406), .Z(n407) );
  NAND2_X1 U478 ( .A1(n408), .A2(n407), .ZN(n410) );
  NAND2_X1 U479 ( .A1(n410), .A2(n409), .ZN(n411) );
  XOR2_X1 U480 ( .A(KEYINPUT64), .B(KEYINPUT10), .Z(n414) );
  XNOR2_X1 U481 ( .A(G162GAT), .B(G106GAT), .ZN(n413) );
  XNOR2_X1 U482 ( .A(n414), .B(n413), .ZN(n434) );
  INV_X1 U483 ( .A(n417), .ZN(n416) );
  INV_X1 U484 ( .A(KEYINPUT9), .ZN(n415) );
  NAND2_X1 U485 ( .A1(n416), .A2(n415), .ZN(n419) );
  NAND2_X1 U486 ( .A1(n417), .A2(KEYINPUT9), .ZN(n418) );
  NAND2_X1 U487 ( .A1(n419), .A2(n418), .ZN(n421) );
  AND2_X1 U488 ( .A1(G232GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U489 ( .A(n421), .B(n420), .ZN(n423) );
  XOR2_X1 U490 ( .A(n423), .B(n422), .Z(n430) );
  XNOR2_X1 U491 ( .A(n425), .B(n424), .ZN(n428) );
  XNOR2_X1 U492 ( .A(G92GAT), .B(KEYINPUT11), .ZN(n431) );
  XNOR2_X1 U493 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U494 ( .A(n434), .B(n433), .ZN(n470) );
  INV_X1 U495 ( .A(n470), .ZN(n558) );
  XNOR2_X1 U496 ( .A(KEYINPUT36), .B(KEYINPUT101), .ZN(n435) );
  XOR2_X1 U497 ( .A(G64GAT), .B(n436), .Z(n438) );
  NAND2_X1 U498 ( .A1(G231GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U499 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U500 ( .A(n440), .B(n439), .Z(n444) );
  XNOR2_X1 U501 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U502 ( .A(n444), .B(n443), .ZN(n452) );
  XOR2_X1 U503 ( .A(KEYINPUT12), .B(G211GAT), .Z(n446) );
  XNOR2_X1 U504 ( .A(G155GAT), .B(G78GAT), .ZN(n445) );
  XNOR2_X1 U505 ( .A(n446), .B(n445), .ZN(n450) );
  XOR2_X1 U506 ( .A(KEYINPUT75), .B(KEYINPUT15), .Z(n448) );
  XNOR2_X1 U507 ( .A(KEYINPUT74), .B(KEYINPUT14), .ZN(n447) );
  XNOR2_X1 U508 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U509 ( .A(n450), .B(n449), .Z(n451) );
  XNOR2_X1 U510 ( .A(n452), .B(n451), .ZN(n496) );
  INV_X1 U511 ( .A(n496), .ZN(n589) );
  NOR2_X1 U512 ( .A1(n593), .A2(n589), .ZN(n453) );
  NAND2_X1 U513 ( .A1(n498), .A2(n453), .ZN(n454) );
  XNOR2_X1 U514 ( .A(KEYINPUT37), .B(n454), .ZN(n455) );
  XOR2_X1 U515 ( .A(KEYINPUT102), .B(n455), .Z(n530) );
  NOR2_X1 U516 ( .A1(n500), .A2(n530), .ZN(n458) );
  INV_X1 U517 ( .A(KEYINPUT103), .ZN(n456) );
  NAND2_X1 U518 ( .A1(n516), .A2(n535), .ZN(n462) );
  XOR2_X1 U519 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n460) );
  INV_X1 U520 ( .A(G43GAT), .ZN(n459) );
  INV_X1 U521 ( .A(KEYINPUT54), .ZN(n478) );
  XNOR2_X1 U522 ( .A(n463), .B(KEYINPUT45), .ZN(n464) );
  NAND2_X1 U523 ( .A1(n464), .A2(n584), .ZN(n465) );
  XNOR2_X1 U524 ( .A(KEYINPUT114), .B(n465), .ZN(n466) );
  NOR2_X1 U525 ( .A1(n466), .A2(n579), .ZN(n474) );
  XNOR2_X1 U526 ( .A(n584), .B(KEYINPUT41), .ZN(n553) );
  NAND2_X1 U527 ( .A1(n579), .A2(n553), .ZN(n467) );
  XNOR2_X1 U528 ( .A(KEYINPUT46), .B(n467), .ZN(n468) );
  XNOR2_X1 U529 ( .A(KEYINPUT112), .B(n496), .ZN(n572) );
  NAND2_X1 U530 ( .A1(n468), .A2(n572), .ZN(n469) );
  XNOR2_X1 U531 ( .A(n469), .B(KEYINPUT113), .ZN(n471) );
  NAND2_X1 U532 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U533 ( .A(n472), .B(KEYINPUT47), .ZN(n473) );
  NOR2_X1 U534 ( .A1(n474), .A2(n473), .ZN(n475) );
  XNOR2_X1 U535 ( .A(n475), .B(KEYINPUT48), .ZN(n488) );
  NOR2_X1 U536 ( .A1(n476), .A2(n488), .ZN(n477) );
  XNOR2_X1 U537 ( .A(n478), .B(n477), .ZN(n575) );
  INV_X1 U538 ( .A(n574), .ZN(n479) );
  NAND2_X1 U539 ( .A1(n480), .A2(n479), .ZN(n481) );
  XOR2_X1 U540 ( .A(KEYINPUT55), .B(n482), .Z(n483) );
  NAND2_X1 U541 ( .A1(n570), .A2(n558), .ZN(n486) );
  NOR2_X1 U542 ( .A1(n488), .A2(n487), .ZN(n551) );
  NAND2_X1 U543 ( .A1(n551), .A2(n535), .ZN(n490) );
  INV_X1 U544 ( .A(KEYINPUT115), .ZN(n489) );
  XNOR2_X1 U545 ( .A(n490), .B(n489), .ZN(n491) );
  NOR2_X1 U546 ( .A1(n491), .A2(n537), .ZN(n492) );
  XNOR2_X1 U547 ( .A(KEYINPUT116), .B(n492), .ZN(n547) );
  INV_X1 U548 ( .A(n547), .ZN(n493) );
  NOR2_X1 U549 ( .A1(n493), .A2(n572), .ZN(n494) );
  XNOR2_X1 U550 ( .A(KEYINPUT50), .B(n494), .ZN(n495) );
  XOR2_X1 U551 ( .A(G127GAT), .B(n495), .Z(G1342GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT34), .B(KEYINPUT98), .Z(n502) );
  NOR2_X1 U553 ( .A1(n558), .A2(n496), .ZN(n497) );
  XNOR2_X1 U554 ( .A(n497), .B(KEYINPUT16), .ZN(n499) );
  NAND2_X1 U555 ( .A1(n499), .A2(n498), .ZN(n520) );
  NOR2_X1 U556 ( .A1(n500), .A2(n520), .ZN(n508) );
  NAND2_X1 U557 ( .A1(n508), .A2(n574), .ZN(n501) );
  XNOR2_X1 U558 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U559 ( .A(G1GAT), .B(n503), .Z(G1324GAT) );
  NAND2_X1 U560 ( .A1(n508), .A2(n533), .ZN(n504) );
  XNOR2_X1 U561 ( .A(n504), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT99), .B(KEYINPUT35), .Z(n506) );
  NAND2_X1 U563 ( .A1(n508), .A2(n535), .ZN(n505) );
  XNOR2_X1 U564 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U565 ( .A(G15GAT), .B(n507), .Z(G1326GAT) );
  NAND2_X1 U566 ( .A1(n508), .A2(n537), .ZN(n509) );
  XNOR2_X1 U567 ( .A(n509), .B(KEYINPUT100), .ZN(n510) );
  XNOR2_X1 U568 ( .A(G22GAT), .B(n510), .ZN(G1327GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT39), .B(KEYINPUT104), .Z(n512) );
  NAND2_X1 U570 ( .A1(n516), .A2(n574), .ZN(n511) );
  XNOR2_X1 U571 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U572 ( .A(G29GAT), .B(n513), .ZN(G1328GAT) );
  XOR2_X1 U573 ( .A(G36GAT), .B(KEYINPUT105), .Z(n515) );
  NAND2_X1 U574 ( .A1(n533), .A2(n516), .ZN(n514) );
  XNOR2_X1 U575 ( .A(n515), .B(n514), .ZN(G1329GAT) );
  NAND2_X1 U576 ( .A1(n516), .A2(n537), .ZN(n517) );
  XNOR2_X1 U577 ( .A(n517), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U578 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n522) );
  XOR2_X1 U579 ( .A(KEYINPUT107), .B(n553), .Z(n567) );
  INV_X1 U580 ( .A(n579), .ZN(n518) );
  NAND2_X1 U581 ( .A1(n567), .A2(n518), .ZN(n519) );
  XNOR2_X1 U582 ( .A(n519), .B(KEYINPUT108), .ZN(n529) );
  NOR2_X1 U583 ( .A1(n529), .A2(n520), .ZN(n526) );
  NAND2_X1 U584 ( .A1(n526), .A2(n574), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n522), .B(n521), .ZN(G1332GAT) );
  NAND2_X1 U586 ( .A1(n526), .A2(n533), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U588 ( .A(G71GAT), .B(KEYINPUT109), .Z(n525) );
  NAND2_X1 U589 ( .A1(n526), .A2(n535), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(G1334GAT) );
  XOR2_X1 U591 ( .A(G78GAT), .B(KEYINPUT43), .Z(n528) );
  NAND2_X1 U592 ( .A1(n526), .A2(n537), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(G1335GAT) );
  NOR2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n538) );
  NAND2_X1 U595 ( .A1(n574), .A2(n538), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n531), .B(KEYINPUT110), .ZN(n532) );
  XNOR2_X1 U597 ( .A(G85GAT), .B(n532), .ZN(G1336GAT) );
  NAND2_X1 U598 ( .A1(n538), .A2(n533), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n534), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U600 ( .A1(n535), .A2(n538), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n536), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n540) );
  NAND2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U605 ( .A(G106GAT), .B(n541), .ZN(G1339GAT) );
  XOR2_X1 U606 ( .A(G113GAT), .B(KEYINPUT117), .Z(n543) );
  NAND2_X1 U607 ( .A1(n579), .A2(n547), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(G1340GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n545) );
  NAND2_X1 U610 ( .A1(n547), .A2(n567), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(G120GAT), .B(n546), .ZN(G1341GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n549) );
  NAND2_X1 U614 ( .A1(n558), .A2(n547), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U616 ( .A(G134GAT), .B(n550), .Z(G1343GAT) );
  AND2_X1 U617 ( .A1(n551), .A2(n576), .ZN(n559) );
  NAND2_X1 U618 ( .A1(n579), .A2(n559), .ZN(n552) );
  XNOR2_X1 U619 ( .A(G141GAT), .B(n552), .ZN(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n555) );
  NAND2_X1 U621 ( .A1(n559), .A2(n553), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(n556), .ZN(G1345GAT) );
  NAND2_X1 U624 ( .A1(n559), .A2(n589), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n557), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(KEYINPUT120), .ZN(n561) );
  XNOR2_X1 U628 ( .A(G162GAT), .B(n561), .ZN(G1347GAT) );
  XOR2_X1 U629 ( .A(G169GAT), .B(KEYINPUT121), .Z(n563) );
  NAND2_X1 U630 ( .A1(n570), .A2(n579), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n563), .B(n562), .ZN(G1348GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n565) );
  XNOR2_X1 U633 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n564) );
  XNOR2_X1 U634 ( .A(n565), .B(n564), .ZN(n566) );
  XOR2_X1 U635 ( .A(KEYINPUT56), .B(n566), .Z(n569) );
  NAND2_X1 U636 ( .A1(n570), .A2(n567), .ZN(n568) );
  XNOR2_X1 U637 ( .A(n569), .B(n568), .ZN(G1349GAT) );
  INV_X1 U638 ( .A(n570), .ZN(n571) );
  NOR2_X1 U639 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U640 ( .A(G183GAT), .B(n573), .Z(G1350GAT) );
  XOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT60), .Z(n581) );
  NOR2_X1 U642 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(KEYINPUT124), .B(n578), .ZN(n592) );
  INV_X1 U645 ( .A(n592), .ZN(n588) );
  NAND2_X1 U646 ( .A1(n579), .A2(n588), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n583) );
  XOR2_X1 U648 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(G1352GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n586) );
  OR2_X1 U651 ( .A1(n592), .A2(n584), .ZN(n585) );
  XNOR2_X1 U652 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U653 ( .A(G204GAT), .B(n587), .ZN(G1353GAT) );
  XOR2_X1 U654 ( .A(G211GAT), .B(KEYINPUT127), .Z(n591) );
  NAND2_X1 U655 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U656 ( .A(n591), .B(n590), .ZN(G1354GAT) );
  NOR2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U658 ( .A(KEYINPUT62), .B(n594), .Z(n595) );
  XNOR2_X1 U659 ( .A(G218GAT), .B(n595), .ZN(G1355GAT) );
endmodule

