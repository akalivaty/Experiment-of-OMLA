//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 0 1 1 0 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 0 1 0 0 0 1 1 0 1 0 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  OR3_X1    g0006(.A1(new_n206), .A2(KEYINPUT64), .A3(G13), .ZN(new_n207));
  OAI21_X1  g0007(.A(KEYINPUT64), .B1(new_n206), .B2(G13), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  AND2_X1   g0011(.A1(new_n211), .A2(KEYINPUT0), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(KEYINPUT0), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G116), .ZN(new_n216));
  INV_X1    g0016(.A(G270), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n214), .B1(new_n202), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n206), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  AND2_X1   g0022(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  INV_X1    g0023(.A(new_n201), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G50), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n226), .A2(G20), .A3(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n229), .B1(new_n222), .B2(KEYINPUT1), .ZN(new_n230));
  NOR4_X1   g0030(.A1(new_n212), .A2(new_n213), .A3(new_n223), .A4(new_n230), .ZN(G361));
  XOR2_X1   g0031(.A(G250), .B(G257), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT66), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n235), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n202), .A2(G68), .ZN(new_n245));
  INV_X1    g0045(.A(G68), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n244), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G41), .ZN(new_n253));
  OAI211_X1 g0053(.A(G1), .B(G13), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n255), .B1(G41), .B2(G45), .ZN(new_n256));
  AND2_X1   g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G226), .ZN(new_n258));
  INV_X1    g0058(.A(G274), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n258), .B1(new_n259), .B2(new_n256), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT3), .B(G33), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(G222), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G77), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(G1698), .ZN(new_n265));
  INV_X1    g0065(.A(G223), .ZN(new_n266));
  OAI221_X1 g0066(.A(new_n263), .B1(new_n264), .B2(new_n261), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT65), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n227), .B(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n252), .A2(new_n253), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n260), .B1(new_n267), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G179), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n274), .B1(G169), .B2(new_n272), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT67), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g0078(.A1(KEYINPUT67), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AND3_X1   g0080(.A1(new_n269), .A2(KEYINPUT68), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(KEYINPUT68), .B1(new_n269), .B2(new_n280), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G20), .A2(G33), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT69), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT69), .ZN(new_n288));
  INV_X1    g0088(.A(G58), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT8), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n252), .A2(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n285), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n255), .A2(G13), .A3(G20), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n283), .A2(new_n294), .B1(new_n202), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT68), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n278), .A2(new_n279), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n298), .B1(new_n299), .B2(new_n228), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n269), .A2(KEYINPUT68), .A3(new_n280), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n255), .A2(G20), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n302), .A2(G50), .A3(new_n295), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n297), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n275), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n272), .A2(G190), .ZN(new_n308));
  INV_X1    g0108(.A(G200), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n308), .B1(new_n309), .B2(new_n272), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n305), .A2(KEYINPUT9), .ZN(new_n311));
  OR2_X1    g0111(.A1(new_n305), .A2(KEYINPUT9), .ZN(new_n312));
  AOI211_X1 g0112(.A(KEYINPUT10), .B(new_n310), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT10), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n311), .ZN(new_n315));
  INV_X1    g0115(.A(new_n310), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n307), .B1(new_n313), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n295), .B(KEYINPUT70), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n302), .A2(new_n320), .A3(new_n303), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n321), .A2(new_n264), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT71), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n322), .B(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G20), .A2(G77), .ZN(new_n325));
  INV_X1    g0125(.A(new_n284), .ZN(new_n326));
  XOR2_X1   g0126(.A(KEYINPUT15), .B(G87), .Z(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  OAI221_X1 g0128(.A(new_n325), .B1(new_n326), .B2(new_n286), .C1(new_n328), .C2(new_n293), .ZN(new_n329));
  INV_X1    g0129(.A(new_n320), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n283), .A2(new_n329), .B1(new_n264), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G238), .ZN(new_n332));
  INV_X1    g0132(.A(G107), .ZN(new_n333));
  OAI22_X1  g0133(.A1(new_n265), .A2(new_n332), .B1(new_n333), .B2(new_n261), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT3), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G33), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NOR3_X1   g0138(.A1(new_n338), .A2(new_n237), .A3(G1698), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n271), .B1(new_n334), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n256), .A2(new_n259), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n341), .B1(new_n257), .B2(G244), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G190), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(G200), .B2(new_n343), .ZN(new_n346));
  AND3_X1   g0146(.A1(new_n324), .A2(new_n331), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G169), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(G179), .B2(new_n343), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n350), .B1(new_n324), .B2(new_n331), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n291), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n302), .A2(new_n295), .A3(new_n303), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n291), .A2(new_n296), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n289), .A2(new_n246), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n358), .A2(new_n201), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G20), .ZN(new_n360));
  INV_X1    g0160(.A(G159), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n360), .B1(new_n361), .B2(new_n326), .ZN(new_n362));
  INV_X1    g0162(.A(G20), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT7), .B1(new_n338), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(KEYINPUT7), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n261), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(G68), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT78), .ZN(new_n368));
  AOI21_X1  g0168(.A(G20), .B1(new_n336), .B2(new_n337), .ZN(new_n369));
  OAI22_X1  g0169(.A1(new_n369), .A2(KEYINPUT7), .B1(new_n261), .B2(new_n365), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT78), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n371), .A3(G68), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n362), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n302), .B1(new_n373), .B2(KEYINPUT16), .ZN(new_n374));
  AND3_X1   g0174(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT79), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT7), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n376), .A2(G20), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n337), .B2(KEYINPUT79), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT80), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n335), .A2(G33), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT79), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n365), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT80), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT79), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n376), .B1(new_n261), .B2(G20), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n379), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n362), .B1(new_n387), .B2(G68), .ZN(new_n388));
  OR2_X1    g0188(.A1(new_n388), .A2(KEYINPUT16), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n357), .B1(new_n374), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n215), .A2(G1698), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(G223), .B2(G1698), .ZN(new_n392));
  INV_X1    g0192(.A(G87), .ZN(new_n393));
  OAI22_X1  g0193(.A1(new_n392), .A2(new_n338), .B1(new_n252), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n271), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n341), .B1(new_n257), .B2(G232), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(G179), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(new_n348), .B2(new_n397), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT18), .B1(new_n390), .B2(new_n400), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n355), .A2(new_n356), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n359), .A2(G20), .B1(G159), .B2(new_n284), .ZN(new_n403));
  AND3_X1   g0203(.A1(new_n370), .A2(new_n371), .A3(G68), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n371), .B1(new_n370), .B2(G68), .ZN(new_n405));
  OAI211_X1 g0205(.A(KEYINPUT16), .B(new_n403), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n283), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n388), .A2(KEYINPUT16), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n402), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT18), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(new_n410), .A3(new_n399), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n309), .B1(new_n395), .B2(new_n396), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(G190), .B2(new_n397), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n413), .B(new_n402), .C1(new_n407), .C2(new_n408), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT17), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n374), .A2(new_n389), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n417), .A2(KEYINPUT17), .A3(new_n402), .A4(new_n413), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n401), .A2(new_n411), .A3(new_n416), .A4(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n246), .B1(new_n321), .B2(KEYINPUT12), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n330), .A2(KEYINPUT12), .A3(new_n246), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(KEYINPUT12), .B2(new_n296), .ZN(new_n423));
  OR3_X1    g0223(.A1(new_n421), .A2(KEYINPUT75), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT75), .B1(new_n421), .B2(new_n423), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n292), .A2(G77), .B1(G20), .B2(new_n246), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n202), .B2(new_n326), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n283), .A2(new_n427), .ZN(new_n428));
  XOR2_X1   g0228(.A(KEYINPUT74), .B(KEYINPUT11), .Z(new_n429));
  XNOR2_X1  g0229(.A(new_n428), .B(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n424), .A2(new_n425), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n341), .B1(new_n257), .B2(G238), .ZN(new_n433));
  NAND2_X1  g0233(.A1(G33), .A2(G97), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT72), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT72), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n436), .A2(G33), .A3(G97), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n336), .A2(new_n337), .A3(G226), .A4(new_n262), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n336), .A2(new_n337), .A3(G232), .A4(G1698), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n441), .A2(KEYINPUT73), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT73), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n438), .A2(new_n439), .A3(new_n440), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n271), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n433), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT13), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n441), .A2(KEYINPUT73), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n448), .A2(new_n271), .A3(new_n444), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT13), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n449), .A2(new_n450), .A3(new_n433), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G200), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n432), .B(new_n453), .C1(new_n344), .C2(new_n452), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n319), .A2(new_n353), .A3(new_n420), .A4(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT77), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n447), .A2(G179), .A3(new_n451), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT76), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT76), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n447), .A2(new_n459), .A3(G179), .A4(new_n451), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n449), .A2(new_n450), .A3(new_n433), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n450), .B1(new_n449), .B2(new_n433), .ZN(new_n463));
  OAI21_X1  g0263(.A(G169), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT14), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT14), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n452), .A2(new_n466), .A3(G169), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n456), .B1(new_n461), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n466), .B1(new_n452), .B2(G169), .ZN(new_n470));
  AOI211_X1 g0270(.A(KEYINPUT14), .B(new_n348), .C1(new_n447), .C2(new_n451), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n458), .A2(new_n460), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(KEYINPUT77), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n432), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n455), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n296), .A2(new_n333), .ZN(new_n477));
  XNOR2_X1  g0277(.A(new_n477), .B(KEYINPUT25), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n255), .A2(G33), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT81), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(KEYINPUT81), .B1(new_n255), .B2(G33), .ZN(new_n483));
  OR2_X1    g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n302), .A2(new_n484), .A3(new_n295), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n479), .B1(new_n485), .B2(new_n333), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n336), .A2(new_n337), .A3(new_n363), .A4(G87), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT22), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT22), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n261), .A2(new_n489), .A3(new_n363), .A4(G87), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT86), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G33), .A2(G116), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n493), .A2(G20), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT23), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(new_n363), .B2(G107), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n333), .A2(KEYINPUT23), .A3(G20), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n494), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n491), .A2(new_n492), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n492), .B1(new_n491), .B2(new_n498), .ZN(new_n500));
  OAI21_X1  g0300(.A(KEYINPUT24), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n491), .A2(new_n498), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT86), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT24), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n491), .A2(new_n492), .A3(new_n498), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n486), .B1(new_n507), .B2(new_n283), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n261), .A2(G250), .A3(new_n262), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n336), .A2(new_n337), .A3(G257), .A4(G1698), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G294), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n255), .B(G45), .C1(new_n253), .C2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT5), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(G41), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n254), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n512), .A2(new_n271), .B1(new_n517), .B2(G264), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT87), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT82), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n514), .B2(G41), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n253), .A2(KEYINPUT82), .A3(KEYINPUT5), .ZN(new_n522));
  INV_X1    g0322(.A(G45), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n523), .A2(G1), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n514), .A2(G41), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n521), .A2(new_n522), .A3(new_n524), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n254), .A2(G274), .ZN(new_n527));
  OR2_X1    g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n518), .A2(new_n519), .A3(G179), .A4(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n512), .A2(new_n271), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n517), .A2(G264), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n531), .A2(new_n532), .A3(new_n528), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G169), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n519), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n518), .A2(G179), .A3(new_n528), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n530), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n508), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n302), .B1(new_n501), .B2(new_n506), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n533), .A2(G190), .ZN(new_n540));
  AOI21_X1  g0340(.A(G200), .B1(new_n518), .B2(new_n528), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR3_X1   g0342(.A1(new_n539), .A2(new_n542), .A3(new_n486), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n302), .A2(G97), .A3(new_n484), .A4(new_n295), .ZN(new_n545));
  INV_X1    g0345(.A(G97), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n296), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT6), .ZN(new_n548));
  NOR3_X1   g0348(.A1(new_n548), .A2(new_n546), .A3(G107), .ZN(new_n549));
  XNOR2_X1  g0349(.A(G97), .B(G107), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n549), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  OAI22_X1  g0351(.A1(new_n551), .A2(new_n363), .B1(new_n264), .B2(new_n326), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n552), .B1(new_n387), .B2(G107), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n545), .B(new_n547), .C1(new_n553), .C2(new_n302), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n336), .A2(new_n337), .A3(G244), .A4(new_n262), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT4), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n261), .A2(KEYINPUT4), .A3(G244), .A4(new_n262), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n261), .A2(G250), .A3(G1698), .ZN(new_n559));
  NAND2_X1  g0359(.A1(G33), .A2(G283), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n557), .A2(new_n558), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n271), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n254), .B(G257), .C1(new_n513), .C2(new_n515), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n527), .B2(new_n526), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT83), .B1(new_n566), .B2(G179), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n564), .B1(new_n561), .B2(new_n271), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT83), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n568), .A2(new_n569), .A3(new_n273), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n566), .A2(new_n348), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n554), .A2(new_n567), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n562), .A2(G190), .A3(new_n565), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n309), .B2(new_n568), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n572), .B1(new_n554), .B2(new_n574), .ZN(new_n575));
  OAI22_X1  g0375(.A1(new_n516), .A2(new_n217), .B1(new_n526), .B2(new_n527), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n336), .A2(new_n337), .A3(G264), .A4(G1698), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n336), .A2(new_n337), .A3(G257), .A4(new_n262), .ZN(new_n579));
  INV_X1    g0379(.A(G303), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n578), .B(new_n579), .C1(new_n580), .C2(new_n261), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n271), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n348), .B1(new_n577), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(G116), .B1(new_n482), .B2(new_n483), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n283), .A2(new_n330), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n330), .A2(new_n216), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n269), .A2(new_n280), .ZN(new_n587));
  AOI21_X1  g0387(.A(G20), .B1(G33), .B2(G283), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n252), .A2(G97), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n588), .A2(new_n589), .B1(G20), .B2(new_n216), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n587), .A2(KEYINPUT20), .A3(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(KEYINPUT20), .B1(new_n587), .B2(new_n590), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n586), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n583), .B1(new_n585), .B2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT85), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n596), .A2(KEYINPUT21), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n597), .ZN(new_n599));
  INV_X1    g0399(.A(new_n582), .ZN(new_n600));
  OAI211_X1 g0400(.A(G169), .B(new_n599), .C1(new_n600), .C2(new_n576), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n577), .A2(G179), .A3(new_n582), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n302), .A2(G116), .A3(new_n484), .A4(new_n320), .ZN(new_n604));
  INV_X1    g0404(.A(new_n593), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n591), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n604), .A2(new_n606), .A3(new_n586), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n577), .A2(new_n582), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(G200), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n605), .A2(new_n591), .B1(new_n216), .B2(new_n330), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n577), .A2(G190), .A3(new_n582), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n604), .A4(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n598), .A2(new_n608), .A3(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n320), .A2(new_n327), .ZN(new_n615));
  NOR2_X1   g0415(.A1(G97), .A2(G107), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n393), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT19), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n618), .B1(new_n435), .B2(new_n437), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n617), .B1(new_n619), .B2(G20), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n261), .A2(new_n363), .A3(G68), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n363), .A2(G33), .A3(G97), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n618), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(KEYINPUT84), .ZN(new_n624));
  OR2_X1    g0424(.A1(new_n623), .A2(KEYINPUT84), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n620), .A2(new_n621), .A3(new_n624), .A4(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n615), .B1(new_n283), .B2(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n302), .A2(new_n484), .A3(new_n295), .A4(new_n327), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n336), .A2(new_n337), .A3(G238), .A4(new_n262), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n336), .A2(new_n337), .A3(G244), .A4(G1698), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(new_n631), .A3(new_n493), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n271), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n255), .A2(G45), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(G250), .ZN(new_n636));
  OAI22_X1  g0436(.A1(new_n634), .A2(new_n636), .B1(new_n259), .B2(new_n635), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n348), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n637), .B1(new_n271), .B2(new_n632), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n273), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n629), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n639), .A2(new_n344), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n302), .A2(G87), .A3(new_n484), .A4(new_n295), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n639), .A2(G200), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n627), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n643), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n575), .A2(new_n614), .A3(new_n648), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n476), .A2(new_n544), .A3(new_n649), .ZN(G372));
  INV_X1    g0450(.A(new_n307), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n418), .A2(new_n416), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n454), .A2(new_n351), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n652), .B1(new_n653), .B2(new_n475), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n409), .A2(new_n410), .A3(new_n399), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n410), .B1(new_n409), .B2(new_n399), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n313), .A2(new_n317), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n651), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n476), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n640), .A2(new_n642), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n662), .B1(new_n627), .B2(new_n628), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT88), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n644), .B1(new_n647), .B2(new_n664), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n627), .A2(new_n645), .A3(new_n646), .A4(KEYINPUT88), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT26), .ZN(new_n668));
  INV_X1    g0468(.A(new_n572), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(KEYINPUT26), .B1(new_n648), .B2(new_n572), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(new_n643), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT87), .B1(new_n533), .B2(G169), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n533), .A2(new_n273), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n529), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n539), .B2(new_n486), .ZN(new_n676));
  AOI22_X1  g0476(.A1(new_n595), .A2(new_n597), .B1(new_n603), .B2(new_n607), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n554), .A2(new_n574), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n568), .A2(new_n569), .A3(new_n273), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n569), .B1(new_n568), .B2(new_n273), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n568), .A2(G169), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n679), .B1(new_n554), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n508), .B1(new_n540), .B2(new_n541), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n678), .A2(new_n684), .A3(new_n685), .A4(new_n667), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT89), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n575), .A2(new_n543), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n689), .A2(KEYINPUT89), .A3(new_n667), .A4(new_n678), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n672), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n660), .B1(new_n661), .B2(new_n691), .ZN(G369));
  NAND3_X1  g0492(.A1(new_n255), .A2(new_n363), .A3(G13), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G213), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(G343), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n607), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n677), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT90), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n677), .A2(new_n613), .A3(new_n699), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n700), .A2(new_n701), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT91), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n706), .B(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n698), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n544), .B1(new_n508), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n538), .A2(new_n698), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n708), .A2(G330), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n538), .A2(new_n709), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n677), .A2(new_n698), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n544), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n713), .A2(new_n714), .A3(new_n716), .ZN(G399));
  INV_X1    g0517(.A(new_n209), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G41), .ZN(new_n719));
  NOR4_X1   g0519(.A1(new_n719), .A2(new_n255), .A3(G116), .A4(new_n617), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n720), .B1(new_n226), .B2(new_n719), .ZN(new_n721));
  XOR2_X1   g0521(.A(new_n721), .B(KEYINPUT28), .Z(new_n722));
  INV_X1    g0522(.A(KEYINPUT29), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(new_n691), .B2(new_n698), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT96), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT96), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n726), .B(new_n723), .C1(new_n691), .C2(new_n698), .ZN(new_n727));
  INV_X1    g0527(.A(new_n667), .ZN(new_n728));
  OAI21_X1  g0528(.A(KEYINPUT26), .B1(new_n728), .B2(new_n572), .ZN(new_n729));
  OR3_X1    g0529(.A1(new_n648), .A2(new_n572), .A3(KEYINPUT26), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n663), .B(KEYINPUT97), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n729), .A2(new_n686), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(KEYINPUT29), .A3(new_n709), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n725), .A2(new_n727), .A3(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT31), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n566), .A2(new_n533), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n609), .A2(new_n273), .A3(new_n639), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n566), .A2(new_n602), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n518), .A2(new_n641), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT92), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n518), .A2(KEYINPUT92), .A3(new_n641), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n739), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n738), .B1(new_n745), .B2(KEYINPUT30), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT30), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  AOI211_X1 g0548(.A(new_n735), .B(new_n709), .C1(new_n746), .C2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n614), .A2(new_n648), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n544), .A2(new_n684), .A3(new_n750), .A4(new_n709), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(KEYINPUT95), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT95), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n649), .A2(new_n753), .A3(new_n544), .A4(new_n709), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n749), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT94), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n744), .A2(new_n747), .B1(new_n737), .B2(new_n736), .ZN(new_n757));
  AOI21_X1  g0557(.A(KEYINPUT93), .B1(new_n744), .B2(new_n747), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n744), .A2(KEYINPUT93), .A3(new_n747), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n709), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n756), .B1(new_n761), .B2(KEYINPUT31), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT93), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n748), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n746), .A2(new_n764), .A3(new_n760), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(new_n698), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n766), .A2(KEYINPUT94), .A3(new_n735), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n762), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n755), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G330), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n734), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n722), .B1(new_n772), .B2(G1), .ZN(G364));
  NAND2_X1  g0573(.A1(new_n708), .A2(G330), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(KEYINPUT98), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT98), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n708), .A2(new_n776), .A3(G330), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n363), .A2(G13), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n255), .B1(new_n779), .B2(G45), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n719), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n778), .B(new_n783), .C1(G330), .C2(new_n708), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n269), .B1(G20), .B2(new_n348), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n363), .A2(G190), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n787), .A2(G179), .A3(new_n309), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n363), .A2(new_n344), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n273), .A2(G200), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n788), .A2(G283), .B1(new_n792), .B2(G322), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n273), .A2(new_n309), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n786), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(KEYINPUT33), .B(G317), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G179), .A2(G200), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n786), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n796), .A2(new_n797), .B1(new_n800), .B2(G329), .ZN(new_n801));
  INV_X1    g0601(.A(new_n789), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n802), .A2(new_n309), .A3(G179), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n338), .B1(new_n804), .B2(new_n580), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n793), .B(new_n801), .C1(new_n805), .C2(KEYINPUT104), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n798), .A2(G190), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G20), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(G294), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n794), .A2(new_n789), .ZN(new_n811));
  INV_X1    g0611(.A(G326), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n809), .A2(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(G311), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n786), .A2(new_n790), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n813), .A2(KEYINPUT102), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(KEYINPUT102), .B2(new_n813), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT103), .Z(new_n818));
  AOI211_X1 g0618(.A(new_n806), .B(new_n818), .C1(KEYINPUT104), .C2(new_n805), .ZN(new_n819));
  INV_X1    g0619(.A(new_n811), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G50), .A2(new_n820), .B1(new_n796), .B2(G68), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n264), .B2(new_n815), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n803), .A2(G87), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n338), .B1(new_n792), .B2(G58), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n788), .A2(G107), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n799), .A2(new_n361), .ZN(new_n827));
  XOR2_X1   g0627(.A(KEYINPUT101), .B(KEYINPUT32), .Z(new_n828));
  XNOR2_X1  g0628(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n809), .A2(new_n546), .ZN(new_n830));
  NOR4_X1   g0630(.A1(new_n822), .A2(new_n826), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n785), .B1(new_n819), .B2(new_n831), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n782), .A2(KEYINPUT99), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n782), .A2(KEYINPUT99), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(G13), .A2(G33), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n837), .A2(G20), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n209), .A2(G355), .A3(new_n261), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n718), .A2(new_n261), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(G45), .B2(new_n225), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n250), .A2(new_n523), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n839), .B1(G116), .B2(new_n209), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n838), .B(new_n785), .C1(new_n843), .C2(KEYINPUT100), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n843), .A2(KEYINPUT100), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n835), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n838), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n832), .B(new_n846), .C1(new_n708), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n784), .A2(new_n848), .ZN(G396));
  NAND2_X1  g0649(.A1(new_n688), .A2(new_n690), .ZN(new_n850));
  INV_X1    g0650(.A(new_n672), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n709), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n709), .B1(new_n324), .B2(new_n331), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n324), .A2(new_n331), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n347), .A2(new_n854), .B1(new_n855), .B2(new_n350), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n351), .A2(new_n709), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n853), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT106), .ZN(new_n860));
  INV_X1    g0660(.A(new_n858), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n852), .A2(new_n861), .A3(new_n709), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n853), .A2(KEYINPUT106), .A3(new_n858), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(G330), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n755), .B2(new_n768), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n863), .A2(new_n770), .A3(new_n864), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n868), .A2(new_n783), .A3(new_n869), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n788), .A2(G87), .B1(G311), .B2(new_n800), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n871), .B(KEYINPUT105), .Z(new_n872));
  INV_X1    g0672(.A(new_n815), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n820), .A2(G303), .B1(new_n873), .B2(G116), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n803), .A2(G107), .B1(G283), .B2(new_n796), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n261), .B(new_n830), .C1(G294), .C2(new_n792), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n872), .A2(new_n874), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(G150), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n795), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(G143), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n791), .A2(new_n880), .B1(new_n815), .B2(new_n361), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n879), .B(new_n881), .C1(G137), .C2(new_n820), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT34), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n261), .B1(new_n804), .B2(new_n202), .ZN(new_n884));
  INV_X1    g0684(.A(new_n788), .ZN(new_n885));
  INV_X1    g0685(.A(G132), .ZN(new_n886));
  OAI22_X1  g0686(.A1(new_n885), .A2(new_n246), .B1(new_n799), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n883), .B(new_n888), .C1(new_n289), .C2(new_n809), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n882), .A2(KEYINPUT34), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n877), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n785), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n785), .A2(new_n836), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n835), .B1(new_n264), .B2(new_n893), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n892), .B(new_n894), .C1(new_n861), .C2(new_n837), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n870), .A2(new_n895), .ZN(G384));
  INV_X1    g0696(.A(new_n551), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n897), .A2(KEYINPUT35), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(KEYINPUT35), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n269), .A2(new_n363), .A3(new_n216), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  XOR2_X1   g0701(.A(new_n901), .B(KEYINPUT107), .Z(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(KEYINPUT36), .ZN(new_n903));
  OR3_X1    g0703(.A1(new_n225), .A2(new_n264), .A3(new_n358), .ZN(new_n904));
  AOI211_X1 g0704(.A(new_n255), .B(G13), .C1(new_n904), .C2(new_n245), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n696), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n657), .A2(new_n907), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n461), .A2(new_n468), .A3(new_n456), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT77), .B1(new_n472), .B2(new_n473), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n431), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT108), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n475), .A2(KEYINPUT108), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n431), .A2(new_n698), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n454), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n909), .A2(new_n910), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n918), .A2(new_n915), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n862), .A2(new_n857), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT38), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT37), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n368), .A2(new_n372), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT16), .B1(new_n924), .B2(new_n403), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n402), .B1(new_n407), .B2(new_n925), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n390), .A2(new_n413), .B1(new_n926), .B2(new_n907), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n399), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n923), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n409), .A2(new_n399), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n409), .A2(new_n907), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n930), .A2(new_n931), .A3(new_n923), .A4(new_n414), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n924), .A2(new_n403), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT16), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n357), .B1(new_n937), .B2(new_n374), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n938), .A2(new_n696), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n657), .B2(new_n652), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n922), .B1(new_n934), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n414), .B1(new_n938), .B2(new_n696), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n938), .A2(new_n400), .ZN(new_n944));
  OAI21_X1  g0744(.A(KEYINPUT37), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n932), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n419), .A2(new_n939), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n946), .A2(new_n947), .A3(KEYINPUT38), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n942), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n908), .B1(new_n921), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n475), .A2(KEYINPUT108), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n912), .B(new_n432), .C1(new_n469), .C2(new_n474), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n709), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT109), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n946), .A2(new_n947), .A3(KEYINPUT38), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT38), .B1(new_n946), .B2(new_n947), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n955), .B(KEYINPUT39), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n930), .A2(new_n931), .A3(new_n414), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(KEYINPUT37), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n932), .ZN(new_n961));
  INV_X1    g0761(.A(new_n931), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n419), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n922), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT39), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n965), .A2(new_n966), .A3(new_n948), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n958), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n955), .B1(new_n949), .B2(KEYINPUT39), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n954), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AND3_X1   g0770(.A1(new_n950), .A2(new_n970), .A3(KEYINPUT110), .ZN(new_n971));
  AOI21_X1  g0771(.A(KEYINPUT110), .B1(new_n950), .B2(new_n970), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n725), .A2(new_n476), .A3(new_n727), .A4(new_n733), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n660), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n973), .B(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n752), .A2(new_n754), .ZN(new_n977));
  AOI211_X1 g0777(.A(new_n735), .B(new_n709), .C1(new_n759), .C2(new_n760), .ZN(new_n978));
  AOI21_X1  g0778(.A(KEYINPUT31), .B1(new_n765), .B2(new_n698), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n858), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n454), .A2(new_n915), .ZN(new_n982));
  NOR3_X1   g0782(.A1(new_n951), .A2(new_n952), .A3(new_n982), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n949), .B(new_n981), .C1(new_n983), .C2(new_n919), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT40), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n917), .A2(new_n920), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n965), .A2(new_n948), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n987), .A2(KEYINPUT40), .A3(new_n988), .A4(new_n981), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n977), .A2(new_n980), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n476), .A2(new_n991), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n990), .A2(new_n992), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n993), .A2(G330), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n976), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n255), .B2(new_n779), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n976), .A2(new_n995), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n906), .B1(new_n997), .B2(new_n998), .ZN(G367));
  INV_X1    g0799(.A(new_n835), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n840), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n235), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n785), .A2(new_n838), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n209), .B2(new_n328), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1000), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n804), .A2(new_n289), .B1(new_n811), .B2(new_n880), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n338), .B(new_n1006), .C1(G150), .C2(new_n792), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n788), .A2(G77), .B1(G137), .B2(new_n800), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G159), .A2(new_n796), .B1(new_n873), .B2(G50), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n808), .A2(G68), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n261), .B1(new_n788), .B2(G97), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n820), .A2(G311), .B1(new_n800), .B2(G317), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1012), .B(new_n1013), .C1(new_n333), .C2(new_n809), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n803), .A2(G116), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT46), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G294), .A2(new_n796), .B1(new_n792), .B2(G303), .ZN(new_n1017));
  INV_X1    g0817(.A(G283), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1016), .B(new_n1017), .C1(new_n1018), .C2(new_n815), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1011), .B1(new_n1014), .B2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT47), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1005), .B1(new_n1021), .B2(new_n785), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT114), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n709), .B1(new_n627), .B2(new_n645), .ZN(new_n1024));
  MUX2_X1   g0824(.A(new_n728), .B(new_n643), .S(new_n1024), .Z(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n838), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT112), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT111), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n554), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n684), .B1(new_n1030), .B2(new_n709), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n669), .A2(new_n698), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n716), .A2(new_n714), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT44), .Z(new_n1037));
  NOR2_X1   g0837(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT45), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1037), .A2(new_n713), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n713), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1029), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n1029), .B2(new_n1042), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n716), .B1(new_n712), .B2(new_n715), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n774), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n778), .B2(new_n1045), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n772), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1028), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1042), .A2(new_n1029), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1042), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n1040), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1050), .B1(new_n1052), .B2(new_n1029), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1053), .A2(KEYINPUT112), .A3(new_n772), .A4(new_n1047), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1049), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n772), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n719), .B(KEYINPUT41), .Z(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1056), .A2(KEYINPUT113), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT113), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n771), .B1(new_n1049), .B2(new_n1054), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1060), .B1(new_n1061), .B2(new_n1057), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n781), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1033), .A2(new_n544), .A3(new_n715), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n572), .B1(new_n676), .B2(new_n679), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n1064), .A2(KEYINPUT42), .B1(new_n709), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(KEYINPUT42), .B2(new_n1064), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT43), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1067), .B1(new_n1068), .B2(new_n1025), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1025), .A2(new_n1068), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1069), .B(new_n1070), .Z(new_n1071));
  OR2_X1    g0871(.A1(new_n713), .A2(new_n1034), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1071), .B(new_n1072), .Z(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1027), .B1(new_n1063), .B2(new_n1074), .ZN(G387));
  NAND3_X1  g0875(.A1(new_n710), .A2(new_n711), .A3(new_n838), .ZN(new_n1076));
  OR3_X1    g0876(.A1(new_n240), .A2(new_n523), .A3(new_n261), .ZN(new_n1077));
  OAI21_X1  g0877(.A(KEYINPUT50), .B1(new_n286), .B2(G50), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1078), .B(new_n523), .C1(new_n246), .C2(new_n264), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n286), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n338), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1081), .A2(new_n393), .A3(new_n216), .A4(new_n616), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n718), .B1(new_n1077), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1003), .B1(new_n333), .B2(new_n209), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1000), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n803), .A2(G77), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n246), .B2(new_n815), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n338), .B(new_n1087), .C1(G97), .C2(new_n788), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n808), .A2(new_n327), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n354), .A2(new_n796), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n791), .A2(new_n202), .B1(new_n799), .B2(new_n878), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(G159), .B2(new_n820), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .A4(new_n1092), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n804), .A2(new_n810), .B1(new_n1018), .B2(new_n809), .ZN(new_n1094));
  XOR2_X1   g0894(.A(KEYINPUT115), .B(G322), .Z(new_n1095));
  INV_X1    g0895(.A(G317), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n811), .A2(new_n1095), .B1(new_n791), .B2(new_n1096), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n795), .A2(new_n814), .B1(new_n815), .B2(new_n580), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1094), .B1(new_n1099), .B2(KEYINPUT48), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1099), .A2(KEYINPUT48), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1100), .A2(KEYINPUT49), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n261), .B1(new_n800), .B2(G326), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1102), .B(new_n1103), .C1(new_n216), .C2(new_n885), .ZN(new_n1104));
  AOI21_X1  g0904(.A(KEYINPUT49), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1093), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1085), .B1(new_n1106), .B2(new_n785), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1047), .A2(new_n781), .B1(new_n1076), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1048), .A2(KEYINPUT116), .A3(new_n719), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n1047), .A2(new_n772), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(KEYINPUT116), .B1(new_n1048), .B2(new_n719), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1108), .B1(new_n1111), .B2(new_n1112), .ZN(G393));
  INV_X1    g0913(.A(new_n719), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n1048), .B2(new_n1052), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1055), .A2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1001), .A2(new_n244), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1003), .B1(new_n546), .B2(new_n209), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1000), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n795), .A2(new_n580), .B1(new_n815), .B2(new_n810), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(G116), .B2(new_n808), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT117), .Z(new_n1122));
  OAI22_X1  g0922(.A1(new_n811), .A2(new_n1096), .B1(new_n791), .B2(new_n814), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT52), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1095), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n803), .A2(G283), .B1(new_n1125), .B2(new_n800), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1124), .A2(new_n338), .A3(new_n825), .A4(new_n1126), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n804), .A2(new_n246), .B1(new_n799), .B2(new_n880), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n808), .A2(G77), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n261), .B(new_n1129), .C1(new_n885), .C2(new_n393), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n795), .A2(new_n202), .B1(new_n815), .B2(new_n286), .ZN(new_n1131));
  OR3_X1    g0931(.A1(new_n1128), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n811), .A2(new_n878), .B1(new_n791), .B2(new_n361), .ZN(new_n1133));
  XOR2_X1   g0933(.A(new_n1133), .B(KEYINPUT51), .Z(new_n1134));
  OAI22_X1  g0934(.A1(new_n1122), .A2(new_n1127), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  XOR2_X1   g0935(.A(new_n1135), .B(KEYINPUT118), .Z(new_n1136));
  AOI21_X1  g0936(.A(new_n1119), .B1(new_n1136), .B2(new_n785), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n1033), .B2(new_n847), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n1052), .B2(new_n780), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1116), .A2(new_n1140), .ZN(G390));
  INV_X1    g0941(.A(new_n893), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1000), .B1(new_n354), .B2(new_n1142), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n788), .A2(G68), .B1(new_n820), .B2(G283), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1144), .A2(new_n338), .A3(new_n823), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(G107), .A2(new_n796), .B1(new_n792), .B2(G116), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G97), .A2(new_n873), .B1(new_n800), .B2(G294), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1145), .A2(new_n1129), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n804), .A2(new_n878), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT53), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1149), .A2(new_n1150), .B1(G159), .B2(new_n808), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(KEYINPUT54), .B(G143), .ZN(new_n1152));
  INV_X1    g0952(.A(G125), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n815), .A2(new_n1152), .B1(new_n799), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1151), .B(new_n1155), .C1(new_n1150), .C2(new_n1149), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n261), .B1(new_n885), .B2(new_n202), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT120), .ZN(new_n1158));
  OR2_X1    g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1160));
  INV_X1    g0960(.A(G128), .ZN(new_n1161));
  INV_X1    g0961(.A(G137), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n811), .A2(new_n1161), .B1(new_n795), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(G132), .B2(new_n792), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1159), .A2(new_n1160), .A3(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1148), .B1(new_n1156), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1143), .B1(new_n1166), .B2(new_n785), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n966), .B1(new_n942), .B2(new_n948), .ZN(new_n1168));
  AOI21_X1  g0968(.A(KEYINPUT38), .B1(new_n961), .B2(new_n963), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n956), .A2(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1168), .A2(new_n955), .B1(new_n1170), .B2(new_n966), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n949), .A2(KEYINPUT39), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(KEYINPUT109), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1167), .B1(new_n1174), .B2(new_n837), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n732), .A2(new_n709), .A3(new_n856), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n857), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n987), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1178), .A2(new_n953), .A3(new_n988), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n987), .A2(new_n867), .A3(new_n861), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n862), .A2(new_n857), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n954), .B1(new_n1181), .B2(new_n987), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1179), .B(new_n1180), .C1(new_n1174), .C2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n953), .A2(new_n988), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n987), .B2(new_n1177), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n862), .A2(new_n857), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n917), .A2(new_n920), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n953), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n968), .A2(new_n969), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1185), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n987), .A2(G330), .A3(new_n981), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1183), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1175), .B1(new_n1192), .B2(new_n780), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n476), .A2(G330), .A3(new_n991), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n974), .A2(new_n660), .A3(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT119), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n974), .A2(new_n660), .A3(KEYINPUT119), .A4(new_n1194), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n991), .A2(G330), .A3(new_n861), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1177), .B1(new_n1187), .B2(new_n1199), .ZN(new_n1200));
  AND2_X1   g1000(.A1(new_n1200), .A2(new_n1180), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1187), .B1(new_n770), .B2(new_n858), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1186), .B1(new_n1202), .B2(new_n1191), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1197), .B(new_n1198), .C1(new_n1201), .C2(new_n1203), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1204), .A2(new_n1192), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1114), .B1(new_n1204), .B2(new_n1192), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1193), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(G378));
  NAND3_X1  g1008(.A1(new_n986), .A2(G330), .A3(new_n989), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n306), .A2(new_n696), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n318), .B(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1211), .B(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1209), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1213), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n986), .A2(new_n1215), .A3(G330), .A4(new_n989), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n973), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(KEYINPUT122), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT123), .ZN(new_n1220));
  AND2_X1   g1020(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n950), .A2(new_n970), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT110), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n950), .A2(new_n970), .A3(KEYINPUT110), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1220), .B1(new_n1221), .B2(new_n1226), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1214), .B(new_n1216), .C1(new_n971), .C2(new_n972), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1228), .A2(KEYINPUT123), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1219), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(KEYINPUT123), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT122), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n973), .B2(new_n1217), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1226), .A2(new_n1220), .A3(new_n1216), .A4(new_n1214), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1231), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1230), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1213), .A2(new_n836), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n782), .B1(new_n1142), .B2(G50), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n811), .A2(new_n1153), .B1(new_n795), .B2(new_n886), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n792), .A2(G128), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n1240), .B1(new_n815), .B2(new_n1162), .C1(new_n804), .C2(new_n1152), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n1239), .B(new_n1241), .C1(G150), .C2(new_n808), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT59), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n788), .A2(G159), .ZN(new_n1246));
  AOI211_X1 g1046(.A(G33), .B(G41), .C1(new_n800), .C2(G124), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n796), .A2(G97), .B1(new_n873), .B2(new_n327), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT121), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(G116), .A2(new_n820), .B1(new_n792), .B2(G107), .ZN(new_n1251));
  OAI221_X1 g1051(.A(new_n1251), .B1(new_n1018), .B2(new_n799), .C1(new_n289), .C2(new_n885), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1086), .A2(new_n253), .A3(new_n338), .A4(new_n1010), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1250), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(KEYINPUT58), .ZN(new_n1255));
  OR2_X1    g1055(.A1(new_n1254), .A2(KEYINPUT58), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n253), .B1(new_n335), .B2(new_n252), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n202), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1248), .A2(new_n1255), .A3(new_n1256), .A4(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1238), .B1(new_n1259), .B2(new_n785), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1236), .A2(new_n781), .B1(new_n1237), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1202), .A2(new_n1191), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1262), .A2(new_n1181), .B1(new_n1180), .B2(new_n1200), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1197), .B(new_n1198), .C1(new_n1192), .C2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT57), .B1(new_n1236), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1218), .A2(new_n1228), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1266), .A2(KEYINPUT57), .A3(new_n1264), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n719), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1261), .B1(new_n1265), .B2(new_n1268), .ZN(G375));
  NAND2_X1  g1069(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1263), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1271), .A2(new_n1058), .A3(new_n1204), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n835), .B1(new_n246), .B2(new_n893), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n785), .ZN(new_n1274));
  OAI22_X1  g1074(.A1(new_n811), .A2(new_n886), .B1(new_n791), .B2(new_n1162), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n261), .B1(new_n885), .B2(new_n289), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n1275), .B(new_n1276), .C1(G50), .C2(new_n808), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n815), .A2(new_n878), .ZN(new_n1278));
  OAI22_X1  g1078(.A1(new_n795), .A2(new_n1152), .B1(new_n799), .B2(new_n1161), .ZN(new_n1279));
  AOI211_X1 g1079(.A(new_n1278), .B(new_n1279), .C1(G159), .C2(new_n803), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(G116), .A2(new_n796), .B1(new_n792), .B2(G283), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n261), .B1(new_n788), .B2(G77), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1281), .A2(new_n1282), .A3(new_n1089), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n811), .A2(new_n810), .ZN(new_n1284));
  OAI22_X1  g1084(.A1(new_n815), .A2(new_n333), .B1(new_n799), .B2(new_n580), .ZN(new_n1285));
  AOI211_X1 g1085(.A(new_n1284), .B(new_n1285), .C1(G97), .C2(new_n803), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(new_n1277), .A2(new_n1280), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1287));
  OAI221_X1 g1087(.A(new_n1273), .B1(new_n1274), .B2(new_n1287), .C1(new_n987), .C2(new_n837), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n780), .B(KEYINPUT124), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1288), .B1(new_n1263), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1272), .A2(new_n1291), .ZN(G381));
  OR2_X1    g1092(.A1(G375), .A2(G378), .ZN(new_n1293));
  INV_X1    g1093(.A(G396), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1294), .B(new_n1108), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1295));
  OR4_X1    g1095(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1295), .ZN(new_n1296));
  OR3_X1    g1096(.A1(new_n1293), .A2(G387), .A3(new_n1296), .ZN(G407));
  OAI211_X1 g1097(.A(G407), .B(G213), .C1(G343), .C2(new_n1293), .ZN(G409));
  NAND3_X1  g1098(.A1(new_n1270), .A2(KEYINPUT60), .A3(new_n1263), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1299), .A2(new_n719), .ZN(new_n1300));
  OAI21_X1  g1100(.A(KEYINPUT60), .B1(new_n1270), .B2(new_n1263), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1271), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1300), .A2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(G384), .B1(new_n1303), .B2(new_n1291), .ZN(new_n1304));
  INV_X1    g1104(.A(G384), .ZN(new_n1305));
  AOI211_X1 g1105(.A(new_n1305), .B(new_n1290), .C1(new_n1300), .C2(new_n1302), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n697), .A2(G213), .A3(G2897), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1304), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1307), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1299), .A2(new_n719), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1310), .B1(new_n1271), .B2(new_n1301), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1305), .B1(new_n1311), .B2(new_n1290), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1303), .A2(G384), .A3(new_n1291), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1309), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1308), .A2(new_n1314), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1231), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1316));
  AOI22_X1  g1116(.A1(new_n1231), .A2(new_n1234), .B1(KEYINPUT122), .B2(new_n1218), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1264), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT57), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1268), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n781), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1237), .A2(new_n1260), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(G378), .B1(new_n1320), .B2(new_n1323), .ZN(new_n1324));
  OAI211_X1 g1124(.A(new_n1058), .B(new_n1264), .C1(new_n1316), .C2(new_n1317), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1289), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1266), .A2(new_n1326), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1207), .A2(new_n1322), .A3(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1325), .A2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n697), .A2(G213), .ZN(new_n1330));
  AND2_X1   g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1315), .B1(new_n1324), .B2(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(KEYINPUT127), .B1(new_n1332), .B2(KEYINPUT61), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT127), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT61), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1336), .B1(G375), .B2(G378), .ZN(new_n1337));
  OAI211_X1 g1137(.A(new_n1334), .B(new_n1335), .C1(new_n1337), .C2(new_n1315), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1324), .A2(new_n1331), .A3(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(KEYINPUT62), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT62), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1337), .A2(new_n1342), .A3(new_n1339), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1333), .A2(new_n1338), .A3(new_n1341), .A4(new_n1343), .ZN(new_n1344));
  AND2_X1   g1144(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1073), .B1(new_n1345), .B2(new_n781), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(G393), .A2(G396), .ZN(new_n1347));
  AND3_X1   g1147(.A1(G390), .A2(new_n1347), .A3(new_n1295), .ZN(new_n1348));
  AOI21_X1  g1148(.A(G390), .B1(new_n1295), .B2(new_n1347), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1346), .A2(new_n1350), .A3(new_n1027), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1349), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(G390), .A2(new_n1347), .A3(new_n1295), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1352), .A2(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1354), .A2(G387), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1351), .A2(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1344), .A2(new_n1356), .ZN(new_n1357));
  AND2_X1   g1157(.A1(new_n1315), .A2(KEYINPUT126), .ZN(new_n1358));
  NOR2_X1   g1158(.A1(new_n1315), .A2(KEYINPUT126), .ZN(new_n1359));
  OR3_X1    g1159(.A1(new_n1358), .A2(new_n1337), .A3(new_n1359), .ZN(new_n1360));
  NOR2_X1   g1160(.A1(new_n1356), .A2(KEYINPUT61), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1340), .A2(KEYINPUT125), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1362), .A2(KEYINPUT63), .ZN(new_n1363));
  INV_X1    g1163(.A(KEYINPUT63), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1340), .A2(KEYINPUT125), .A3(new_n1364), .ZN(new_n1365));
  NAND4_X1  g1165(.A1(new_n1360), .A2(new_n1361), .A3(new_n1363), .A4(new_n1365), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1357), .A2(new_n1366), .ZN(G405));
  NAND2_X1  g1167(.A1(new_n1293), .A2(new_n1324), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1368), .A2(new_n1339), .ZN(new_n1369));
  INV_X1    g1169(.A(new_n1356), .ZN(new_n1370));
  OAI211_X1 g1170(.A(new_n1293), .B(new_n1324), .C1(new_n1304), .C2(new_n1306), .ZN(new_n1371));
  AND3_X1   g1171(.A1(new_n1369), .A2(new_n1370), .A3(new_n1371), .ZN(new_n1372));
  AOI21_X1  g1172(.A(new_n1370), .B1(new_n1369), .B2(new_n1371), .ZN(new_n1373));
  NOR2_X1   g1173(.A1(new_n1372), .A2(new_n1373), .ZN(G402));
endmodule


