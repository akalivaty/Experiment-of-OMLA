//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 0 0 0 0 1 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n819, new_n820, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921;
  INV_X1    g000(.A(KEYINPUT6), .ZN(new_n202));
  XNOR2_X1  g001(.A(G1gat), .B(G29gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT0), .ZN(new_n204));
  XNOR2_X1  g003(.A(G57gat), .B(G85gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  NAND2_X1  g005(.A1(G225gat), .A2(G233gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G127gat), .B(G134gat), .ZN(new_n209));
  INV_X1    g008(.A(G113gat), .ZN(new_n210));
  INV_X1    g009(.A(G120gat), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT1), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  OR2_X1    g012(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n211), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AND2_X1   g015(.A1(G113gat), .A2(G120gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(G113gat), .A2(G120gat), .ZN(new_n218));
  NOR3_X1   g017(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT1), .ZN(new_n219));
  OAI22_X1  g018(.A1(new_n213), .A2(new_n216), .B1(new_n219), .B2(new_n209), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT2), .ZN(new_n223));
  INV_X1    g022(.A(G141gat), .ZN(new_n224));
  INV_X1    g023(.A(G148gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G141gat), .A2(G148gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n223), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT79), .ZN(new_n229));
  XNOR2_X1  g028(.A(G155gat), .B(G162gat), .ZN(new_n230));
  AND3_X1   g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n230), .B1(new_n228), .B2(new_n229), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n221), .B1(new_n233), .B2(KEYINPUT3), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n228), .A2(new_n229), .ZN(new_n235));
  INV_X1    g034(.A(new_n230), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n208), .B1(new_n234), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT80), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n243), .B1(new_n233), .B2(new_n220), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT4), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n239), .A2(new_n221), .A3(KEYINPUT80), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n233), .A2(new_n220), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT4), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n242), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT81), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n251), .B1(new_n233), .B2(new_n220), .ZN(new_n252));
  AND4_X1   g051(.A1(new_n251), .A2(new_n220), .A3(new_n237), .A4(new_n238), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n244), .A2(new_n246), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n208), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n250), .A2(new_n256), .A3(KEYINPUT5), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n244), .A2(KEYINPUT4), .A3(new_n246), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT82), .B1(new_n248), .B2(new_n245), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT5), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n244), .A2(new_n246), .A3(KEYINPUT82), .A4(KEYINPUT4), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n260), .A2(new_n261), .A3(new_n242), .A4(new_n262), .ZN(new_n263));
  AOI211_X1 g062(.A(new_n202), .B(new_n206), .C1(new_n257), .C2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT89), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n257), .A2(new_n263), .ZN(new_n267));
  INV_X1    g066(.A(new_n206), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT6), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n257), .A2(new_n206), .A3(new_n263), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n264), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n266), .B1(new_n271), .B2(KEYINPUT89), .ZN(new_n272));
  XOR2_X1   g071(.A(KEYINPUT90), .B(KEYINPUT35), .Z(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  OR2_X1    g074(.A1(G183gat), .A2(G190gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n276), .B(new_n277), .C1(new_n278), .C2(KEYINPUT64), .ZN(new_n279));
  NAND2_X1  g078(.A1(G183gat), .A2(G190gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT24), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT64), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT65), .B1(new_n279), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286));
  AND2_X1   g085(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n286), .B1(new_n287), .B2(G190gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n282), .A2(new_n283), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT65), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n278), .A2(KEYINPUT64), .ZN(new_n291));
  NAND4_X1  g090(.A1(new_n288), .A2(new_n289), .A3(new_n290), .A4(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT23), .ZN(new_n294));
  NAND2_X1  g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT23), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n296), .B1(G169gat), .B2(G176gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n294), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n285), .A2(new_n292), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT25), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n294), .A2(KEYINPUT25), .A3(new_n297), .A4(new_n295), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n281), .A2(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n304), .B1(KEYINPUT66), .B2(new_n281), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n303), .B1(new_n305), .B2(new_n288), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(KEYINPUT27), .B(G183gat), .ZN(new_n309));
  INV_X1    g108(.A(G190gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT28), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(KEYINPUT67), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(KEYINPUT67), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n309), .A2(new_n310), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n293), .A2(KEYINPUT26), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(new_n280), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT26), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n295), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n320), .A2(new_n293), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G226gat), .A2(G233gat), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G197gat), .B(G204gat), .ZN(new_n328));
  INV_X1    g127(.A(G211gat), .ZN(new_n329));
  INV_X1    g128(.A(G218gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n328), .B1(KEYINPUT22), .B2(new_n331), .ZN(new_n332));
  XOR2_X1   g131(.A(G211gat), .B(G218gat), .Z(new_n333));
  XNOR2_X1  g132(.A(new_n332), .B(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n327), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT29), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT75), .B1(new_n308), .B2(new_n323), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n306), .B1(new_n300), .B2(new_n301), .ZN(new_n339));
  AOI211_X1 g138(.A(new_n321), .B(new_n318), .C1(new_n313), .C2(new_n315), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n341));
  NOR3_X1   g140(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n337), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT76), .B1(new_n343), .B2(new_n325), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n341), .B1(new_n339), .B2(new_n340), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n288), .A2(new_n289), .A3(new_n291), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n298), .B1(new_n346), .B2(KEYINPUT65), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT25), .B1(new_n347), .B2(new_n292), .ZN(new_n348));
  OAI211_X1 g147(.A(KEYINPUT75), .B(new_n323), .C1(new_n348), .C2(new_n306), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT29), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT76), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n350), .A2(new_n351), .A3(new_n326), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n336), .B1(new_n344), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n345), .A2(new_n349), .A3(new_n326), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n324), .A2(new_n337), .A3(new_n325), .ZN(new_n355));
  INV_X1    g154(.A(new_n334), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G8gat), .B(G36gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(G64gat), .B(G92gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n361), .B(new_n362), .Z(new_n363));
  NAND4_X1  g162(.A1(new_n353), .A2(KEYINPUT30), .A3(new_n358), .A4(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n363), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n343), .A2(KEYINPUT76), .A3(new_n325), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n351), .B1(new_n350), .B2(new_n326), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n335), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n365), .B1(new_n368), .B2(new_n357), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n364), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n366), .A2(new_n367), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n357), .B1(new_n371), .B2(new_n336), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT30), .B1(new_n372), .B2(new_n363), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT85), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n353), .A2(new_n358), .A3(new_n363), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT30), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT85), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n377), .A2(new_n378), .A3(new_n369), .A4(new_n364), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n275), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT72), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n221), .B1(new_n339), .B2(new_n340), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n220), .B(new_n323), .C1(new_n348), .C2(new_n306), .ZN(new_n383));
  NAND2_X1  g182(.A1(G227gat), .A2(G233gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n382), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT32), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT33), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G15gat), .B(G43gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(KEYINPUT69), .ZN(new_n391));
  XNOR2_X1  g190(.A(G71gat), .B(G99gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT70), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n387), .B1(new_n393), .B2(KEYINPUT33), .ZN(new_n396));
  AND3_X1   g195(.A1(new_n386), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n395), .B1(new_n386), .B2(new_n396), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n394), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n383), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n384), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT34), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n402), .B1(new_n384), .B2(KEYINPUT71), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n400), .B(new_n384), .C1(KEYINPUT71), .C2(new_n402), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n381), .B1(new_n399), .B2(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n404), .A2(new_n405), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n386), .A2(new_n396), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT70), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n386), .A2(new_n395), .A3(new_n396), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n408), .A2(new_n412), .A3(KEYINPUT72), .A4(new_n394), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n407), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT73), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT73), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n407), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n399), .A2(new_n406), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n415), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n334), .A2(new_n337), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n239), .B1(new_n420), .B2(new_n240), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n334), .B1(new_n241), .B2(new_n337), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(G228gat), .A2(G233gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(G22gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n423), .B(new_n424), .ZN(new_n427));
  INV_X1    g226(.A(G22gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n426), .A2(new_n429), .A3(KEYINPUT83), .ZN(new_n430));
  XNOR2_X1  g229(.A(G78gat), .B(G106gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(KEYINPUT31), .B(G50gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n427), .A2(new_n428), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT83), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n430), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n426), .A2(new_n429), .A3(new_n433), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT84), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n426), .A2(new_n429), .A3(KEYINPUT84), .A4(new_n433), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n437), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n419), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n437), .A2(new_n440), .A3(new_n441), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n370), .A2(new_n373), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n267), .A2(new_n268), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n446), .A2(new_n202), .A3(new_n270), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n265), .ZN(new_n448));
  INV_X1    g247(.A(new_n418), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n449), .B1(new_n407), .B2(new_n413), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n444), .A2(new_n445), .A3(new_n448), .A4(new_n450), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n380), .A2(new_n443), .B1(new_n451), .B2(KEYINPUT35), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n444), .B1(new_n445), .B2(new_n448), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT38), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n327), .A2(new_n356), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n455), .B1(new_n366), .B2(new_n367), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n354), .A2(new_n334), .A3(new_n355), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT37), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n454), .B(new_n365), .C1(new_n456), .C2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT37), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n353), .A2(new_n460), .A3(new_n358), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT88), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n372), .A2(KEYINPUT88), .A3(new_n460), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n459), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n375), .B(new_n266), .C1(new_n271), .C2(KEYINPUT89), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n353), .A2(new_n358), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n363), .B1(new_n468), .B2(KEYINPUT37), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT88), .B1(new_n372), .B2(new_n460), .ZN(new_n470));
  NOR4_X1   g269(.A1(new_n368), .A2(new_n462), .A3(KEYINPUT37), .A4(new_n357), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT38), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n442), .B1(new_n467), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT87), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n234), .A2(new_n241), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n260), .A2(new_n476), .A3(new_n262), .ZN(new_n477));
  XOR2_X1   g276(.A(KEYINPUT86), .B(KEYINPUT39), .Z(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n208), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n206), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n220), .A2(new_n237), .A3(new_n238), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n481), .B(KEYINPUT81), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n482), .A2(new_n244), .A3(new_n246), .A4(new_n207), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT39), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n484), .B1(new_n208), .B2(new_n477), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n475), .B1(new_n480), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT40), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT40), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n475), .B(new_n488), .C1(new_n480), .C2(new_n485), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n487), .A2(new_n446), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n374), .A2(new_n490), .A3(new_n379), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n453), .B1(new_n474), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT36), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n419), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT74), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n449), .B1(new_n414), .B2(KEYINPUT73), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT36), .B1(new_n496), .B2(new_n417), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT74), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n450), .A2(KEYINPUT36), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n495), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n452), .B1(new_n492), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(KEYINPUT91), .B(G29gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(G36gat), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT14), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(G29gat), .B2(G36gat), .ZN(new_n506));
  OR3_X1    g305(.A1(new_n505), .A2(G29gat), .A3(G36gat), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n504), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT15), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n504), .A2(KEYINPUT15), .A3(new_n506), .A4(new_n507), .ZN(new_n511));
  XNOR2_X1  g310(.A(G43gat), .B(G50gat), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n511), .A2(new_n512), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G15gat), .B(G22gat), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT16), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n517), .B1(new_n518), .B2(G1gat), .ZN(new_n519));
  INV_X1    g318(.A(G8gat), .ZN(new_n520));
  OAI221_X1 g319(.A(new_n519), .B1(KEYINPUT92), .B2(new_n520), .C1(G1gat), .C2(new_n517), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(KEYINPUT92), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n521), .B(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n516), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n521), .B(new_n522), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n515), .A2(KEYINPUT17), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT17), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n513), .A2(new_n528), .A3(new_n514), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n526), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT93), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n525), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G229gat), .A2(G233gat), .ZN(new_n533));
  INV_X1    g332(.A(new_n529), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n528), .B1(new_n513), .B2(new_n514), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n524), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT93), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n532), .A2(new_n533), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT94), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n532), .A2(new_n537), .A3(KEYINPUT94), .A4(new_n533), .ZN(new_n541));
  XOR2_X1   g340(.A(KEYINPUT95), .B(KEYINPUT18), .Z(new_n542));
  NAND3_X1  g341(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G113gat), .B(G141gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(G197gat), .ZN(new_n545));
  XOR2_X1   g344(.A(KEYINPUT11), .B(G169gat), .Z(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT12), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n526), .B(new_n515), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n533), .B(KEYINPUT13), .Z(new_n550));
  AND2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n532), .A2(new_n533), .A3(new_n537), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n551), .B1(new_n552), .B2(KEYINPUT18), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n543), .A2(new_n548), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n548), .B1(new_n543), .B2(new_n553), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n502), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT9), .ZN(new_n558));
  XNOR2_X1  g357(.A(G57gat), .B(G64gat), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n558), .B1(new_n559), .B2(KEYINPUT97), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n560), .B1(KEYINPUT97), .B2(new_n559), .ZN(new_n561));
  NAND2_X1  g360(.A1(G71gat), .A2(G78gat), .ZN(new_n562));
  NOR2_X1   g361(.A1(G71gat), .A2(G78gat), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT96), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n565), .B1(new_n564), .B2(new_n563), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n568));
  AND2_X1   g367(.A1(new_n568), .A2(new_n562), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n569), .A2(new_n559), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT21), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(G127gat), .ZN(new_n576));
  XOR2_X1   g375(.A(G183gat), .B(G211gat), .Z(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n571), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n526), .B1(KEYINPUT21), .B2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT99), .ZN(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT98), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(G155gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n581), .B(new_n584), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n578), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n578), .A2(new_n585), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(G230gat), .ZN(new_n589));
  INV_X1    g388(.A(G233gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(KEYINPUT100), .A2(G85gat), .A3(G92gat), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT7), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n593), .ZN(new_n595));
  NAND2_X1  g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  INV_X1    g395(.A(G85gat), .ZN(new_n597));
  INV_X1    g396(.A(G92gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(KEYINPUT8), .A2(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n594), .A2(new_n595), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G99gat), .B(G106gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n579), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT10), .ZN(new_n604));
  INV_X1    g403(.A(new_n602), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n571), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n579), .A2(KEYINPUT10), .A3(new_n602), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n591), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n603), .A2(new_n606), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n609), .B1(new_n610), .B2(new_n591), .ZN(new_n611));
  XOR2_X1   g410(.A(G120gat), .B(G148gat), .Z(new_n612));
  XNOR2_X1  g411(.A(G176gat), .B(G204gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n611), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n602), .B1(new_n527), .B2(new_n529), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT41), .ZN(new_n621));
  NAND2_X1  g420(.A1(G232gat), .A2(G233gat), .ZN(new_n622));
  OAI22_X1  g421(.A1(new_n516), .A2(new_n605), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT101), .ZN(new_n624));
  XNOR2_X1  g423(.A(G190gat), .B(G218gat), .ZN(new_n625));
  OAI22_X1  g424(.A1(new_n620), .A2(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G134gat), .B(G162gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n624), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n622), .A2(new_n621), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n628), .A2(new_n632), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NOR3_X1   g435(.A1(new_n588), .A2(new_n619), .A3(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n557), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n271), .B(KEYINPUT104), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G1gat), .ZN(G1324gat));
  INV_X1    g440(.A(new_n638), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n374), .A2(new_n379), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT16), .B(G8gat), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n643), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n520), .B1(new_n638), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(KEYINPUT42), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n648), .B1(KEYINPUT42), .B2(new_n645), .ZN(G1325gat));
  OAI21_X1  g448(.A(G15gat), .B1(new_n642), .B2(new_n501), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n419), .A2(G15gat), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n650), .B1(new_n642), .B2(new_n651), .ZN(G1326gat));
  NAND2_X1  g451(.A1(new_n638), .A2(new_n442), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT105), .ZN(new_n654));
  XOR2_X1   g453(.A(KEYINPUT43), .B(G22gat), .Z(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(G1327gat));
  INV_X1    g455(.A(new_n588), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n657), .A2(new_n619), .A3(new_n635), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n557), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n639), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n659), .A2(new_n660), .A3(new_n503), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n661), .B(KEYINPUT45), .Z(new_n662));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n663), .B1(new_n502), .B2(new_n635), .ZN(new_n664));
  INV_X1    g463(.A(new_n459), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n665), .B1(new_n470), .B2(new_n471), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT89), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n264), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n668), .B1(new_n448), .B2(new_n667), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n666), .A2(new_n375), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n463), .A2(new_n464), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n454), .B1(new_n671), .B2(new_n469), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n491), .B(new_n444), .C1(new_n670), .C2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n453), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n500), .B1(new_n497), .B2(new_n498), .ZN(new_n675));
  AOI211_X1 g474(.A(KEYINPUT74), .B(KEYINPUT36), .C1(new_n496), .C2(new_n417), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n673), .B(new_n674), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n380), .A2(new_n443), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n451), .A2(KEYINPUT35), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n681), .A2(KEYINPUT44), .A3(new_n636), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n664), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT106), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n588), .B(new_n684), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n685), .A2(new_n556), .A3(new_n619), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n503), .B1(new_n687), .B2(new_n660), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n662), .A2(new_n688), .ZN(G1328gat));
  AND2_X1   g488(.A1(new_n683), .A2(new_n686), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n690), .A2(KEYINPUT108), .A3(new_n646), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT108), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n692), .B1(new_n687), .B2(new_n643), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n691), .A2(G36gat), .A3(new_n693), .ZN(new_n694));
  OR3_X1    g493(.A1(new_n659), .A2(G36gat), .A3(new_n643), .ZN(new_n695));
  AND2_X1   g494(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n696));
  NOR2_X1   g495(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n695), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n694), .B(new_n698), .C1(new_n696), .C2(new_n695), .ZN(G1329gat));
  INV_X1    g498(.A(KEYINPUT109), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT47), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n659), .A2(new_n419), .ZN(new_n702));
  INV_X1    g501(.A(new_n501), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(G43gat), .ZN(new_n704));
  OAI221_X1 g503(.A(new_n701), .B1(new_n702), .B2(G43gat), .C1(new_n687), .C2(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n700), .A2(KEYINPUT47), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n705), .B(new_n706), .Z(G1330gat));
  OAI21_X1  g506(.A(G50gat), .B1(new_n687), .B2(new_n444), .ZN(new_n708));
  OR3_X1    g507(.A1(new_n659), .A2(G50gat), .A3(new_n444), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n710), .B(KEYINPUT48), .Z(G1331gat));
  INV_X1    g510(.A(new_n556), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n712), .A2(new_n588), .A3(new_n636), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n619), .ZN(new_n714));
  XOR2_X1   g513(.A(new_n714), .B(KEYINPUT110), .Z(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(new_n502), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n639), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g517(.A1(new_n715), .A2(new_n643), .A3(new_n502), .ZN(new_n719));
  NOR2_X1   g518(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n720));
  AND2_X1   g519(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(new_n719), .B2(new_n720), .ZN(G1333gat));
  NAND2_X1  g522(.A1(new_n716), .A2(new_n703), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n419), .A2(G71gat), .ZN(new_n725));
  AOI22_X1  g524(.A1(new_n724), .A2(G71gat), .B1(new_n716), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g526(.A1(new_n716), .A2(new_n442), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G78gat), .ZN(G1335gat));
  INV_X1    g528(.A(new_n619), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n502), .A2(new_n635), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n657), .A2(new_n712), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT51), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n731), .A2(KEYINPUT51), .A3(new_n732), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n730), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n737), .A2(new_n597), .A3(new_n639), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n657), .A2(new_n712), .A3(new_n730), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n664), .A2(new_n682), .A3(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n664), .A2(new_n682), .A3(KEYINPUT111), .A4(new_n739), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n742), .A2(new_n639), .A3(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n738), .B1(new_n597), .B2(new_n744), .ZN(G1336gat));
  NOR2_X1   g544(.A1(new_n643), .A2(G92gat), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n737), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n747), .A2(KEYINPUT52), .ZN(new_n748));
  OAI21_X1  g547(.A(G92gat), .B1(new_n740), .B2(new_n643), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n742), .A2(new_n646), .A3(new_n743), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT112), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n751), .A2(new_n752), .A3(G92gat), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n752), .B1(new_n751), .B2(G92gat), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n753), .A2(new_n754), .A3(new_n747), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT52), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n750), .B1(new_n755), .B2(new_n756), .ZN(G1337gat));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n703), .A3(new_n743), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(G99gat), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n735), .A2(new_n736), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n419), .A2(G99gat), .A3(new_n730), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT113), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n759), .A2(new_n763), .ZN(G1338gat));
  NOR2_X1   g563(.A1(new_n444), .A2(G106gat), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT53), .B1(new_n737), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT115), .ZN(new_n767));
  XOR2_X1   g566(.A(KEYINPUT114), .B(G106gat), .Z(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n740), .B2(new_n444), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n767), .B1(new_n766), .B2(new_n769), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n742), .A2(new_n442), .A3(new_n743), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n773), .A2(new_n768), .B1(new_n737), .B2(new_n765), .ZN(new_n774));
  OAI22_X1  g573(.A1(new_n770), .A2(new_n771), .B1(new_n772), .B2(new_n774), .ZN(G1339gat));
  AND2_X1   g574(.A1(new_n713), .A2(new_n730), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n543), .A2(new_n553), .A3(new_n548), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n533), .B1(new_n532), .B2(new_n537), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n549), .A2(new_n550), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n547), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n777), .A2(new_n619), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n609), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n607), .A2(new_n608), .A3(new_n591), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n784), .A2(KEYINPUT54), .A3(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n616), .B1(new_n609), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(KEYINPUT55), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n618), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT55), .B1(new_n786), .B2(new_n788), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(new_n554), .B2(new_n555), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n777), .A2(KEYINPUT116), .A3(new_n619), .A4(new_n780), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n783), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n635), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n777), .A2(new_n780), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n797), .A2(new_n636), .A3(new_n792), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n685), .B1(new_n799), .B2(KEYINPUT117), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT117), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n796), .A2(new_n801), .A3(new_n798), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n776), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n803), .A2(new_n419), .A3(new_n442), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n646), .A2(new_n660), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(G113gat), .B1(new_n806), .B2(new_n556), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n803), .A2(new_n660), .A3(new_n646), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n444), .A2(new_n450), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n712), .A2(new_n214), .A3(new_n215), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT118), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n807), .B1(new_n811), .B2(new_n813), .ZN(G1340gat));
  OAI21_X1  g613(.A(G120gat), .B1(new_n806), .B2(new_n730), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n619), .A2(new_n211), .ZN(new_n816));
  XOR2_X1   g615(.A(new_n816), .B(KEYINPUT119), .Z(new_n817));
  OAI21_X1  g616(.A(new_n815), .B1(new_n811), .B2(new_n817), .ZN(G1341gat));
  INV_X1    g617(.A(new_n685), .ZN(new_n819));
  OAI21_X1  g618(.A(G127gat), .B1(new_n806), .B2(new_n819), .ZN(new_n820));
  OR2_X1    g619(.A1(new_n588), .A2(G127gat), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n820), .B1(new_n811), .B2(new_n821), .ZN(G1342gat));
  OR3_X1    g621(.A1(new_n811), .A2(G134gat), .A3(new_n635), .ZN(new_n823));
  OR2_X1    g622(.A1(new_n823), .A2(KEYINPUT56), .ZN(new_n824));
  OAI21_X1  g623(.A(G134gat), .B1(new_n806), .B2(new_n635), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(KEYINPUT56), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(G1343gat));
  NOR2_X1   g626(.A1(new_n803), .A2(new_n444), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT57), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n501), .A2(new_n805), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n793), .A2(new_n781), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n635), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n657), .B1(new_n833), .B2(new_n798), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n442), .B1(new_n776), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n831), .B1(new_n835), .B2(KEYINPUT57), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n830), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(G141gat), .B1(new_n837), .B2(new_n556), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n703), .A2(new_n444), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n808), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n840), .A2(new_n224), .A3(new_n712), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g642(.A1(new_n840), .A2(new_n225), .A3(new_n619), .ZN(new_n844));
  INV_X1    g643(.A(new_n837), .ZN(new_n845));
  AOI211_X1 g644(.A(KEYINPUT59), .B(new_n225), .C1(new_n845), .C2(new_n619), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT59), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT57), .B1(new_n803), .B2(new_n444), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n636), .A2(new_n792), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(KEYINPUT120), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n797), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n657), .B1(new_n851), .B2(new_n833), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n829), .B(new_n442), .C1(new_n852), .C2(new_n776), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n848), .A2(new_n619), .A3(new_n853), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n854), .A2(new_n831), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n847), .B1(new_n855), .B2(G148gat), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n844), .B1(new_n846), .B2(new_n856), .ZN(G1345gat));
  OAI21_X1  g656(.A(G155gat), .B1(new_n837), .B2(new_n819), .ZN(new_n858));
  INV_X1    g657(.A(G155gat), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n840), .A2(new_n859), .A3(new_n657), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n860), .ZN(G1346gat));
  AOI21_X1  g660(.A(G162gat), .B1(new_n840), .B2(new_n636), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n636), .A2(G162gat), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n845), .B2(new_n863), .ZN(G1347gat));
  INV_X1    g663(.A(G169gat), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n646), .A2(new_n660), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n803), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n810), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n865), .B1(new_n868), .B2(new_n556), .ZN(new_n869));
  XOR2_X1   g668(.A(new_n866), .B(KEYINPUT121), .Z(new_n870));
  NAND4_X1  g669(.A1(new_n804), .A2(G169gat), .A3(new_n712), .A4(new_n870), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n869), .A2(new_n871), .ZN(G1348gat));
  NAND2_X1  g671(.A1(new_n804), .A2(new_n870), .ZN(new_n873));
  OAI21_X1  g672(.A(G176gat), .B1(new_n873), .B2(new_n730), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n730), .A2(G176gat), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n874), .B1(new_n868), .B2(new_n875), .ZN(G1349gat));
  OAI21_X1  g675(.A(G183gat), .B1(new_n873), .B2(new_n819), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n657), .A2(new_n309), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n877), .B1(new_n868), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(KEYINPUT123), .B1(KEYINPUT122), .B2(KEYINPUT60), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(KEYINPUT123), .A2(KEYINPUT60), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n877), .B(new_n880), .C1(new_n868), .C2(new_n878), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(G1350gat));
  NOR3_X1   g684(.A1(new_n868), .A2(G190gat), .A3(new_n635), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT124), .ZN(new_n887));
  OAI21_X1  g686(.A(G190gat), .B1(new_n873), .B2(new_n635), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT61), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n889), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n887), .A2(new_n890), .A3(new_n891), .ZN(G1351gat));
  NAND2_X1  g691(.A1(new_n867), .A2(new_n839), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n893), .A2(G197gat), .A3(new_n556), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT125), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n870), .A2(new_n501), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n848), .A2(new_n853), .A3(new_n896), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n897), .A2(new_n712), .ZN(new_n898));
  INV_X1    g697(.A(G197gat), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n895), .B1(new_n898), .B2(new_n899), .ZN(G1352gat));
  NOR2_X1   g699(.A1(new_n730), .A2(G204gat), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n867), .A2(new_n839), .A3(new_n901), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n902), .A2(KEYINPUT126), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(KEYINPUT126), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n903), .A2(KEYINPUT62), .A3(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n896), .ZN(new_n906));
  OAI21_X1  g705(.A(G204gat), .B1(new_n854), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(KEYINPUT62), .B1(new_n903), .B2(new_n904), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n908), .A2(new_n909), .ZN(G1353gat));
  NAND4_X1  g709(.A1(new_n867), .A2(new_n329), .A3(new_n657), .A4(new_n839), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n848), .A2(new_n657), .A3(new_n853), .A4(new_n896), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n912), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT63), .B1(new_n912), .B2(G211gat), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(KEYINPUT127), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n917), .B(new_n911), .C1(new_n913), .C2(new_n914), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1354gat));
  AND2_X1   g718(.A1(new_n897), .A2(new_n636), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n636), .A2(new_n330), .ZN(new_n921));
  OAI22_X1  g720(.A1(new_n920), .A2(new_n330), .B1(new_n893), .B2(new_n921), .ZN(G1355gat));
endmodule


