

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U557 ( .A1(n525), .A2(G2105), .ZN(n539) );
  BUF_X2 U558 ( .A(n623), .Z(n523) );
  NOR2_X1 U559 ( .A1(n790), .A2(n777), .ZN(n778) );
  BUF_X1 U560 ( .A(n697), .Z(G160) );
  INV_X1 U561 ( .A(KEYINPUT100), .ZN(n710) );
  XNOR2_X1 U562 ( .A(KEYINPUT30), .B(KEYINPUT102), .ZN(n745) );
  XNOR2_X1 U563 ( .A(n746), .B(n745), .ZN(n747) );
  INV_X1 U564 ( .A(KEYINPUT31), .ZN(n752) );
  NAND2_X1 U565 ( .A1(n755), .A2(n754), .ZN(n769) );
  INV_X1 U566 ( .A(n969), .ZN(n777) );
  AND2_X1 U567 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U568 ( .A(G2104), .B(KEYINPUT64), .ZN(n524) );
  XNOR2_X1 U569 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U570 ( .A(KEYINPUT70), .B(n603), .ZN(n964) );
  NAND2_X1 U571 ( .A1(n594), .A2(n593), .ZN(n971) );
  NOR2_X1 U572 ( .A1(n535), .A2(n534), .ZN(n697) );
  NOR2_X1 U573 ( .A1(n543), .A2(n542), .ZN(G164) );
  AND2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n897) );
  NAND2_X1 U575 ( .A1(n897), .A2(G113), .ZN(n529) );
  INV_X1 U576 ( .A(n524), .ZN(n525) );
  NAND2_X1 U577 ( .A1(n539), .A2(G101), .ZN(n527) );
  INV_X1 U578 ( .A(KEYINPUT23), .ZN(n526) );
  NAND2_X1 U579 ( .A1(n529), .A2(n528), .ZN(n535) );
  XOR2_X1 U580 ( .A(G2104), .B(KEYINPUT64), .Z(n530) );
  AND2_X2 U581 ( .A1(n530), .A2(G2105), .ZN(n898) );
  NAND2_X1 U582 ( .A1(G125), .A2(n898), .ZN(n533) );
  NOR2_X1 U583 ( .A1(G2104), .A2(G2105), .ZN(n531) );
  XOR2_X1 U584 ( .A(KEYINPUT17), .B(n531), .Z(n623) );
  NAND2_X1 U585 ( .A1(G137), .A2(n523), .ZN(n532) );
  NAND2_X1 U586 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U587 ( .A1(G114), .A2(n897), .ZN(n537) );
  NAND2_X1 U588 ( .A1(G126), .A2(n898), .ZN(n536) );
  NAND2_X1 U589 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U590 ( .A(KEYINPUT86), .B(n538), .ZN(n543) );
  BUF_X1 U591 ( .A(n539), .Z(n902) );
  NAND2_X1 U592 ( .A1(n902), .A2(G102), .ZN(n541) );
  NAND2_X1 U593 ( .A1(n523), .A2(G138), .ZN(n540) );
  NAND2_X1 U594 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U595 ( .A(G2443), .B(G2446), .Z(n545) );
  XNOR2_X1 U596 ( .A(G2427), .B(G2451), .ZN(n544) );
  XNOR2_X1 U597 ( .A(n545), .B(n544), .ZN(n551) );
  XOR2_X1 U598 ( .A(G2430), .B(G2454), .Z(n547) );
  XNOR2_X1 U599 ( .A(G1341), .B(G1348), .ZN(n546) );
  XNOR2_X1 U600 ( .A(n547), .B(n546), .ZN(n549) );
  XOR2_X1 U601 ( .A(G2435), .B(G2438), .Z(n548) );
  XNOR2_X1 U602 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U603 ( .A(n551), .B(n550), .Z(n552) );
  AND2_X1 U604 ( .A1(G14), .A2(n552), .ZN(G401) );
  AND2_X1 U605 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U606 ( .A(G57), .ZN(G237) );
  INV_X1 U607 ( .A(G82), .ZN(G220) );
  NOR2_X1 U608 ( .A1(G651), .A2(G543), .ZN(n663) );
  NAND2_X1 U609 ( .A1(G88), .A2(n663), .ZN(n554) );
  XOR2_X1 U610 ( .A(KEYINPUT0), .B(G543), .Z(n642) );
  INV_X1 U611 ( .A(G651), .ZN(n555) );
  NOR2_X2 U612 ( .A1(n642), .A2(n555), .ZN(n664) );
  NAND2_X1 U613 ( .A1(G75), .A2(n664), .ZN(n553) );
  NAND2_X1 U614 ( .A1(n554), .A2(n553), .ZN(n560) );
  NOR2_X1 U615 ( .A1(G543), .A2(n555), .ZN(n556) );
  XOR2_X2 U616 ( .A(KEYINPUT1), .B(n556), .Z(n659) );
  NAND2_X1 U617 ( .A1(G62), .A2(n659), .ZN(n558) );
  NOR2_X2 U618 ( .A1(G651), .A2(n642), .ZN(n660) );
  NAND2_X1 U619 ( .A1(G50), .A2(n660), .ZN(n557) );
  NAND2_X1 U620 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U621 ( .A1(n560), .A2(n559), .ZN(G166) );
  NAND2_X1 U622 ( .A1(G64), .A2(n659), .ZN(n562) );
  NAND2_X1 U623 ( .A1(G52), .A2(n660), .ZN(n561) );
  NAND2_X1 U624 ( .A1(n562), .A2(n561), .ZN(n567) );
  NAND2_X1 U625 ( .A1(G90), .A2(n663), .ZN(n564) );
  NAND2_X1 U626 ( .A1(G77), .A2(n664), .ZN(n563) );
  NAND2_X1 U627 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U628 ( .A(KEYINPUT9), .B(n565), .Z(n566) );
  NOR2_X1 U629 ( .A1(n567), .A2(n566), .ZN(G171) );
  NAND2_X1 U630 ( .A1(G63), .A2(n659), .ZN(n569) );
  NAND2_X1 U631 ( .A1(G51), .A2(n660), .ZN(n568) );
  NAND2_X1 U632 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U633 ( .A(KEYINPUT6), .B(n570), .ZN(n578) );
  NAND2_X1 U634 ( .A1(n664), .A2(G76), .ZN(n571) );
  XNOR2_X1 U635 ( .A(KEYINPUT72), .B(n571), .ZN(n575) );
  XOR2_X1 U636 ( .A(KEYINPUT4), .B(KEYINPUT71), .Z(n573) );
  NAND2_X1 U637 ( .A1(G89), .A2(n663), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  NAND2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U640 ( .A(n576), .B(KEYINPUT5), .Z(n577) );
  NOR2_X1 U641 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U642 ( .A(KEYINPUT73), .B(n579), .Z(n580) );
  XOR2_X1 U643 ( .A(KEYINPUT7), .B(n580), .Z(G168) );
  XOR2_X1 U644 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U645 ( .A(KEYINPUT10), .B(KEYINPUT67), .Z(n582) );
  NAND2_X1 U646 ( .A1(G7), .A2(G661), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G223) );
  INV_X1 U648 ( .A(G223), .ZN(n853) );
  NAND2_X1 U649 ( .A1(n853), .A2(G567), .ZN(n583) );
  XOR2_X1 U650 ( .A(KEYINPUT11), .B(n583), .Z(G234) );
  NAND2_X1 U651 ( .A1(n664), .A2(G68), .ZN(n584) );
  XNOR2_X1 U652 ( .A(KEYINPUT68), .B(n584), .ZN(n587) );
  NAND2_X1 U653 ( .A1(n663), .A2(G81), .ZN(n585) );
  XNOR2_X1 U654 ( .A(KEYINPUT12), .B(n585), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U656 ( .A(n588), .B(KEYINPUT13), .ZN(n591) );
  NAND2_X1 U657 ( .A1(n659), .A2(G56), .ZN(n589) );
  XNOR2_X1 U658 ( .A(KEYINPUT14), .B(n589), .ZN(n590) );
  NAND2_X1 U659 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U660 ( .A(n592), .B(KEYINPUT69), .ZN(n594) );
  NAND2_X1 U661 ( .A1(G43), .A2(n660), .ZN(n593) );
  INV_X1 U662 ( .A(n971), .ZN(n595) );
  NAND2_X1 U663 ( .A1(n595), .A2(G860), .ZN(G153) );
  INV_X1 U664 ( .A(G171), .ZN(G301) );
  NAND2_X1 U665 ( .A1(G66), .A2(n659), .ZN(n597) );
  NAND2_X1 U666 ( .A1(G92), .A2(n663), .ZN(n596) );
  NAND2_X1 U667 ( .A1(n597), .A2(n596), .ZN(n601) );
  NAND2_X1 U668 ( .A1(G79), .A2(n664), .ZN(n599) );
  NAND2_X1 U669 ( .A1(G54), .A2(n660), .ZN(n598) );
  NAND2_X1 U670 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U671 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U672 ( .A(KEYINPUT15), .B(n602), .Z(n603) );
  INV_X1 U673 ( .A(G868), .ZN(n679) );
  AND2_X1 U674 ( .A1(n964), .A2(n679), .ZN(n605) );
  NOR2_X1 U675 ( .A1(n679), .A2(G301), .ZN(n604) );
  NOR2_X1 U676 ( .A1(n605), .A2(n604), .ZN(G284) );
  NAND2_X1 U677 ( .A1(G65), .A2(n659), .ZN(n607) );
  NAND2_X1 U678 ( .A1(G53), .A2(n660), .ZN(n606) );
  NAND2_X1 U679 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U680 ( .A1(G91), .A2(n663), .ZN(n609) );
  NAND2_X1 U681 ( .A1(G78), .A2(n664), .ZN(n608) );
  NAND2_X1 U682 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U683 ( .A1(n611), .A2(n610), .ZN(n961) );
  INV_X1 U684 ( .A(n961), .ZN(G299) );
  NOR2_X1 U685 ( .A1(G868), .A2(G299), .ZN(n612) );
  XNOR2_X1 U686 ( .A(n612), .B(KEYINPUT74), .ZN(n614) );
  NOR2_X1 U687 ( .A1(n679), .A2(G286), .ZN(n613) );
  NOR2_X1 U688 ( .A1(n614), .A2(n613), .ZN(G297) );
  INV_X1 U689 ( .A(G559), .ZN(n615) );
  NOR2_X1 U690 ( .A1(G860), .A2(n615), .ZN(n616) );
  XNOR2_X1 U691 ( .A(KEYINPUT75), .B(n616), .ZN(n617) );
  NAND2_X1 U692 ( .A1(n617), .A2(n964), .ZN(n618) );
  XNOR2_X1 U693 ( .A(n618), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U694 ( .A1(G868), .A2(n971), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n964), .A2(G868), .ZN(n619) );
  NOR2_X1 U696 ( .A1(G559), .A2(n619), .ZN(n620) );
  NOR2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U698 ( .A(KEYINPUT76), .B(n622), .ZN(G282) );
  NAND2_X1 U699 ( .A1(G111), .A2(n897), .ZN(n625) );
  NAND2_X1 U700 ( .A1(G135), .A2(n523), .ZN(n624) );
  NAND2_X1 U701 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U702 ( .A1(n898), .A2(G123), .ZN(n626) );
  XOR2_X1 U703 ( .A(KEYINPUT18), .B(n626), .Z(n627) );
  NOR2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n630) );
  NAND2_X1 U705 ( .A1(n902), .A2(G99), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n630), .A2(n629), .ZN(n995) );
  XNOR2_X1 U707 ( .A(G2096), .B(n995), .ZN(n631) );
  NOR2_X1 U708 ( .A1(n631), .A2(G2100), .ZN(n632) );
  XNOR2_X1 U709 ( .A(n632), .B(KEYINPUT77), .ZN(G156) );
  NAND2_X1 U710 ( .A1(G559), .A2(n964), .ZN(n676) );
  XNOR2_X1 U711 ( .A(n971), .B(n676), .ZN(n633) );
  NOR2_X1 U712 ( .A1(n633), .A2(G860), .ZN(n641) );
  NAND2_X1 U713 ( .A1(G67), .A2(n659), .ZN(n635) );
  NAND2_X1 U714 ( .A1(G55), .A2(n660), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n663), .A2(G93), .ZN(n636) );
  XOR2_X1 U717 ( .A(KEYINPUT78), .B(n636), .Z(n637) );
  NOR2_X1 U718 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n664), .A2(G80), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n640), .A2(n639), .ZN(n678) );
  XOR2_X1 U721 ( .A(n641), .B(n678), .Z(G145) );
  NAND2_X1 U722 ( .A1(n642), .A2(G87), .ZN(n647) );
  NAND2_X1 U723 ( .A1(G49), .A2(n660), .ZN(n644) );
  NAND2_X1 U724 ( .A1(G74), .A2(G651), .ZN(n643) );
  NAND2_X1 U725 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U726 ( .A1(n659), .A2(n645), .ZN(n646) );
  NAND2_X1 U727 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U728 ( .A(KEYINPUT79), .B(n648), .Z(G288) );
  NAND2_X1 U729 ( .A1(G61), .A2(n659), .ZN(n649) );
  XNOR2_X1 U730 ( .A(n649), .B(KEYINPUT80), .ZN(n658) );
  NAND2_X1 U731 ( .A1(G73), .A2(n664), .ZN(n650) );
  XNOR2_X1 U732 ( .A(n650), .B(KEYINPUT82), .ZN(n651) );
  XNOR2_X1 U733 ( .A(n651), .B(KEYINPUT2), .ZN(n653) );
  NAND2_X1 U734 ( .A1(G48), .A2(n660), .ZN(n652) );
  NAND2_X1 U735 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U736 ( .A1(G86), .A2(n663), .ZN(n654) );
  XNOR2_X1 U737 ( .A(KEYINPUT81), .B(n654), .ZN(n655) );
  NOR2_X1 U738 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U739 ( .A1(n658), .A2(n657), .ZN(G305) );
  NAND2_X1 U740 ( .A1(G60), .A2(n659), .ZN(n662) );
  NAND2_X1 U741 ( .A1(G47), .A2(n660), .ZN(n661) );
  NAND2_X1 U742 ( .A1(n662), .A2(n661), .ZN(n668) );
  NAND2_X1 U743 ( .A1(G85), .A2(n663), .ZN(n666) );
  NAND2_X1 U744 ( .A1(G72), .A2(n664), .ZN(n665) );
  NAND2_X1 U745 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U746 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U747 ( .A(n669), .B(KEYINPUT65), .ZN(G290) );
  XOR2_X1 U748 ( .A(n971), .B(G305), .Z(n670) );
  XNOR2_X1 U749 ( .A(G288), .B(n670), .ZN(n671) );
  XNOR2_X1 U750 ( .A(KEYINPUT19), .B(n671), .ZN(n673) );
  XNOR2_X1 U751 ( .A(G290), .B(G166), .ZN(n672) );
  XNOR2_X1 U752 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U753 ( .A(n961), .B(n674), .ZN(n675) );
  XNOR2_X1 U754 ( .A(n675), .B(n678), .ZN(n919) );
  XOR2_X1 U755 ( .A(n919), .B(n676), .Z(n677) );
  NOR2_X1 U756 ( .A1(n679), .A2(n677), .ZN(n681) );
  AND2_X1 U757 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U758 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U759 ( .A(KEYINPUT83), .B(n682), .ZN(G295) );
  NAND2_X1 U760 ( .A1(G2078), .A2(G2084), .ZN(n683) );
  XOR2_X1 U761 ( .A(KEYINPUT20), .B(n683), .Z(n684) );
  NAND2_X1 U762 ( .A1(G2090), .A2(n684), .ZN(n686) );
  XNOR2_X1 U763 ( .A(KEYINPUT84), .B(KEYINPUT21), .ZN(n685) );
  XNOR2_X1 U764 ( .A(n686), .B(n685), .ZN(n687) );
  NAND2_X1 U765 ( .A1(G2072), .A2(n687), .ZN(G158) );
  XNOR2_X1 U766 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U767 ( .A(KEYINPUT66), .B(G132), .Z(G219) );
  NOR2_X1 U768 ( .A1(G219), .A2(G220), .ZN(n688) );
  XOR2_X1 U769 ( .A(KEYINPUT22), .B(n688), .Z(n689) );
  NOR2_X1 U770 ( .A1(G218), .A2(n689), .ZN(n690) );
  NAND2_X1 U771 ( .A1(G96), .A2(n690), .ZN(n857) );
  NAND2_X1 U772 ( .A1(n857), .A2(G2106), .ZN(n694) );
  NAND2_X1 U773 ( .A1(G69), .A2(G120), .ZN(n691) );
  NOR2_X1 U774 ( .A1(G237), .A2(n691), .ZN(n692) );
  NAND2_X1 U775 ( .A1(G108), .A2(n692), .ZN(n858) );
  NAND2_X1 U776 ( .A1(n858), .A2(G567), .ZN(n693) );
  NAND2_X1 U777 ( .A1(n694), .A2(n693), .ZN(n930) );
  NAND2_X1 U778 ( .A1(G661), .A2(G483), .ZN(n695) );
  NOR2_X1 U779 ( .A1(n930), .A2(n695), .ZN(n856) );
  NAND2_X1 U780 ( .A1(G36), .A2(n856), .ZN(n696) );
  XOR2_X1 U781 ( .A(KEYINPUT85), .B(n696), .Z(G176) );
  INV_X1 U782 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U783 ( .A(KEYINPUT40), .B(KEYINPUT108), .ZN(n852) );
  NOR2_X1 U784 ( .A1(G164), .A2(G1384), .ZN(n816) );
  INV_X1 U785 ( .A(KEYINPUT94), .ZN(n698) );
  NAND2_X1 U786 ( .A1(n697), .A2(G40), .ZN(n815) );
  XNOR2_X1 U787 ( .A(n698), .B(n815), .ZN(n699) );
  NAND2_X1 U788 ( .A1(n816), .A2(n699), .ZN(n757) );
  NAND2_X1 U789 ( .A1(G8), .A2(n757), .ZN(n790) );
  NOR2_X1 U790 ( .A1(G1976), .A2(G288), .ZN(n775) );
  NAND2_X1 U791 ( .A1(n775), .A2(KEYINPUT33), .ZN(n700) );
  NOR2_X1 U792 ( .A1(n790), .A2(n700), .ZN(n782) );
  INV_X1 U793 ( .A(G1996), .ZN(n1017) );
  NOR2_X1 U794 ( .A1(n757), .A2(n1017), .ZN(n702) );
  INV_X1 U795 ( .A(KEYINPUT26), .ZN(n701) );
  XNOR2_X1 U796 ( .A(n702), .B(n701), .ZN(n704) );
  NAND2_X1 U797 ( .A1(n757), .A2(G1341), .ZN(n703) );
  NAND2_X1 U798 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U799 ( .A1(n971), .A2(n705), .ZN(n712) );
  NAND2_X1 U800 ( .A1(n712), .A2(n964), .ZN(n709) );
  INV_X1 U801 ( .A(n757), .ZN(n732) );
  NOR2_X1 U802 ( .A1(n732), .A2(G1348), .ZN(n707) );
  NOR2_X1 U803 ( .A1(G2067), .A2(n757), .ZN(n706) );
  NOR2_X1 U804 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U805 ( .A1(n709), .A2(n708), .ZN(n711) );
  XNOR2_X1 U806 ( .A(n711), .B(n710), .ZN(n714) );
  NOR2_X1 U807 ( .A1(n712), .A2(n964), .ZN(n713) );
  NOR2_X1 U808 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U809 ( .A(n715), .B(KEYINPUT101), .ZN(n721) );
  NAND2_X1 U810 ( .A1(G1956), .A2(n757), .ZN(n716) );
  XNOR2_X1 U811 ( .A(KEYINPUT99), .B(n716), .ZN(n719) );
  NAND2_X1 U812 ( .A1(n732), .A2(G2072), .ZN(n717) );
  XNOR2_X1 U813 ( .A(KEYINPUT27), .B(n717), .ZN(n718) );
  NOR2_X1 U814 ( .A1(n719), .A2(n718), .ZN(n722) );
  NAND2_X1 U815 ( .A1(n722), .A2(n961), .ZN(n720) );
  NAND2_X1 U816 ( .A1(n721), .A2(n720), .ZN(n725) );
  NOR2_X1 U817 ( .A1(n722), .A2(n961), .ZN(n723) );
  XOR2_X1 U818 ( .A(n723), .B(KEYINPUT28), .Z(n724) );
  NAND2_X1 U819 ( .A1(n725), .A2(n724), .ZN(n727) );
  INV_X1 U820 ( .A(KEYINPUT29), .ZN(n726) );
  XNOR2_X1 U821 ( .A(n727), .B(n726), .ZN(n741) );
  XNOR2_X1 U822 ( .A(G1961), .B(KEYINPUT96), .ZN(n945) );
  NOR2_X1 U823 ( .A1(n732), .A2(n945), .ZN(n728) );
  NAND2_X1 U824 ( .A1(KEYINPUT98), .A2(n728), .ZN(n729) );
  NAND2_X1 U825 ( .A1(n729), .A2(KEYINPUT97), .ZN(n739) );
  XNOR2_X1 U826 ( .A(KEYINPUT25), .B(G2078), .ZN(n1020) );
  NAND2_X1 U827 ( .A1(KEYINPUT98), .A2(n1020), .ZN(n730) );
  NOR2_X1 U828 ( .A1(n757), .A2(n730), .ZN(n734) );
  AND2_X1 U829 ( .A1(KEYINPUT98), .A2(n945), .ZN(n731) );
  NOR2_X1 U830 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U831 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U832 ( .A1(KEYINPUT97), .A2(n735), .ZN(n737) );
  NOR2_X1 U833 ( .A1(KEYINPUT98), .A2(n1020), .ZN(n736) );
  NOR2_X1 U834 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U835 ( .A1(n739), .A2(n738), .ZN(n748) );
  NAND2_X1 U836 ( .A1(n748), .A2(G171), .ZN(n740) );
  NAND2_X1 U837 ( .A1(n741), .A2(n740), .ZN(n755) );
  NOR2_X1 U838 ( .A1(G1966), .A2(n790), .ZN(n742) );
  XOR2_X1 U839 ( .A(KEYINPUT95), .B(n742), .Z(n771) );
  NOR2_X1 U840 ( .A1(G2084), .A2(n757), .ZN(n767) );
  INV_X1 U841 ( .A(n767), .ZN(n743) );
  NAND2_X1 U842 ( .A1(G8), .A2(n743), .ZN(n744) );
  OR2_X1 U843 ( .A1(n771), .A2(n744), .ZN(n746) );
  NOR2_X1 U844 ( .A1(n747), .A2(G168), .ZN(n751) );
  NOR2_X1 U845 ( .A1(G171), .A2(n748), .ZN(n749) );
  XOR2_X1 U846 ( .A(KEYINPUT103), .B(n749), .Z(n750) );
  NOR2_X1 U847 ( .A1(n751), .A2(n750), .ZN(n753) );
  XNOR2_X1 U848 ( .A(n753), .B(n752), .ZN(n754) );
  AND2_X1 U849 ( .A1(G286), .A2(G8), .ZN(n756) );
  NAND2_X1 U850 ( .A1(n769), .A2(n756), .ZN(n764) );
  INV_X1 U851 ( .A(G8), .ZN(n762) );
  NOR2_X1 U852 ( .A1(G1971), .A2(n790), .ZN(n759) );
  NOR2_X1 U853 ( .A1(G2090), .A2(n757), .ZN(n758) );
  NOR2_X1 U854 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U855 ( .A1(n760), .A2(G303), .ZN(n761) );
  OR2_X1 U856 ( .A1(n762), .A2(n761), .ZN(n763) );
  AND2_X1 U857 ( .A1(n764), .A2(n763), .ZN(n766) );
  XOR2_X1 U858 ( .A(KEYINPUT32), .B(KEYINPUT104), .Z(n765) );
  XNOR2_X1 U859 ( .A(n766), .B(n765), .ZN(n773) );
  NAND2_X1 U860 ( .A1(G8), .A2(n767), .ZN(n768) );
  NAND2_X1 U861 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X1 U862 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X2 U863 ( .A1(n773), .A2(n772), .ZN(n788) );
  INV_X1 U864 ( .A(n788), .ZN(n776) );
  NOR2_X1 U865 ( .A1(G1971), .A2(G303), .ZN(n774) );
  NOR2_X1 U866 ( .A1(n775), .A2(n774), .ZN(n965) );
  NAND2_X1 U867 ( .A1(n776), .A2(n965), .ZN(n779) );
  NAND2_X1 U868 ( .A1(G1976), .A2(G288), .ZN(n969) );
  NOR2_X1 U869 ( .A1(KEYINPUT33), .A2(n780), .ZN(n781) );
  NOR2_X1 U870 ( .A1(n782), .A2(n781), .ZN(n783) );
  XOR2_X1 U871 ( .A(G1981), .B(G305), .Z(n976) );
  NAND2_X1 U872 ( .A1(n783), .A2(n976), .ZN(n795) );
  NOR2_X1 U873 ( .A1(G1981), .A2(G305), .ZN(n784) );
  XOR2_X1 U874 ( .A(n784), .B(KEYINPUT24), .Z(n785) );
  OR2_X1 U875 ( .A1(n790), .A2(n785), .ZN(n793) );
  NAND2_X1 U876 ( .A1(G166), .A2(G8), .ZN(n786) );
  NOR2_X1 U877 ( .A1(G2090), .A2(n786), .ZN(n787) );
  NOR2_X1 U878 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U879 ( .A(n789), .B(KEYINPUT105), .ZN(n791) );
  NAND2_X1 U880 ( .A1(n791), .A2(n790), .ZN(n792) );
  AND2_X1 U881 ( .A1(n793), .A2(n792), .ZN(n794) );
  AND2_X1 U882 ( .A1(n795), .A2(n794), .ZN(n797) );
  INV_X1 U883 ( .A(KEYINPUT106), .ZN(n796) );
  XNOR2_X1 U884 ( .A(n797), .B(n796), .ZN(n836) );
  NAND2_X1 U885 ( .A1(n898), .A2(G129), .ZN(n804) );
  NAND2_X1 U886 ( .A1(G117), .A2(n897), .ZN(n799) );
  NAND2_X1 U887 ( .A1(G141), .A2(n523), .ZN(n798) );
  NAND2_X1 U888 ( .A1(n799), .A2(n798), .ZN(n802) );
  NAND2_X1 U889 ( .A1(n902), .A2(G105), .ZN(n800) );
  XOR2_X1 U890 ( .A(KEYINPUT38), .B(n800), .Z(n801) );
  NOR2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U892 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U893 ( .A(KEYINPUT91), .B(n805), .Z(n908) );
  NAND2_X1 U894 ( .A1(G1996), .A2(n908), .ZN(n806) );
  XOR2_X1 U895 ( .A(KEYINPUT92), .B(n806), .Z(n814) );
  NAND2_X1 U896 ( .A1(G131), .A2(n523), .ZN(n808) );
  NAND2_X1 U897 ( .A1(G95), .A2(n902), .ZN(n807) );
  NAND2_X1 U898 ( .A1(n808), .A2(n807), .ZN(n812) );
  NAND2_X1 U899 ( .A1(G107), .A2(n897), .ZN(n810) );
  NAND2_X1 U900 ( .A1(G119), .A2(n898), .ZN(n809) );
  NAND2_X1 U901 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U902 ( .A1(n812), .A2(n811), .ZN(n911) );
  INV_X1 U903 ( .A(G1991), .ZN(n1014) );
  NOR2_X1 U904 ( .A1(n911), .A2(n1014), .ZN(n813) );
  NOR2_X1 U905 ( .A1(n814), .A2(n813), .ZN(n1003) );
  NOR2_X1 U906 ( .A1(n816), .A2(n815), .ZN(n847) );
  INV_X1 U907 ( .A(n847), .ZN(n817) );
  NOR2_X1 U908 ( .A1(n1003), .A2(n817), .ZN(n839) );
  INV_X1 U909 ( .A(n839), .ZN(n831) );
  NAND2_X1 U910 ( .A1(G140), .A2(n523), .ZN(n819) );
  NAND2_X1 U911 ( .A1(G104), .A2(n902), .ZN(n818) );
  NAND2_X1 U912 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U913 ( .A(KEYINPUT34), .B(n820), .ZN(n826) );
  NAND2_X1 U914 ( .A1(n897), .A2(G116), .ZN(n821) );
  XNOR2_X1 U915 ( .A(n821), .B(KEYINPUT88), .ZN(n823) );
  NAND2_X1 U916 ( .A1(G128), .A2(n898), .ZN(n822) );
  NAND2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n824) );
  XOR2_X1 U918 ( .A(n824), .B(KEYINPUT35), .Z(n825) );
  NOR2_X1 U919 ( .A1(n826), .A2(n825), .ZN(n827) );
  XOR2_X1 U920 ( .A(KEYINPUT36), .B(n827), .Z(n828) );
  XNOR2_X1 U921 ( .A(KEYINPUT89), .B(n828), .ZN(n916) );
  XOR2_X1 U922 ( .A(G2067), .B(KEYINPUT37), .Z(n829) );
  XNOR2_X1 U923 ( .A(KEYINPUT87), .B(n829), .ZN(n845) );
  NOR2_X1 U924 ( .A1(n916), .A2(n845), .ZN(n998) );
  NAND2_X1 U925 ( .A1(n847), .A2(n998), .ZN(n830) );
  XNOR2_X1 U926 ( .A(KEYINPUT90), .B(n830), .ZN(n843) );
  NAND2_X1 U927 ( .A1(n831), .A2(n843), .ZN(n832) );
  XNOR2_X1 U928 ( .A(KEYINPUT93), .B(n832), .ZN(n834) );
  XNOR2_X1 U929 ( .A(G1986), .B(G290), .ZN(n960) );
  NAND2_X1 U930 ( .A1(n960), .A2(n847), .ZN(n833) );
  AND2_X1 U931 ( .A1(n834), .A2(n833), .ZN(n835) );
  NAND2_X1 U932 ( .A1(n836), .A2(n835), .ZN(n850) );
  NOR2_X1 U933 ( .A1(G1996), .A2(n908), .ZN(n989) );
  AND2_X1 U934 ( .A1(n1014), .A2(n911), .ZN(n994) );
  NOR2_X1 U935 ( .A1(G1986), .A2(G290), .ZN(n837) );
  XOR2_X1 U936 ( .A(n837), .B(KEYINPUT107), .Z(n838) );
  NOR2_X1 U937 ( .A1(n994), .A2(n838), .ZN(n840) );
  NOR2_X1 U938 ( .A1(n840), .A2(n839), .ZN(n841) );
  NOR2_X1 U939 ( .A1(n989), .A2(n841), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n842), .B(KEYINPUT39), .ZN(n844) );
  NAND2_X1 U941 ( .A1(n844), .A2(n843), .ZN(n846) );
  NAND2_X1 U942 ( .A1(n916), .A2(n845), .ZN(n991) );
  NAND2_X1 U943 ( .A1(n846), .A2(n991), .ZN(n848) );
  NAND2_X1 U944 ( .A1(n848), .A2(n847), .ZN(n849) );
  NAND2_X1 U945 ( .A1(n850), .A2(n849), .ZN(n851) );
  XNOR2_X1 U946 ( .A(n852), .B(n851), .ZN(G329) );
  NAND2_X1 U947 ( .A1(G2106), .A2(n853), .ZN(G217) );
  AND2_X1 U948 ( .A1(G15), .A2(G2), .ZN(n854) );
  NAND2_X1 U949 ( .A1(G661), .A2(n854), .ZN(G259) );
  NAND2_X1 U950 ( .A1(G3), .A2(G1), .ZN(n855) );
  NAND2_X1 U951 ( .A1(n856), .A2(n855), .ZN(G188) );
  NOR2_X1 U952 ( .A1(n858), .A2(n857), .ZN(G325) );
  XNOR2_X1 U953 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  INV_X1 U955 ( .A(G120), .ZN(G236) );
  INV_X1 U956 ( .A(G96), .ZN(G221) );
  INV_X1 U957 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U958 ( .A(G1996), .B(G2474), .ZN(n868) );
  XOR2_X1 U959 ( .A(G1956), .B(G1961), .Z(n860) );
  XNOR2_X1 U960 ( .A(G1991), .B(G1986), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U962 ( .A(G1976), .B(G1981), .Z(n862) );
  XNOR2_X1 U963 ( .A(G1971), .B(G1966), .ZN(n861) );
  XNOR2_X1 U964 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U965 ( .A(n864), .B(n863), .Z(n866) );
  XNOR2_X1 U966 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n865) );
  XNOR2_X1 U967 ( .A(n866), .B(n865), .ZN(n867) );
  XNOR2_X1 U968 ( .A(n868), .B(n867), .ZN(G229) );
  XOR2_X1 U969 ( .A(G2100), .B(G2096), .Z(n870) );
  XNOR2_X1 U970 ( .A(KEYINPUT42), .B(G2678), .ZN(n869) );
  XNOR2_X1 U971 ( .A(n870), .B(n869), .ZN(n874) );
  XOR2_X1 U972 ( .A(KEYINPUT43), .B(G2072), .Z(n872) );
  XNOR2_X1 U973 ( .A(G2067), .B(G2090), .ZN(n871) );
  XNOR2_X1 U974 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U975 ( .A(n874), .B(n873), .Z(n876) );
  XNOR2_X1 U976 ( .A(G2078), .B(G2084), .ZN(n875) );
  XNOR2_X1 U977 ( .A(n876), .B(n875), .ZN(G227) );
  NAND2_X1 U978 ( .A1(G112), .A2(n897), .ZN(n878) );
  NAND2_X1 U979 ( .A1(G136), .A2(n523), .ZN(n877) );
  NAND2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n883) );
  NAND2_X1 U981 ( .A1(n898), .A2(G124), .ZN(n879) );
  XNOR2_X1 U982 ( .A(n879), .B(KEYINPUT44), .ZN(n881) );
  NAND2_X1 U983 ( .A1(G100), .A2(n902), .ZN(n880) );
  NAND2_X1 U984 ( .A1(n881), .A2(n880), .ZN(n882) );
  NOR2_X1 U985 ( .A1(n883), .A2(n882), .ZN(G162) );
  NAND2_X1 U986 ( .A1(G115), .A2(n897), .ZN(n885) );
  NAND2_X1 U987 ( .A1(G127), .A2(n898), .ZN(n884) );
  NAND2_X1 U988 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U989 ( .A(n886), .B(KEYINPUT47), .ZN(n888) );
  NAND2_X1 U990 ( .A1(G139), .A2(n523), .ZN(n887) );
  NAND2_X1 U991 ( .A1(n888), .A2(n887), .ZN(n891) );
  NAND2_X1 U992 ( .A1(G103), .A2(n902), .ZN(n889) );
  XNOR2_X1 U993 ( .A(KEYINPUT113), .B(n889), .ZN(n890) );
  NOR2_X1 U994 ( .A1(n891), .A2(n890), .ZN(n983) );
  XNOR2_X1 U995 ( .A(G164), .B(n983), .ZN(n915) );
  XOR2_X1 U996 ( .A(G160), .B(G162), .Z(n892) );
  XNOR2_X1 U997 ( .A(n995), .B(n892), .ZN(n896) );
  XOR2_X1 U998 ( .A(KEYINPUT112), .B(KEYINPUT114), .Z(n894) );
  XNOR2_X1 U999 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n893) );
  XNOR2_X1 U1000 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U1001 ( .A(n896), .B(n895), .Z(n913) );
  NAND2_X1 U1002 ( .A1(G118), .A2(n897), .ZN(n900) );
  NAND2_X1 U1003 ( .A1(G130), .A2(n898), .ZN(n899) );
  NAND2_X1 U1004 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U1005 ( .A(KEYINPUT111), .B(n901), .Z(n907) );
  NAND2_X1 U1006 ( .A1(G142), .A2(n523), .ZN(n904) );
  NAND2_X1 U1007 ( .A1(G106), .A2(n902), .ZN(n903) );
  NAND2_X1 U1008 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U1009 ( .A(n905), .B(KEYINPUT45), .Z(n906) );
  NOR2_X1 U1010 ( .A1(n907), .A2(n906), .ZN(n909) );
  XNOR2_X1 U1011 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1012 ( .A(n911), .B(n910), .ZN(n912) );
  XNOR2_X1 U1013 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1014 ( .A(n915), .B(n914), .ZN(n917) );
  XOR2_X1 U1015 ( .A(n917), .B(n916), .Z(n918) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n918), .ZN(G395) );
  XNOR2_X1 U1017 ( .A(G171), .B(n964), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(n920), .B(n919), .ZN(n921) );
  XOR2_X1 U1019 ( .A(G286), .B(n921), .Z(n922) );
  NOR2_X1 U1020 ( .A1(G37), .A2(n922), .ZN(G397) );
  XNOR2_X1 U1021 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(G229), .A2(G227), .ZN(n923) );
  XNOR2_X1 U1023 ( .A(n924), .B(n923), .ZN(n927) );
  NOR2_X1 U1024 ( .A1(G401), .A2(n930), .ZN(n925) );
  XNOR2_X1 U1025 ( .A(KEYINPUT115), .B(n925), .ZN(n926) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n929) );
  NOR2_X1 U1027 ( .A1(G395), .A2(G397), .ZN(n928) );
  NAND2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(G225) );
  INV_X1 U1029 ( .A(G225), .ZN(G308) );
  INV_X1 U1030 ( .A(n930), .ZN(G319) );
  INV_X1 U1031 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1032 ( .A(G1966), .B(G21), .ZN(n943) );
  XNOR2_X1 U1033 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n931) );
  XNOR2_X1 U1034 ( .A(n931), .B(KEYINPUT60), .ZN(n941) );
  XNOR2_X1 U1035 ( .A(G1348), .B(KEYINPUT59), .ZN(n932) );
  XNOR2_X1 U1036 ( .A(n932), .B(G4), .ZN(n936) );
  XNOR2_X1 U1037 ( .A(G1956), .B(G20), .ZN(n934) );
  XNOR2_X1 U1038 ( .A(G1981), .B(G6), .ZN(n933) );
  NOR2_X1 U1039 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1040 ( .A1(n936), .A2(n935), .ZN(n939) );
  XNOR2_X1 U1041 ( .A(KEYINPUT122), .B(G1341), .ZN(n937) );
  XNOR2_X1 U1042 ( .A(G19), .B(n937), .ZN(n938) );
  NOR2_X1 U1043 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1044 ( .A(n941), .B(n940), .ZN(n942) );
  NOR2_X1 U1045 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1046 ( .A(KEYINPUT125), .B(n944), .Z(n947) );
  XOR2_X1 U1047 ( .A(n945), .B(G5), .Z(n946) );
  NAND2_X1 U1048 ( .A1(n947), .A2(n946), .ZN(n955) );
  XNOR2_X1 U1049 ( .A(G1971), .B(G22), .ZN(n949) );
  XNOR2_X1 U1050 ( .A(G23), .B(G1976), .ZN(n948) );
  NOR2_X1 U1051 ( .A1(n949), .A2(n948), .ZN(n952) );
  XOR2_X1 U1052 ( .A(G1986), .B(KEYINPUT126), .Z(n950) );
  XNOR2_X1 U1053 ( .A(G24), .B(n950), .ZN(n951) );
  NAND2_X1 U1054 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1055 ( .A(KEYINPUT58), .B(n953), .ZN(n954) );
  NOR2_X1 U1056 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1057 ( .A(KEYINPUT61), .B(n956), .Z(n957) );
  NOR2_X1 U1058 ( .A1(G16), .A2(n957), .ZN(n958) );
  XNOR2_X1 U1059 ( .A(KEYINPUT127), .B(n958), .ZN(n1013) );
  XNOR2_X1 U1060 ( .A(G1961), .B(G301), .ZN(n959) );
  NOR2_X1 U1061 ( .A1(n960), .A2(n959), .ZN(n975) );
  XNOR2_X1 U1062 ( .A(G1956), .B(n961), .ZN(n963) );
  NAND2_X1 U1063 ( .A1(G1971), .A2(G303), .ZN(n962) );
  NAND2_X1 U1064 ( .A1(n963), .A2(n962), .ZN(n968) );
  XNOR2_X1 U1065 ( .A(G1348), .B(n964), .ZN(n966) );
  NAND2_X1 U1066 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1067 ( .A1(n968), .A2(n967), .ZN(n970) );
  NAND2_X1 U1068 ( .A1(n970), .A2(n969), .ZN(n973) );
  XNOR2_X1 U1069 ( .A(G1341), .B(n971), .ZN(n972) );
  NOR2_X1 U1070 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(G168), .B(G1966), .ZN(n977) );
  NAND2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1074 ( .A(KEYINPUT57), .B(n978), .Z(n979) );
  NOR2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n982) );
  XOR2_X1 U1076 ( .A(KEYINPUT56), .B(G16), .Z(n981) );
  NOR2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n1011) );
  XNOR2_X1 U1078 ( .A(G2072), .B(n983), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(G164), .B(G2078), .ZN(n984) );
  XNOR2_X1 U1080 ( .A(n984), .B(KEYINPUT118), .ZN(n985) );
  NAND2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1082 ( .A(n987), .B(KEYINPUT50), .ZN(n1005) );
  XOR2_X1 U1083 ( .A(G2090), .B(G162), .Z(n988) );
  NOR2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n990) );
  XOR2_X1 U1085 ( .A(KEYINPUT51), .B(n990), .Z(n992) );
  NAND2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n1001) );
  XOR2_X1 U1087 ( .A(G160), .B(G2084), .Z(n993) );
  NOR2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n996) );
  NAND2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1091 ( .A(KEYINPUT117), .B(n999), .ZN(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1095 ( .A(KEYINPUT52), .B(n1006), .Z(n1007) );
  NOR2_X1 U1096 ( .A1(KEYINPUT55), .A2(n1007), .ZN(n1009) );
  INV_X1 U1097 ( .A(G29), .ZN(n1008) );
  NOR2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1039) );
  XNOR2_X1 U1101 ( .A(G29), .B(KEYINPUT121), .ZN(n1036) );
  XOR2_X1 U1102 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n1034) );
  XNOR2_X1 U1103 ( .A(G2090), .B(G35), .ZN(n1029) );
  XNOR2_X1 U1104 ( .A(G25), .B(n1014), .ZN(n1015) );
  NAND2_X1 U1105 ( .A1(n1015), .A2(G28), .ZN(n1026) );
  XNOR2_X1 U1106 ( .A(KEYINPUT119), .B(G2072), .ZN(n1016) );
  XNOR2_X1 U1107 ( .A(n1016), .B(G33), .ZN(n1024) );
  XOR2_X1 U1108 ( .A(G2067), .B(G26), .Z(n1019) );
  XNOR2_X1 U1109 ( .A(n1017), .B(G32), .ZN(n1018) );
  NAND2_X1 U1110 ( .A1(n1019), .A2(n1018), .ZN(n1022) );
  XOR2_X1 U1111 ( .A(G27), .B(n1020), .Z(n1021) );
  NOR2_X1 U1112 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1113 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1115 ( .A(KEYINPUT53), .B(n1027), .ZN(n1028) );
  NOR2_X1 U1116 ( .A1(n1029), .A2(n1028), .ZN(n1032) );
  XOR2_X1 U1117 ( .A(G2084), .B(G34), .Z(n1030) );
  XNOR2_X1 U1118 ( .A(KEYINPUT54), .B(n1030), .ZN(n1031) );
  NAND2_X1 U1119 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1120 ( .A(n1034), .B(n1033), .ZN(n1035) );
  NAND2_X1 U1121 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NAND2_X1 U1122 ( .A1(n1037), .A2(G11), .ZN(n1038) );
  NOR2_X1 U1123 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  XNOR2_X1 U1124 ( .A(n1040), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1125 ( .A(G311), .ZN(G150) );
endmodule

