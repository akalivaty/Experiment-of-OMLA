//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 1 0 0 0 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G128), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT24), .B(G110), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n194), .B1(new_n187), .B2(G128), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n189), .A2(KEYINPUT23), .A3(G119), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(new_n188), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n193), .B1(G110), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G140), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G125), .ZN(new_n200));
  INV_X1    g014(.A(G125), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G140), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(new_n202), .A3(KEYINPUT16), .ZN(new_n203));
  OR3_X1    g017(.A1(new_n201), .A2(KEYINPUT16), .A3(G140), .ZN(new_n204));
  AOI21_X1  g018(.A(G146), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT72), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n203), .A2(new_n204), .A3(G146), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n209), .B1(new_n205), .B2(new_n206), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n198), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n191), .A2(new_n192), .ZN(new_n212));
  INV_X1    g026(.A(G110), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n195), .A2(new_n196), .A3(new_n213), .A4(new_n188), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  XNOR2_X1  g029(.A(G125), .B(G140), .ZN(new_n216));
  AOI22_X1  g030(.A1(new_n212), .A2(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n209), .A2(KEYINPUT73), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT73), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n203), .A2(new_n204), .A3(new_n219), .A4(G146), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n217), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT74), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT74), .A4(new_n220), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n211), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G953), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(G221), .A3(G234), .ZN(new_n227));
  XOR2_X1   g041(.A(new_n227), .B(KEYINPUT75), .Z(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT22), .B(G137), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n228), .A2(new_n229), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n225), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G902), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n232), .A2(new_n211), .A3(new_n223), .A4(new_n224), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT25), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT25), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n234), .A2(new_n239), .A3(new_n235), .A4(new_n236), .ZN(new_n240));
  NAND2_X1  g054(.A1(G217), .A2(G902), .ZN(new_n241));
  INV_X1    g055(.A(G217), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n241), .B1(new_n242), .B2(G234), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n243), .B(KEYINPUT71), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n238), .A2(new_n240), .A3(new_n244), .ZN(new_n245));
  AND2_X1   g059(.A1(new_n234), .A2(new_n236), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n244), .A2(G902), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  XOR2_X1   g063(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n250));
  NOR2_X1   g064(.A1(G237), .A2(G953), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G210), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n250), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT26), .B(G101), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n253), .B(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n187), .A2(G116), .ZN(new_n256));
  INV_X1    g070(.A(G116), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G119), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT2), .B(G113), .ZN(new_n260));
  OR2_X1    g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n260), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OR2_X1    g077(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n264));
  NAND2_X1  g078(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n265));
  INV_X1    g079(.A(G137), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n264), .A2(new_n265), .B1(G134), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(G134), .ZN(new_n269));
  INV_X1    g083(.A(G134), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G137), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n268), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(G131), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n269), .B1(new_n274), .B2(new_n268), .ZN(new_n275));
  INV_X1    g089(.A(G131), .ZN(new_n276));
  XNOR2_X1  g090(.A(G134), .B(G137), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n275), .B(new_n276), .C1(new_n268), .C2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n273), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(G143), .B(G146), .ZN(new_n280));
  NAND2_X1  g094(.A1(KEYINPUT0), .A2(G128), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XOR2_X1   g096(.A(KEYINPUT0), .B(G128), .Z(new_n283));
  OAI21_X1  g097(.A(new_n282), .B1(new_n283), .B2(new_n280), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n263), .B1(new_n279), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G143), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(KEYINPUT1), .A3(G146), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n287), .B1(new_n280), .B2(G128), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n189), .A2(KEYINPUT1), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n215), .A2(G143), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n286), .A2(G146), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT66), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n280), .A2(KEYINPUT66), .A3(new_n289), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n288), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  OR2_X1    g110(.A1(new_n277), .A2(new_n276), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n278), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT67), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n290), .A2(new_n291), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n215), .A2(G143), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n300), .A2(new_n189), .B1(KEYINPUT1), .B2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT66), .B1(new_n280), .B2(new_n289), .ZN(new_n303));
  AND4_X1   g117(.A1(KEYINPUT66), .A2(new_n289), .A3(new_n290), .A4(new_n291), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT67), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n305), .A2(new_n306), .A3(new_n278), .A4(new_n297), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n285), .A2(new_n299), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT68), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT68), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n285), .A2(new_n299), .A3(new_n307), .A4(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT65), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n294), .A2(new_n295), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n298), .A2(new_n313), .B1(new_n314), .B2(new_n302), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n278), .A2(KEYINPUT65), .A3(new_n297), .ZN(new_n316));
  AOI22_X1  g130(.A1(new_n315), .A2(new_n316), .B1(new_n279), .B2(new_n284), .ZN(new_n317));
  INV_X1    g131(.A(new_n263), .ZN(new_n318));
  OR2_X1    g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n312), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT28), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n285), .B1(new_n298), .B2(new_n296), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT28), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n255), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT31), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n279), .A2(new_n284), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n299), .A2(new_n307), .A3(KEYINPUT30), .A4(new_n327), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n263), .B(new_n328), .C1(new_n317), .C2(KEYINPUT30), .ZN(new_n329));
  INV_X1    g143(.A(new_n255), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n330), .B1(new_n309), .B2(new_n311), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT70), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n329), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AOI211_X1 g147(.A(KEYINPUT70), .B(new_n330), .C1(new_n309), .C2(new_n311), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n326), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n312), .A2(new_n255), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT70), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n331), .A2(new_n332), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n337), .A2(KEYINPUT31), .A3(new_n338), .A4(new_n329), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n325), .B1(new_n335), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(G472), .A2(G902), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT32), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n321), .A2(new_n324), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n330), .ZN(new_n345));
  INV_X1    g159(.A(new_n329), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n346), .B1(new_n336), .B2(KEYINPUT70), .ZN(new_n347));
  AOI21_X1  g161(.A(KEYINPUT31), .B1(new_n347), .B2(new_n338), .ZN(new_n348));
  NOR3_X1   g162(.A1(new_n333), .A2(new_n326), .A3(new_n334), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n345), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT32), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n351), .A3(new_n341), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n343), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G472), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n299), .A2(new_n307), .A3(new_n327), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n263), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n312), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT28), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n358), .A2(new_n324), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n255), .A2(KEYINPUT29), .ZN(new_n360));
  AOI21_X1  g174(.A(G902), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n312), .A2(new_n329), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT29), .B1(new_n362), .B2(new_n330), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n363), .B1(new_n344), .B2(new_n330), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n354), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n249), .B1(new_n353), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(KEYINPUT9), .B(G234), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n368), .B(KEYINPUT76), .ZN(new_n369));
  OAI21_X1  g183(.A(G221), .B1(new_n369), .B2(G902), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n279), .ZN(new_n372));
  INV_X1    g186(.A(G104), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT3), .B1(new_n373), .B2(G107), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT3), .ZN(new_n375));
  INV_X1    g189(.A(G107), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(G104), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n373), .A2(G107), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n374), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT4), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(G101), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT77), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n379), .A2(new_n382), .A3(G101), .ZN(new_n383));
  INV_X1    g197(.A(G101), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n374), .A2(new_n377), .A3(new_n384), .A4(new_n378), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n383), .A2(KEYINPUT4), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n382), .B1(new_n379), .B2(G101), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n284), .B(new_n381), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT10), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n373), .A2(G107), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n376), .A2(G104), .ZN(new_n391));
  OAI21_X1  g205(.A(G101), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n385), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n389), .B1(new_n296), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n393), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n305), .A2(KEYINPUT10), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n388), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT81), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n372), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n388), .A2(new_n394), .A3(KEYINPUT81), .A4(new_n396), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n388), .A2(new_n394), .A3(new_n372), .A4(new_n396), .ZN(new_n401));
  XNOR2_X1  g215(.A(G110), .B(G140), .ZN(new_n402));
  INV_X1    g216(.A(G227), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(G953), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n402), .B(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n401), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT80), .ZN(new_n408));
  AOI22_X1  g222(.A1(new_n399), .A2(new_n400), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n401), .A2(KEYINPUT80), .A3(new_n406), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT78), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n305), .A2(new_n395), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n393), .B1(new_n314), .B2(new_n302), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n411), .B(new_n279), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT79), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n415), .A3(KEYINPUT12), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n296), .A2(new_n393), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n305), .A2(new_n395), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n372), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT79), .B1(new_n419), .B2(new_n411), .ZN(new_n420));
  OAI211_X1 g234(.A(KEYINPUT79), .B(new_n279), .C1(new_n412), .C2(new_n413), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT12), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n401), .B(new_n416), .C1(new_n420), .C2(new_n423), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n409), .A2(new_n410), .B1(new_n424), .B2(new_n405), .ZN(new_n425));
  OAI21_X1  g239(.A(G469), .B1(new_n425), .B2(G902), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n414), .A2(new_n415), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(new_n422), .A3(new_n421), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n416), .ZN(new_n429));
  INV_X1    g243(.A(new_n401), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n430), .B1(new_n399), .B2(new_n400), .ZN(new_n431));
  OAI22_X1  g245(.A1(new_n429), .A2(new_n407), .B1(new_n431), .B2(new_n406), .ZN(new_n432));
  XOR2_X1   g246(.A(KEYINPUT82), .B(G469), .Z(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n235), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n371), .B1(new_n426), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n251), .A2(G143), .A3(G214), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(G143), .B1(new_n251), .B2(G214), .ZN(new_n438));
  AND2_X1   g252(.A1(KEYINPUT18), .A2(G131), .ZN(new_n439));
  OR3_X1    g253(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n251), .A2(G214), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n286), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n436), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n439), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n216), .B(new_n215), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n440), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  OR2_X1    g260(.A1(new_n205), .A2(new_n206), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(new_n209), .A3(new_n207), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n443), .A2(KEYINPUT17), .A3(G131), .ZN(new_n449));
  OAI21_X1  g263(.A(G131), .B1(new_n437), .B2(new_n438), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n442), .A2(new_n276), .A3(new_n436), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n449), .B1(new_n452), .B2(KEYINPUT17), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n446), .B1(new_n448), .B2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G113), .B(G122), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(G104), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G475), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n446), .A2(new_n456), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n216), .B(KEYINPUT19), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n215), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n462), .A2(new_n218), .A3(new_n220), .A4(new_n452), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n458), .A2(new_n459), .A3(new_n235), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT20), .ZN(new_n466));
  AOI22_X1  g280(.A1(new_n454), .A2(new_n457), .B1(new_n460), .B2(new_n463), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT20), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n467), .A2(new_n468), .A3(new_n459), .A4(new_n235), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G952), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n471), .A2(G953), .ZN(new_n472));
  INV_X1    g286(.A(G234), .ZN(new_n473));
  INV_X1    g287(.A(G237), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  AOI211_X1 g290(.A(new_n235), .B(new_n226), .C1(G234), .C2(G237), .ZN(new_n477));
  XNOR2_X1  g291(.A(KEYINPUT21), .B(G898), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  OR2_X1    g294(.A1(new_n457), .A2(KEYINPUT88), .ZN(new_n481));
  AOI21_X1  g295(.A(G902), .B1(new_n454), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n482), .B1(new_n454), .B2(new_n481), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G475), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n470), .A2(new_n480), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n286), .A2(G128), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n189), .A2(G143), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(new_n487), .A3(new_n270), .ZN(new_n488));
  INV_X1    g302(.A(G122), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(G116), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n257), .A2(G122), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n490), .A2(new_n491), .A3(new_n376), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n376), .B1(new_n490), .B2(new_n491), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n488), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT13), .B1(new_n286), .B2(G128), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n286), .A2(G128), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n286), .A2(KEYINPUT13), .A3(G128), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n270), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT89), .B1(new_n494), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n493), .ZN(new_n501));
  XNOR2_X1  g315(.A(G116), .B(G122), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n376), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT13), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n486), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(new_n498), .A3(new_n487), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G134), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT89), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n504), .A2(new_n508), .A3(new_n509), .A4(new_n488), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n500), .A2(new_n510), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n369), .A2(new_n242), .A3(G953), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n376), .B1(new_n490), .B2(KEYINPUT14), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(new_n502), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n486), .A2(new_n487), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(G134), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n516), .A2(KEYINPUT90), .A3(new_n488), .ZN(new_n517));
  AOI21_X1  g331(.A(KEYINPUT90), .B1(new_n516), .B2(new_n488), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n511), .A2(new_n512), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n512), .B1(new_n511), .B2(new_n519), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n235), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT91), .ZN(new_n523));
  INV_X1    g337(.A(G478), .ZN(new_n524));
  NOR2_X1   g338(.A1(KEYINPUT92), .A2(KEYINPUT15), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(KEYINPUT92), .A2(KEYINPUT15), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT91), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n529), .B(new_n235), .C1(new_n520), .C2(new_n521), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n523), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  OR2_X1    g345(.A1(new_n522), .A2(new_n528), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT93), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT93), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n531), .A2(new_n535), .A3(new_n532), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n485), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(G214), .B1(G237), .B2(G902), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(G210), .B1(G237), .B2(G902), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n284), .A2(G125), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n296), .B2(G125), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n226), .A2(G224), .ZN(new_n544));
  XOR2_X1   g358(.A(new_n544), .B(KEYINPUT84), .Z(new_n545));
  XNOR2_X1  g359(.A(new_n543), .B(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n256), .A2(new_n258), .A3(KEYINPUT5), .ZN(new_n548));
  OAI21_X1  g362(.A(G113), .B1(new_n256), .B2(KEYINPUT5), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n259), .A2(new_n260), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n395), .ZN(new_n553));
  XNOR2_X1  g367(.A(G110), .B(G122), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n386), .A2(new_n387), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n263), .A2(new_n381), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n553), .B(new_n554), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT6), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n553), .B1(new_n555), .B2(new_n556), .ZN(new_n559));
  XOR2_X1   g373(.A(G110), .B(G122), .Z(new_n560));
  AND2_X1   g374(.A1(new_n560), .A2(KEYINPUT83), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n559), .A2(KEYINPUT6), .A3(new_n561), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n547), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT85), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n554), .B(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n552), .A2(new_n393), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n548), .A2(KEYINPUT86), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(new_n549), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n548), .A2(KEYINPUT86), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n551), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n568), .B(new_n569), .C1(new_n573), .C2(new_n393), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT87), .ZN(new_n575));
  OAI211_X1 g389(.A(KEYINPUT7), .B(new_n544), .C1(new_n543), .C2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n305), .A2(new_n201), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n544), .A2(new_n575), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n544), .A2(KEYINPUT7), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n577), .A2(new_n542), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n574), .A2(new_n576), .A3(new_n557), .A4(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n235), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n541), .B1(new_n565), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n557), .A2(KEYINPUT6), .B1(new_n559), .B2(new_n561), .ZN(new_n584));
  INV_X1    g398(.A(new_n564), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n546), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n586), .A2(new_n235), .A3(new_n540), .A4(new_n581), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n539), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n435), .A2(new_n537), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n367), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(G101), .ZN(G3));
  NAND2_X1  g405(.A1(new_n350), .A2(new_n341), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n588), .A2(new_n480), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n470), .A2(new_n484), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n524), .A2(G902), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(KEYINPUT94), .B1(new_n520), .B2(new_n521), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT33), .ZN(new_n598));
  OR2_X1    g412(.A1(new_n512), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n598), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  OR2_X1    g415(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n597), .A2(new_n601), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n596), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n523), .A2(new_n524), .A3(new_n530), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n594), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n593), .A2(new_n607), .ZN(new_n608));
  AOI211_X1 g422(.A(new_n371), .B(new_n249), .C1(new_n426), .C2(new_n434), .ZN(new_n609));
  OAI21_X1  g423(.A(G472), .B1(new_n340), .B2(G902), .ZN(new_n610));
  AND4_X1   g424(.A1(new_n592), .A2(new_n608), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(new_n373), .ZN(new_n612));
  XNOR2_X1  g426(.A(KEYINPUT95), .B(KEYINPUT34), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G6));
  AND2_X1   g428(.A1(new_n610), .A2(new_n592), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT96), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n470), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n466), .A2(new_n469), .A3(KEYINPUT96), .ZN(new_n618));
  AOI22_X1  g432(.A1(new_n617), .A2(new_n618), .B1(G475), .B2(new_n483), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n619), .A2(new_n536), .A3(new_n534), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n620), .A2(new_n593), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n615), .A2(new_n609), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT35), .B(G107), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G9));
  NAND2_X1  g438(.A1(new_n610), .A2(new_n592), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT36), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n225), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n626), .A2(new_n224), .A3(new_n211), .A4(new_n223), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n628), .A2(new_n247), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT97), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT98), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n631), .A2(new_n632), .A3(new_n245), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n632), .B1(new_n631), .B2(new_n245), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n635), .A2(new_n435), .A3(new_n537), .A4(new_n588), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n625), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT37), .B(G110), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G12));
  AOI21_X1  g453(.A(new_n351), .B1(new_n350), .B2(new_n341), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n340), .A2(KEYINPUT32), .A3(new_n342), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n366), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n635), .A2(new_n435), .A3(new_n588), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(G900), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n476), .B1(new_n477), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n620), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n642), .A2(new_n644), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G128), .ZN(G30));
  XOR2_X1   g463(.A(new_n646), .B(KEYINPUT39), .Z(new_n650));
  NAND2_X1  g464(.A1(new_n435), .A2(new_n650), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n651), .A2(KEYINPUT40), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n583), .A2(new_n587), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n631), .A2(new_n245), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n539), .B1(new_n470), .B2(new_n484), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n534), .A2(new_n536), .A3(new_n657), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n655), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n652), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(KEYINPUT40), .B2(new_n651), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n357), .A2(new_n330), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n662), .B1(new_n333), .B2(new_n334), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT100), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI211_X1 g479(.A(KEYINPUT100), .B(new_n662), .C1(new_n333), .C2(new_n334), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n665), .A2(new_n235), .A3(new_n666), .ZN(new_n667));
  AOI221_X4 g481(.A(KEYINPUT101), .B1(G472), .B2(new_n667), .C1(new_n343), .C2(new_n352), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT101), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n667), .A2(G472), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n669), .B1(new_n353), .B2(new_n670), .ZN(new_n671));
  OR2_X1    g485(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n661), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G143), .ZN(G45));
  NOR2_X1   g488(.A1(new_n607), .A2(new_n646), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n642), .A2(new_n644), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G146), .ZN(G48));
  INV_X1    g491(.A(new_n249), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n432), .A2(new_n235), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(G469), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n680), .A2(new_n370), .A3(new_n434), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n681), .A2(new_n593), .A3(new_n607), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n642), .A2(new_n678), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT41), .B(G113), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G15));
  NOR3_X1   g499(.A1(new_n620), .A2(new_n681), .A3(new_n593), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n642), .A2(new_n678), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G116), .ZN(G18));
  NAND2_X1  g502(.A1(new_n635), .A2(new_n537), .ZN(new_n689));
  INV_X1    g503(.A(new_n588), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n689), .A2(new_n690), .A3(new_n681), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n642), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G119), .ZN(G21));
  NAND2_X1  g507(.A1(new_n358), .A2(new_n324), .ZN(new_n694));
  AOI22_X1  g508(.A1(new_n335), .A2(new_n339), .B1(new_n330), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g509(.A(KEYINPUT102), .B1(new_n695), .B2(new_n342), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n694), .A2(new_n330), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n697), .B1(new_n348), .B2(new_n349), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT102), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n698), .A2(new_n699), .A3(new_n341), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n610), .A2(new_n696), .A3(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n534), .A2(new_n653), .A3(new_n657), .A4(new_n536), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n681), .A2(new_n702), .A3(new_n479), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n701), .A2(new_n678), .A3(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(KEYINPUT103), .B(G122), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G24));
  NOR2_X1   g520(.A1(new_n681), .A2(new_n690), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n701), .A2(new_n656), .A3(new_n675), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G125), .ZN(G27));
  NOR2_X1   g523(.A1(new_n653), .A2(new_n539), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n675), .A2(new_n435), .A3(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g526(.A(KEYINPUT42), .B1(new_n367), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n365), .B1(new_n343), .B2(new_n352), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT42), .ZN(new_n715));
  NOR4_X1   g529(.A1(new_n714), .A2(new_n715), .A3(new_n711), .A4(new_n249), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n713), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n642), .A2(new_n678), .A3(new_n712), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n715), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n367), .A2(KEYINPUT42), .A3(new_n712), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT104), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G131), .ZN(G33));
  NAND2_X1  g538(.A1(new_n435), .A2(new_n710), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n725), .A2(new_n620), .A3(new_n646), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n367), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G134), .ZN(G36));
  INV_X1    g542(.A(G469), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n235), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT105), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n399), .A2(new_n400), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n407), .A2(new_n408), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(new_n410), .A3(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n424), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n734), .B1(new_n735), .B2(new_n406), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT45), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n731), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n425), .A2(KEYINPUT105), .A3(KEYINPUT45), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n729), .B1(new_n736), .B2(new_n737), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n730), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n742), .A2(KEYINPUT46), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n434), .B1(new_n742), .B2(KEYINPUT46), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n370), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n746));
  INV_X1    g560(.A(new_n650), .ZN(new_n747));
  OR3_X1    g561(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n746), .B1(new_n745), .B2(new_n747), .ZN(new_n749));
  INV_X1    g563(.A(new_n604), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n605), .ZN(new_n751));
  INV_X1    g565(.A(new_n594), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT43), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(new_n625), .A3(new_n656), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n756), .A2(KEYINPUT44), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(KEYINPUT44), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n710), .B(KEYINPUT107), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n748), .A2(new_n749), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G137), .ZN(G39));
  INV_X1    g576(.A(new_n675), .ZN(new_n763));
  INV_X1    g577(.A(new_n710), .ZN(new_n764));
  NOR4_X1   g578(.A1(new_n642), .A2(new_n678), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n745), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n370), .B(new_n766), .C1(new_n743), .C2(new_n744), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n765), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G140), .ZN(G42));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n635), .A2(new_n435), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n533), .A2(new_n646), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n710), .A2(new_n619), .A3(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n710), .A2(new_n619), .A3(KEYINPUT112), .A4(new_n777), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n776), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AOI22_X1  g596(.A1(new_n367), .A2(new_n726), .B1(new_n782), .B2(new_n642), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n615), .A2(new_n589), .A3(new_n635), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n752), .A2(new_n533), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n593), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n615), .A2(new_n609), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT111), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n784), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n611), .B1(new_n367), .B2(new_n589), .ZN(new_n790));
  AND4_X1   g604(.A1(new_n592), .A2(new_n786), .A3(new_n609), .A4(new_n610), .ZN(new_n791));
  OAI21_X1  g605(.A(KEYINPUT111), .B1(new_n791), .B2(new_n637), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n783), .A2(new_n789), .A3(new_n790), .A4(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n610), .A2(new_n696), .A3(new_n700), .A4(new_n656), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n763), .ZN(new_n796));
  INV_X1    g610(.A(new_n725), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n794), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR4_X1   g612(.A1(new_n795), .A2(KEYINPUT113), .A3(new_n763), .A4(new_n725), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n793), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n683), .A2(new_n704), .A3(new_n687), .A4(new_n692), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT110), .ZN(new_n803));
  AOI22_X1  g617(.A1(new_n367), .A2(new_n682), .B1(new_n691), .B2(new_n642), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT110), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n804), .A2(new_n805), .A3(new_n687), .A4(new_n704), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n801), .A2(new_n723), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n435), .ZN(new_n809));
  NOR4_X1   g623(.A1(new_n809), .A2(new_n702), .A3(new_n656), .A4(new_n646), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n810), .B1(new_n668), .B2(new_n671), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n811), .A2(new_n648), .A3(new_n676), .A4(new_n708), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n708), .A2(new_n648), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(KEYINPUT52), .A3(new_n811), .A4(new_n676), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n775), .B1(new_n808), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT53), .B1(new_n713), .B2(new_n716), .ZN(new_n819));
  NOR4_X1   g633(.A1(new_n793), .A2(new_n800), .A3(new_n819), .A4(new_n802), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n708), .A2(new_n648), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT114), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n708), .A2(new_n648), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n822), .A2(new_n676), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n811), .A2(KEYINPUT52), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n814), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n820), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n818), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n774), .B1(new_n829), .B2(KEYINPUT54), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n814), .A2(new_n816), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n723), .A3(new_n801), .A4(new_n807), .ZN(new_n832));
  AOI22_X1  g646(.A1(new_n832), .A2(new_n775), .B1(new_n827), .B2(new_n820), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n833), .A2(KEYINPUT115), .A3(new_n834), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n801), .A2(new_n723), .A3(new_n807), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(new_n775), .A3(new_n827), .ZN(new_n837));
  INV_X1    g651(.A(new_n832), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n837), .B(KEYINPUT54), .C1(new_n838), .C2(new_n775), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n830), .A2(new_n835), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n367), .ZN(new_n841));
  INV_X1    g655(.A(new_n681), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n710), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n475), .B1(new_n843), .B2(KEYINPUT117), .ZN(new_n844));
  OR3_X1    g658(.A1(new_n681), .A2(new_n764), .A3(KEYINPUT117), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n844), .A2(new_n755), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n844), .A2(KEYINPUT118), .A3(new_n755), .A4(new_n845), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n841), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT48), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT120), .ZN(new_n852));
  OR2_X1    g666(.A1(new_n851), .A2(KEYINPUT120), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n850), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n854), .B1(new_n850), .B2(new_n852), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n678), .A2(new_n701), .A3(new_n755), .A4(new_n476), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n707), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT119), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n672), .A2(new_n249), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n844), .A2(new_n845), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n859), .A2(new_n594), .A3(new_n751), .A4(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n858), .A2(new_n472), .A3(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n855), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT51), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT50), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n842), .A2(new_n655), .A3(new_n539), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n856), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n865), .B1(new_n856), .B2(new_n866), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n751), .A2(new_n594), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n859), .A2(new_n860), .A3(new_n870), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n848), .A2(new_n849), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n869), .B(new_n871), .C1(new_n795), .C2(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n680), .A2(new_n434), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT109), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n768), .B(new_n770), .C1(new_n370), .C2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n856), .A2(new_n760), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT116), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT116), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n856), .A2(new_n879), .A3(new_n760), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n876), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n864), .B1(new_n873), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n863), .A2(new_n882), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n873), .A2(new_n881), .A3(new_n864), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI22_X1  g699(.A1(new_n840), .A2(new_n885), .B1(G952), .B2(G953), .ZN(new_n886));
  INV_X1    g700(.A(new_n753), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n655), .A2(new_n887), .A3(new_n370), .A4(new_n538), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(new_n875), .B2(KEYINPUT49), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n859), .B(new_n889), .C1(KEYINPUT49), .C2(new_n875), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n886), .A2(new_n890), .ZN(G75));
  INV_X1    g705(.A(KEYINPUT56), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n829), .A2(G902), .ZN(new_n893));
  INV_X1    g707(.A(G210), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n584), .A2(new_n585), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(new_n546), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT55), .Z(new_n898));
  NAND2_X1  g712(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n898), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n892), .B(new_n900), .C1(new_n893), .C2(new_n894), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n226), .A2(G952), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n899), .A2(new_n901), .A3(new_n903), .ZN(G51));
  XNOR2_X1  g718(.A(new_n730), .B(KEYINPUT57), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n818), .A2(new_n834), .A3(new_n828), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n834), .B1(new_n818), .B2(new_n828), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n432), .ZN(new_n909));
  INV_X1    g723(.A(new_n893), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n910), .A2(new_n740), .A3(new_n741), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n902), .B1(new_n909), .B2(new_n911), .ZN(G54));
  AND2_X1   g726(.A1(KEYINPUT58), .A2(G475), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n910), .A2(new_n467), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n467), .B1(new_n910), .B2(new_n913), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n914), .A2(new_n915), .A3(new_n902), .ZN(G60));
  NAND2_X1  g730(.A1(G478), .A2(G902), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT59), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n602), .A2(new_n603), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT121), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n918), .B(new_n920), .C1(new_n906), .C2(new_n907), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n903), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n840), .A2(new_n918), .ZN(new_n923));
  INV_X1    g737(.A(new_n920), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(G63));
  INV_X1    g739(.A(new_n246), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n241), .B(KEYINPUT60), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n926), .B1(new_n833), .B2(new_n927), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n628), .A2(new_n629), .ZN(new_n929));
  INV_X1    g743(.A(new_n927), .ZN(new_n930));
  AOI21_X1  g744(.A(KEYINPUT53), .B1(new_n836), .B2(new_n831), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n820), .A2(new_n827), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n929), .B(new_n930), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n928), .A2(new_n933), .A3(new_n903), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT122), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n933), .A2(new_n935), .A3(new_n903), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n934), .A2(new_n936), .A3(KEYINPUT61), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n927), .B1(new_n818), .B2(new_n828), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n902), .B1(new_n938), .B2(new_n929), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT61), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n939), .B(new_n928), .C1(new_n935), .C2(new_n940), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n937), .A2(new_n941), .ZN(G66));
  AND2_X1   g756(.A1(new_n790), .A2(new_n792), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n807), .A2(new_n789), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(G224), .A2(G953), .ZN(new_n945));
  OAI22_X1  g759(.A1(new_n944), .A2(G953), .B1(new_n478), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n896), .B1(G898), .B2(new_n226), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n946), .B(new_n947), .Z(G69));
  INV_X1    g762(.A(KEYINPUT123), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n328), .B1(new_n317), .B2(KEYINPUT30), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(new_n461), .Z(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n825), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n953), .A2(KEYINPUT62), .A3(new_n673), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n955));
  INV_X1    g769(.A(new_n673), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n955), .B1(new_n825), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n764), .B1(new_n785), .B2(new_n607), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n367), .A2(new_n435), .A3(new_n650), .A4(new_n959), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n761), .A2(new_n772), .A3(new_n960), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n949), .B(new_n952), .C1(new_n962), .C2(G953), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n952), .B1(G900), .B2(G953), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n841), .A2(new_n702), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n748), .A2(new_n749), .A3(new_n965), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT124), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n723), .A2(new_n772), .A3(new_n727), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n967), .A2(new_n968), .A3(new_n761), .A4(new_n953), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n964), .B1(new_n969), .B2(G953), .ZN(new_n970));
  AOI21_X1  g784(.A(G953), .B1(new_n958), .B2(new_n961), .ZN(new_n971));
  OAI21_X1  g785(.A(KEYINPUT123), .B1(new_n971), .B2(new_n951), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n963), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(G953), .B1(new_n403), .B2(new_n645), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT125), .Z(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n963), .A2(new_n970), .A3(new_n972), .A4(new_n975), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(G72));
  NAND2_X1  g793(.A1(G472), .A2(G902), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT63), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT126), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n982), .B1(new_n969), .B2(new_n944), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n362), .A2(new_n255), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n362), .A2(new_n255), .ZN(new_n986));
  INV_X1    g800(.A(new_n944), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n962), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n986), .B1(new_n988), .B2(new_n982), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n837), .B1(new_n838), .B2(new_n775), .ZN(new_n990));
  AOI22_X1  g804(.A1(new_n347), .A2(new_n338), .B1(new_n330), .B2(new_n362), .ZN(new_n991));
  NOR3_X1   g805(.A1(new_n990), .A2(new_n981), .A3(new_n991), .ZN(new_n992));
  NOR4_X1   g806(.A1(new_n985), .A2(new_n989), .A3(new_n992), .A4(new_n902), .ZN(G57));
endmodule


