

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U550 ( .A1(G8), .A2(n664), .ZN(n705) );
  OR2_X2 U551 ( .A1(n537), .A2(n555), .ZN(n535) );
  NOR2_X2 U552 ( .A1(G2104), .A2(n530), .ZN(n879) );
  NAND2_X1 U553 ( .A1(n720), .A2(n593), .ZN(n664) );
  NOR2_X2 U554 ( .A1(n530), .A2(n547), .ZN(n878) );
  INV_X1 U555 ( .A(G2104), .ZN(n547) );
  NOR2_X1 U556 ( .A1(n614), .A2(n613), .ZN(n616) );
  OR2_X1 U557 ( .A1(n629), .A2(n781), .ZN(n628) );
  NOR2_X1 U558 ( .A1(G651), .A2(G543), .ZN(n541) );
  XNOR2_X2 U559 ( .A(KEYINPUT69), .B(n535), .ZN(n601) );
  OR2_X1 U560 ( .A1(n696), .A2(n695), .ZN(n515) );
  AND2_X1 U561 ( .A1(n742), .A2(n741), .ZN(n516) );
  XOR2_X1 U562 ( .A(KEYINPUT23), .B(n526), .Z(n517) );
  AND2_X1 U563 ( .A1(n758), .A2(n976), .ZN(n518) );
  XOR2_X1 U564 ( .A(n707), .B(KEYINPUT92), .Z(n519) );
  AND2_X1 U565 ( .A1(n708), .A2(n519), .ZN(n520) );
  OR2_X1 U566 ( .A1(n612), .A2(n1015), .ZN(n613) );
  INV_X1 U567 ( .A(KEYINPUT64), .ZN(n615) );
  XNOR2_X1 U568 ( .A(n616), .B(n615), .ZN(n629) );
  NOR2_X1 U569 ( .A1(n740), .A2(n518), .ZN(n741) );
  XNOR2_X1 U570 ( .A(KEYINPUT12), .B(KEYINPUT72), .ZN(n599) );
  NOR2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n528) );
  INV_X1 U572 ( .A(KEYINPUT101), .ZN(n743) );
  XNOR2_X1 U573 ( .A(n600), .B(n599), .ZN(n603) );
  NOR2_X1 U574 ( .A1(n534), .A2(n533), .ZN(n592) );
  BUF_X1 U575 ( .A(n592), .Z(G160) );
  INV_X1 U576 ( .A(G2105), .ZN(n530) );
  NAND2_X1 U577 ( .A1(G113), .A2(n878), .ZN(n521) );
  XNOR2_X1 U578 ( .A(n521), .B(KEYINPUT68), .ZN(n527) );
  XOR2_X1 U579 ( .A(KEYINPUT67), .B(KEYINPUT66), .Z(n525) );
  INV_X1 U580 ( .A(G101), .ZN(n522) );
  NOR2_X1 U581 ( .A1(n547), .A2(n522), .ZN(n523) );
  NAND2_X1 U582 ( .A1(n530), .A2(n523), .ZN(n524) );
  XNOR2_X1 U583 ( .A(n525), .B(n524), .ZN(n526) );
  NAND2_X1 U584 ( .A1(n527), .A2(n517), .ZN(n534) );
  XOR2_X1 U585 ( .A(KEYINPUT17), .B(n528), .Z(n529) );
  BUF_X2 U586 ( .A(n529), .Z(n874) );
  NAND2_X1 U587 ( .A1(G137), .A2(n874), .ZN(n532) );
  NAND2_X1 U588 ( .A1(G125), .A2(n879), .ZN(n531) );
  NAND2_X1 U589 ( .A1(n532), .A2(n531), .ZN(n533) );
  INV_X1 U590 ( .A(G651), .ZN(n537) );
  XOR2_X1 U591 ( .A(KEYINPUT0), .B(G543), .Z(n555) );
  NAND2_X1 U592 ( .A1(G73), .A2(n601), .ZN(n536) );
  XNOR2_X1 U593 ( .A(n536), .B(KEYINPUT2), .ZN(n546) );
  NOR2_X1 U594 ( .A1(G543), .A2(n537), .ZN(n538) );
  XOR2_X1 U595 ( .A(KEYINPUT1), .B(n538), .Z(n605) );
  BUF_X1 U596 ( .A(n605), .Z(n790) );
  NAND2_X1 U597 ( .A1(G61), .A2(n790), .ZN(n540) );
  NOR2_X2 U598 ( .A1(G651), .A2(n555), .ZN(n794) );
  NAND2_X1 U599 ( .A1(G48), .A2(n794), .ZN(n539) );
  NAND2_X1 U600 ( .A1(n540), .A2(n539), .ZN(n544) );
  XOR2_X2 U601 ( .A(KEYINPUT65), .B(n541), .Z(n787) );
  NAND2_X1 U602 ( .A1(G86), .A2(n787), .ZN(n542) );
  XNOR2_X1 U603 ( .A(KEYINPUT79), .B(n542), .ZN(n543) );
  NOR2_X1 U604 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U605 ( .A1(n546), .A2(n545), .ZN(G305) );
  NAND2_X1 U606 ( .A1(G138), .A2(n874), .ZN(n549) );
  NOR2_X1 U607 ( .A1(G2105), .A2(n547), .ZN(n875) );
  NAND2_X1 U608 ( .A1(G102), .A2(n875), .ZN(n548) );
  NAND2_X1 U609 ( .A1(n549), .A2(n548), .ZN(n553) );
  NAND2_X1 U610 ( .A1(G114), .A2(n878), .ZN(n551) );
  NAND2_X1 U611 ( .A1(G126), .A2(n879), .ZN(n550) );
  NAND2_X1 U612 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U613 ( .A1(n553), .A2(n552), .ZN(G164) );
  NAND2_X1 U614 ( .A1(G49), .A2(n794), .ZN(n554) );
  XNOR2_X1 U615 ( .A(n554), .B(KEYINPUT78), .ZN(n560) );
  NAND2_X1 U616 ( .A1(G87), .A2(n555), .ZN(n557) );
  NAND2_X1 U617 ( .A1(G74), .A2(G651), .ZN(n556) );
  NAND2_X1 U618 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U619 ( .A1(n790), .A2(n558), .ZN(n559) );
  NAND2_X1 U620 ( .A1(n560), .A2(n559), .ZN(G288) );
  NAND2_X1 U621 ( .A1(G64), .A2(n790), .ZN(n562) );
  NAND2_X1 U622 ( .A1(G52), .A2(n794), .ZN(n561) );
  NAND2_X1 U623 ( .A1(n562), .A2(n561), .ZN(n568) );
  NAND2_X1 U624 ( .A1(G90), .A2(n787), .ZN(n564) );
  NAND2_X1 U625 ( .A1(G77), .A2(n601), .ZN(n563) );
  NAND2_X1 U626 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U627 ( .A(KEYINPUT70), .B(n565), .Z(n566) );
  XNOR2_X1 U628 ( .A(KEYINPUT9), .B(n566), .ZN(n567) );
  NOR2_X1 U629 ( .A1(n568), .A2(n567), .ZN(G171) );
  INV_X1 U630 ( .A(G171), .ZN(G301) );
  NAND2_X1 U631 ( .A1(n787), .A2(G89), .ZN(n569) );
  XNOR2_X1 U632 ( .A(n569), .B(KEYINPUT4), .ZN(n571) );
  NAND2_X1 U633 ( .A1(G76), .A2(n601), .ZN(n570) );
  NAND2_X1 U634 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U635 ( .A(n572), .B(KEYINPUT5), .ZN(n577) );
  NAND2_X1 U636 ( .A1(G63), .A2(n790), .ZN(n574) );
  NAND2_X1 U637 ( .A1(G51), .A2(n794), .ZN(n573) );
  NAND2_X1 U638 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U639 ( .A(KEYINPUT6), .B(n575), .Z(n576) );
  NAND2_X1 U640 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U641 ( .A(n578), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U642 ( .A1(G88), .A2(n787), .ZN(n580) );
  NAND2_X1 U643 ( .A1(G75), .A2(n601), .ZN(n579) );
  NAND2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n584) );
  NAND2_X1 U645 ( .A1(G62), .A2(n790), .ZN(n582) );
  NAND2_X1 U646 ( .A1(G50), .A2(n794), .ZN(n581) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(G166) );
  XOR2_X1 U649 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U650 ( .A(G166), .ZN(G303) );
  AND2_X1 U651 ( .A1(n601), .A2(G72), .ZN(n588) );
  NAND2_X1 U652 ( .A1(G85), .A2(n787), .ZN(n586) );
  NAND2_X1 U653 ( .A1(G47), .A2(n794), .ZN(n585) );
  NAND2_X1 U654 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U655 ( .A1(n588), .A2(n587), .ZN(n590) );
  NAND2_X1 U656 ( .A1(n790), .A2(G60), .ZN(n589) );
  NAND2_X1 U657 ( .A1(n590), .A2(n589), .ZN(G290) );
  XOR2_X1 U658 ( .A(KEYINPUT100), .B(G1981), .Z(n591) );
  XNOR2_X1 U659 ( .A(G305), .B(n591), .ZN(n1001) );
  NOR2_X1 U660 ( .A1(G164), .A2(G1384), .ZN(n720) );
  NAND2_X1 U661 ( .A1(n592), .A2(G40), .ZN(n719) );
  INV_X1 U662 ( .A(n719), .ZN(n593) );
  NOR2_X1 U663 ( .A1(G1976), .A2(G288), .ZN(n687) );
  NAND2_X1 U664 ( .A1(n687), .A2(KEYINPUT33), .ZN(n594) );
  NOR2_X1 U665 ( .A1(n705), .A2(n594), .ZN(n595) );
  XNOR2_X1 U666 ( .A(n595), .B(KEYINPUT99), .ZN(n596) );
  NAND2_X1 U667 ( .A1(n1001), .A2(n596), .ZN(n696) );
  INV_X1 U668 ( .A(G1996), .ZN(n597) );
  NOR2_X1 U669 ( .A1(n664), .A2(n597), .ZN(n598) );
  XNOR2_X1 U670 ( .A(n598), .B(KEYINPUT26), .ZN(n614) );
  AND2_X1 U671 ( .A1(n664), .A2(G1341), .ZN(n612) );
  NAND2_X1 U672 ( .A1(G81), .A2(n787), .ZN(n600) );
  NAND2_X1 U673 ( .A1(G68), .A2(n601), .ZN(n602) );
  NAND2_X1 U674 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U675 ( .A(KEYINPUT13), .B(n604), .ZN(n611) );
  NAND2_X1 U676 ( .A1(G56), .A2(n605), .ZN(n606) );
  XOR2_X1 U677 ( .A(KEYINPUT14), .B(n606), .Z(n609) );
  NAND2_X1 U678 ( .A1(G43), .A2(n794), .ZN(n607) );
  XNOR2_X1 U679 ( .A(KEYINPUT73), .B(n607), .ZN(n608) );
  NOR2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U681 ( .A1(n611), .A2(n610), .ZN(n1015) );
  NAND2_X1 U682 ( .A1(n790), .A2(G66), .ZN(n623) );
  NAND2_X1 U683 ( .A1(G92), .A2(n787), .ZN(n618) );
  NAND2_X1 U684 ( .A1(G79), .A2(n601), .ZN(n617) );
  NAND2_X1 U685 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U686 ( .A1(G54), .A2(n794), .ZN(n619) );
  XNOR2_X1 U687 ( .A(KEYINPUT75), .B(n619), .ZN(n620) );
  NOR2_X1 U688 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U689 ( .A1(n623), .A2(n622), .ZN(n624) );
  XOR2_X1 U690 ( .A(KEYINPUT15), .B(n624), .Z(n781) );
  INV_X1 U691 ( .A(n664), .ZN(n649) );
  NOR2_X1 U692 ( .A1(n649), .A2(G1348), .ZN(n626) );
  NOR2_X1 U693 ( .A1(G2067), .A2(n664), .ZN(n625) );
  NOR2_X1 U694 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U695 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U696 ( .A1(n629), .A2(n781), .ZN(n630) );
  NAND2_X1 U697 ( .A1(n631), .A2(n630), .ZN(n642) );
  NAND2_X1 U698 ( .A1(G65), .A2(n790), .ZN(n633) );
  NAND2_X1 U699 ( .A1(G53), .A2(n794), .ZN(n632) );
  NAND2_X1 U700 ( .A1(n633), .A2(n632), .ZN(n637) );
  NAND2_X1 U701 ( .A1(G91), .A2(n787), .ZN(n635) );
  NAND2_X1 U702 ( .A1(G78), .A2(n601), .ZN(n634) );
  NAND2_X1 U703 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U704 ( .A1(n637), .A2(n636), .ZN(n1004) );
  NAND2_X1 U705 ( .A1(n649), .A2(G2072), .ZN(n638) );
  XNOR2_X1 U706 ( .A(n638), .B(KEYINPUT27), .ZN(n640) );
  INV_X1 U707 ( .A(G1956), .ZN(n1005) );
  NOR2_X1 U708 ( .A1(n1005), .A2(n649), .ZN(n639) );
  NOR2_X1 U709 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U710 ( .A1(n1004), .A2(n643), .ZN(n641) );
  NAND2_X1 U711 ( .A1(n642), .A2(n641), .ZN(n646) );
  NOR2_X1 U712 ( .A1(n1004), .A2(n643), .ZN(n644) );
  XOR2_X1 U713 ( .A(n644), .B(KEYINPUT28), .Z(n645) );
  NAND2_X1 U714 ( .A1(n646), .A2(n645), .ZN(n648) );
  XOR2_X1 U715 ( .A(KEYINPUT29), .B(KEYINPUT94), .Z(n647) );
  XNOR2_X1 U716 ( .A(n648), .B(n647), .ZN(n653) );
  XOR2_X1 U717 ( .A(KEYINPUT25), .B(G2078), .Z(n956) );
  NOR2_X1 U718 ( .A1(n956), .A2(n664), .ZN(n651) );
  NOR2_X1 U719 ( .A1(n649), .A2(G1961), .ZN(n650) );
  NOR2_X1 U720 ( .A1(n651), .A2(n650), .ZN(n659) );
  OR2_X1 U721 ( .A1(n659), .A2(G301), .ZN(n652) );
  NAND2_X1 U722 ( .A1(n653), .A2(n652), .ZN(n678) );
  NOR2_X1 U723 ( .A1(G2084), .A2(n664), .ZN(n679) );
  NOR2_X1 U724 ( .A1(n705), .A2(G1966), .ZN(n654) );
  XNOR2_X1 U725 ( .A(n654), .B(KEYINPUT93), .ZN(n681) );
  NAND2_X1 U726 ( .A1(G8), .A2(n681), .ZN(n655) );
  NOR2_X1 U727 ( .A1(n679), .A2(n655), .ZN(n656) );
  XNOR2_X1 U728 ( .A(KEYINPUT30), .B(n656), .ZN(n658) );
  INV_X1 U729 ( .A(G168), .ZN(n657) );
  NAND2_X1 U730 ( .A1(n658), .A2(n657), .ZN(n661) );
  NAND2_X1 U731 ( .A1(n659), .A2(G301), .ZN(n660) );
  NAND2_X1 U732 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U733 ( .A(n662), .B(KEYINPUT31), .ZN(n677) );
  INV_X1 U734 ( .A(G8), .ZN(n669) );
  NOR2_X1 U735 ( .A1(G1971), .A2(n705), .ZN(n663) );
  XNOR2_X1 U736 ( .A(KEYINPUT95), .B(n663), .ZN(n667) );
  NOR2_X1 U737 ( .A1(G2090), .A2(n664), .ZN(n665) );
  NOR2_X1 U738 ( .A1(G166), .A2(n665), .ZN(n666) );
  NAND2_X1 U739 ( .A1(n667), .A2(n666), .ZN(n668) );
  OR2_X1 U740 ( .A1(n669), .A2(n668), .ZN(n671) );
  AND2_X1 U741 ( .A1(n677), .A2(n671), .ZN(n670) );
  NAND2_X1 U742 ( .A1(n678), .A2(n670), .ZN(n675) );
  INV_X1 U743 ( .A(n671), .ZN(n673) );
  AND2_X1 U744 ( .A1(G286), .A2(G8), .ZN(n672) );
  OR2_X1 U745 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U746 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U747 ( .A(n676), .B(KEYINPUT32), .ZN(n697) );
  NAND2_X1 U748 ( .A1(n678), .A2(n677), .ZN(n683) );
  NAND2_X1 U749 ( .A1(G8), .A2(n679), .ZN(n680) );
  AND2_X1 U750 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U751 ( .A1(n683), .A2(n682), .ZN(n698) );
  NAND2_X1 U752 ( .A1(G288), .A2(G1976), .ZN(n684) );
  XNOR2_X1 U753 ( .A(n684), .B(KEYINPUT96), .ZN(n1014) );
  AND2_X1 U754 ( .A1(n698), .A2(n1014), .ZN(n685) );
  NAND2_X1 U755 ( .A1(n697), .A2(n685), .ZN(n690) );
  INV_X1 U756 ( .A(n1014), .ZN(n688) );
  NOR2_X1 U757 ( .A1(G1971), .A2(G303), .ZN(n686) );
  NOR2_X1 U758 ( .A1(n687), .A2(n686), .ZN(n1010) );
  OR2_X1 U759 ( .A1(n688), .A2(n1010), .ZN(n689) );
  NAND2_X1 U760 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U761 ( .A(n691), .B(KEYINPUT97), .ZN(n692) );
  NOR2_X1 U762 ( .A1(n705), .A2(n692), .ZN(n693) );
  NOR2_X1 U763 ( .A1(n693), .A2(KEYINPUT33), .ZN(n694) );
  XNOR2_X1 U764 ( .A(n694), .B(KEYINPUT98), .ZN(n695) );
  NAND2_X1 U765 ( .A1(n698), .A2(n697), .ZN(n701) );
  NOR2_X1 U766 ( .A1(G2090), .A2(G303), .ZN(n699) );
  NAND2_X1 U767 ( .A1(G8), .A2(n699), .ZN(n700) );
  NAND2_X1 U768 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U769 ( .A1(n705), .A2(n702), .ZN(n708) );
  NOR2_X1 U770 ( .A1(G1981), .A2(G305), .ZN(n703) );
  XNOR2_X1 U771 ( .A(n703), .B(KEYINPUT24), .ZN(n704) );
  XNOR2_X1 U772 ( .A(n704), .B(KEYINPUT91), .ZN(n706) );
  NOR2_X1 U773 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U774 ( .A1(n515), .A2(n520), .ZN(n742) );
  NAND2_X1 U775 ( .A1(G116), .A2(n878), .ZN(n710) );
  NAND2_X1 U776 ( .A1(G128), .A2(n879), .ZN(n709) );
  NAND2_X1 U777 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U778 ( .A(n711), .B(KEYINPUT35), .ZN(n716) );
  NAND2_X1 U779 ( .A1(G140), .A2(n874), .ZN(n713) );
  NAND2_X1 U780 ( .A1(G104), .A2(n875), .ZN(n712) );
  NAND2_X1 U781 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U782 ( .A(KEYINPUT34), .B(n714), .Z(n715) );
  NAND2_X1 U783 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U784 ( .A(n717), .B(KEYINPUT36), .Z(n887) );
  XNOR2_X1 U785 ( .A(G2067), .B(KEYINPUT37), .ZN(n756) );
  OR2_X1 U786 ( .A1(n887), .A2(n756), .ZN(n718) );
  XOR2_X1 U787 ( .A(KEYINPUT86), .B(n718), .Z(n989) );
  NOR2_X1 U788 ( .A1(n720), .A2(n719), .ZN(n758) );
  NAND2_X1 U789 ( .A1(n989), .A2(n758), .ZN(n721) );
  XOR2_X1 U790 ( .A(KEYINPUT87), .B(n721), .Z(n754) );
  INV_X1 U791 ( .A(n754), .ZN(n740) );
  NAND2_X1 U792 ( .A1(n879), .A2(G129), .ZN(n722) );
  XOR2_X1 U793 ( .A(KEYINPUT89), .B(n722), .Z(n724) );
  NAND2_X1 U794 ( .A1(n878), .A2(G117), .ZN(n723) );
  NAND2_X1 U795 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U796 ( .A(KEYINPUT90), .B(n725), .ZN(n728) );
  NAND2_X1 U797 ( .A1(n875), .A2(G105), .ZN(n726) );
  XOR2_X1 U798 ( .A(KEYINPUT38), .B(n726), .Z(n727) );
  NOR2_X1 U799 ( .A1(n728), .A2(n727), .ZN(n730) );
  NAND2_X1 U800 ( .A1(n874), .A2(G141), .ZN(n729) );
  NAND2_X1 U801 ( .A1(n730), .A2(n729), .ZN(n893) );
  NAND2_X1 U802 ( .A1(G1996), .A2(n893), .ZN(n739) );
  NAND2_X1 U803 ( .A1(G131), .A2(n874), .ZN(n732) );
  NAND2_X1 U804 ( .A1(G95), .A2(n875), .ZN(n731) );
  NAND2_X1 U805 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U806 ( .A(KEYINPUT88), .B(n733), .Z(n737) );
  NAND2_X1 U807 ( .A1(G107), .A2(n878), .ZN(n735) );
  NAND2_X1 U808 ( .A1(G119), .A2(n879), .ZN(n734) );
  AND2_X1 U809 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U810 ( .A1(n737), .A2(n736), .ZN(n900) );
  NAND2_X1 U811 ( .A1(G1991), .A2(n900), .ZN(n738) );
  NAND2_X1 U812 ( .A1(n739), .A2(n738), .ZN(n976) );
  XNOR2_X1 U813 ( .A(n516), .B(n743), .ZN(n745) );
  XNOR2_X1 U814 ( .A(G1986), .B(G290), .ZN(n1012) );
  NAND2_X1 U815 ( .A1(n1012), .A2(n758), .ZN(n744) );
  NAND2_X1 U816 ( .A1(n745), .A2(n744), .ZN(n761) );
  XOR2_X1 U817 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n753) );
  NOR2_X1 U818 ( .A1(G1991), .A2(n900), .ZN(n972) );
  NOR2_X1 U819 ( .A1(G1986), .A2(G290), .ZN(n746) );
  XOR2_X1 U820 ( .A(n746), .B(KEYINPUT103), .Z(n747) );
  NOR2_X1 U821 ( .A1(n972), .A2(n747), .ZN(n748) );
  XNOR2_X1 U822 ( .A(n748), .B(KEYINPUT104), .ZN(n749) );
  NOR2_X1 U823 ( .A1(n976), .A2(n749), .ZN(n751) );
  NOR2_X1 U824 ( .A1(n893), .A2(G1996), .ZN(n750) );
  XNOR2_X1 U825 ( .A(n750), .B(KEYINPUT102), .ZN(n982) );
  NOR2_X1 U826 ( .A1(n751), .A2(n982), .ZN(n752) );
  XNOR2_X1 U827 ( .A(n753), .B(n752), .ZN(n755) );
  NAND2_X1 U828 ( .A1(n755), .A2(n754), .ZN(n757) );
  NAND2_X1 U829 ( .A1(n756), .A2(n887), .ZN(n973) );
  NAND2_X1 U830 ( .A1(n757), .A2(n973), .ZN(n759) );
  NAND2_X1 U831 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U832 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U833 ( .A(n762), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U834 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U835 ( .A1(G135), .A2(n874), .ZN(n764) );
  NAND2_X1 U836 ( .A1(G111), .A2(n878), .ZN(n763) );
  NAND2_X1 U837 ( .A1(n764), .A2(n763), .ZN(n767) );
  NAND2_X1 U838 ( .A1(n879), .A2(G123), .ZN(n765) );
  XOR2_X1 U839 ( .A(KEYINPUT18), .B(n765), .Z(n766) );
  NOR2_X1 U840 ( .A1(n767), .A2(n766), .ZN(n769) );
  NAND2_X1 U841 ( .A1(n875), .A2(G99), .ZN(n768) );
  NAND2_X1 U842 ( .A1(n769), .A2(n768), .ZN(n969) );
  XNOR2_X1 U843 ( .A(G2096), .B(n969), .ZN(n770) );
  OR2_X1 U844 ( .A1(G2100), .A2(n770), .ZN(G156) );
  INV_X1 U845 ( .A(G132), .ZN(G219) );
  INV_X1 U846 ( .A(G82), .ZN(G220) );
  INV_X1 U847 ( .A(G57), .ZN(G237) );
  NAND2_X1 U848 ( .A1(G7), .A2(G661), .ZN(n771) );
  XNOR2_X1 U849 ( .A(n771), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U850 ( .A(G223), .ZN(n829) );
  NAND2_X1 U851 ( .A1(n829), .A2(G567), .ZN(n772) );
  XNOR2_X1 U852 ( .A(n772), .B(KEYINPUT11), .ZN(n773) );
  XNOR2_X1 U853 ( .A(KEYINPUT71), .B(n773), .ZN(G234) );
  INV_X1 U854 ( .A(G860), .ZN(n780) );
  OR2_X1 U855 ( .A1(n1015), .A2(n780), .ZN(G153) );
  NAND2_X1 U856 ( .A1(G301), .A2(G868), .ZN(n774) );
  XNOR2_X1 U857 ( .A(n774), .B(KEYINPUT74), .ZN(n776) );
  INV_X1 U858 ( .A(G868), .ZN(n810) );
  NAND2_X1 U859 ( .A1(n810), .A2(n781), .ZN(n775) );
  NAND2_X1 U860 ( .A1(n776), .A2(n775), .ZN(G284) );
  INV_X1 U861 ( .A(n1004), .ZN(G299) );
  XNOR2_X1 U862 ( .A(KEYINPUT76), .B(n810), .ZN(n777) );
  NOR2_X1 U863 ( .A1(G286), .A2(n777), .ZN(n779) );
  NOR2_X1 U864 ( .A1(G868), .A2(G299), .ZN(n778) );
  NOR2_X1 U865 ( .A1(n779), .A2(n778), .ZN(G297) );
  NAND2_X1 U866 ( .A1(n780), .A2(G559), .ZN(n782) );
  INV_X1 U867 ( .A(n781), .ZN(n998) );
  NAND2_X1 U868 ( .A1(n782), .A2(n998), .ZN(n783) );
  XNOR2_X1 U869 ( .A(n783), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U870 ( .A1(G868), .A2(n1015), .ZN(n786) );
  NAND2_X1 U871 ( .A1(G868), .A2(n998), .ZN(n784) );
  NOR2_X1 U872 ( .A1(G559), .A2(n784), .ZN(n785) );
  NOR2_X1 U873 ( .A1(n786), .A2(n785), .ZN(G282) );
  NAND2_X1 U874 ( .A1(G93), .A2(n787), .ZN(n789) );
  NAND2_X1 U875 ( .A1(G80), .A2(n601), .ZN(n788) );
  NAND2_X1 U876 ( .A1(n789), .A2(n788), .ZN(n793) );
  NAND2_X1 U877 ( .A1(G67), .A2(n790), .ZN(n791) );
  XNOR2_X1 U878 ( .A(KEYINPUT77), .B(n791), .ZN(n792) );
  NOR2_X1 U879 ( .A1(n793), .A2(n792), .ZN(n796) );
  NAND2_X1 U880 ( .A1(n794), .A2(G55), .ZN(n795) );
  NAND2_X1 U881 ( .A1(n796), .A2(n795), .ZN(n809) );
  NAND2_X1 U882 ( .A1(n998), .A2(G559), .ZN(n807) );
  XNOR2_X1 U883 ( .A(n1015), .B(n807), .ZN(n797) );
  NOR2_X1 U884 ( .A1(G860), .A2(n797), .ZN(n798) );
  XOR2_X1 U885 ( .A(n809), .B(n798), .Z(G145) );
  XNOR2_X1 U886 ( .A(KEYINPUT81), .B(KEYINPUT80), .ZN(n800) );
  XNOR2_X1 U887 ( .A(G288), .B(KEYINPUT19), .ZN(n799) );
  XNOR2_X1 U888 ( .A(n800), .B(n799), .ZN(n801) );
  XNOR2_X1 U889 ( .A(n1004), .B(n801), .ZN(n803) );
  XNOR2_X1 U890 ( .A(G305), .B(G166), .ZN(n802) );
  XNOR2_X1 U891 ( .A(n803), .B(n802), .ZN(n804) );
  XNOR2_X1 U892 ( .A(n804), .B(G290), .ZN(n805) );
  XNOR2_X1 U893 ( .A(n805), .B(n809), .ZN(n806) );
  XNOR2_X1 U894 ( .A(n806), .B(n1015), .ZN(n904) );
  XNOR2_X1 U895 ( .A(n807), .B(n904), .ZN(n808) );
  NAND2_X1 U896 ( .A1(n808), .A2(G868), .ZN(n812) );
  NAND2_X1 U897 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U898 ( .A1(n812), .A2(n811), .ZN(G295) );
  XNOR2_X1 U899 ( .A(KEYINPUT20), .B(KEYINPUT83), .ZN(n815) );
  NAND2_X1 U900 ( .A1(G2078), .A2(G2084), .ZN(n813) );
  XNOR2_X1 U901 ( .A(n813), .B(KEYINPUT82), .ZN(n814) );
  XNOR2_X1 U902 ( .A(n815), .B(n814), .ZN(n816) );
  NAND2_X1 U903 ( .A1(G2090), .A2(n816), .ZN(n817) );
  XNOR2_X1 U904 ( .A(KEYINPUT21), .B(n817), .ZN(n818) );
  NAND2_X1 U905 ( .A1(n818), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U906 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U907 ( .A1(G120), .A2(G108), .ZN(n819) );
  NOR2_X1 U908 ( .A1(G237), .A2(n819), .ZN(n820) );
  NAND2_X1 U909 ( .A1(G69), .A2(n820), .ZN(n835) );
  NAND2_X1 U910 ( .A1(n835), .A2(G567), .ZN(n826) );
  NOR2_X1 U911 ( .A1(G220), .A2(G219), .ZN(n821) );
  XNOR2_X1 U912 ( .A(KEYINPUT22), .B(n821), .ZN(n822) );
  NAND2_X1 U913 ( .A1(n822), .A2(G96), .ZN(n823) );
  NOR2_X1 U914 ( .A1(G218), .A2(n823), .ZN(n824) );
  XOR2_X1 U915 ( .A(KEYINPUT84), .B(n824), .Z(n836) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n836), .ZN(n825) );
  NAND2_X1 U917 ( .A1(n826), .A2(n825), .ZN(n837) );
  NAND2_X1 U918 ( .A1(G483), .A2(G661), .ZN(n827) );
  NOR2_X1 U919 ( .A1(n837), .A2(n827), .ZN(n832) );
  NAND2_X1 U920 ( .A1(n832), .A2(G36), .ZN(n828) );
  XOR2_X1 U921 ( .A(KEYINPUT85), .B(n828), .Z(G176) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n829), .ZN(G217) );
  NAND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n830) );
  XOR2_X1 U924 ( .A(KEYINPUT106), .B(n830), .Z(n831) );
  NAND2_X1 U925 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U927 ( .A1(n833), .A2(n832), .ZN(n834) );
  XOR2_X1 U928 ( .A(KEYINPUT107), .B(n834), .Z(G188) );
  XOR2_X1 U929 ( .A(G96), .B(KEYINPUT108), .Z(G221) );
  XNOR2_X1 U930 ( .A(G108), .B(KEYINPUT119), .ZN(G238) );
  INV_X1 U932 ( .A(G120), .ZN(G236) );
  NOR2_X1 U933 ( .A1(n836), .A2(n835), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  INV_X1 U935 ( .A(n837), .ZN(G319) );
  XOR2_X1 U936 ( .A(G2100), .B(G2096), .Z(n839) );
  XNOR2_X1 U937 ( .A(KEYINPUT42), .B(G2678), .ZN(n838) );
  XNOR2_X1 U938 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U939 ( .A(KEYINPUT43), .B(G2090), .Z(n841) );
  XNOR2_X1 U940 ( .A(G2067), .B(G2072), .ZN(n840) );
  XNOR2_X1 U941 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U942 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U943 ( .A(G2078), .B(G2084), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(G227) );
  XOR2_X1 U945 ( .A(G1956), .B(G1961), .Z(n847) );
  XNOR2_X1 U946 ( .A(G1976), .B(G1971), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U948 ( .A(n848), .B(G2474), .Z(n850) );
  XNOR2_X1 U949 ( .A(G1981), .B(G1966), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U951 ( .A(KEYINPUT41), .B(G1986), .Z(n852) );
  XNOR2_X1 U952 ( .A(G1996), .B(G1991), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n854), .B(n853), .ZN(G229) );
  NAND2_X1 U955 ( .A1(G124), .A2(n879), .ZN(n855) );
  XOR2_X1 U956 ( .A(KEYINPUT109), .B(n855), .Z(n856) );
  XNOR2_X1 U957 ( .A(n856), .B(KEYINPUT44), .ZN(n858) );
  NAND2_X1 U958 ( .A1(G112), .A2(n878), .ZN(n857) );
  NAND2_X1 U959 ( .A1(n858), .A2(n857), .ZN(n862) );
  NAND2_X1 U960 ( .A1(G136), .A2(n874), .ZN(n860) );
  NAND2_X1 U961 ( .A1(G100), .A2(n875), .ZN(n859) );
  NAND2_X1 U962 ( .A1(n860), .A2(n859), .ZN(n861) );
  NOR2_X1 U963 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U964 ( .A(KEYINPUT110), .B(n863), .ZN(G162) );
  NAND2_X1 U965 ( .A1(G118), .A2(n878), .ZN(n873) );
  NAND2_X1 U966 ( .A1(n879), .A2(G130), .ZN(n864) );
  XNOR2_X1 U967 ( .A(KEYINPUT111), .B(n864), .ZN(n871) );
  NAND2_X1 U968 ( .A1(n874), .A2(G142), .ZN(n865) );
  XNOR2_X1 U969 ( .A(n865), .B(KEYINPUT112), .ZN(n867) );
  NAND2_X1 U970 ( .A1(G106), .A2(n875), .ZN(n866) );
  NAND2_X1 U971 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U972 ( .A(KEYINPUT113), .B(n868), .ZN(n869) );
  XNOR2_X1 U973 ( .A(KEYINPUT45), .B(n869), .ZN(n870) );
  NOR2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n872) );
  NAND2_X1 U975 ( .A1(n873), .A2(n872), .ZN(n902) );
  NAND2_X1 U976 ( .A1(G139), .A2(n874), .ZN(n877) );
  NAND2_X1 U977 ( .A1(G103), .A2(n875), .ZN(n876) );
  NAND2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n886) );
  XNOR2_X1 U979 ( .A(KEYINPUT116), .B(KEYINPUT47), .ZN(n884) );
  NAND2_X1 U980 ( .A1(n878), .A2(G115), .ZN(n882) );
  NAND2_X1 U981 ( .A1(n879), .A2(G127), .ZN(n880) );
  XOR2_X1 U982 ( .A(KEYINPUT115), .B(n880), .Z(n881) );
  NAND2_X1 U983 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U984 ( .A(n884), .B(n883), .Z(n885) );
  NOR2_X1 U985 ( .A1(n886), .A2(n885), .ZN(n977) );
  XNOR2_X1 U986 ( .A(G164), .B(n887), .ZN(n888) );
  XNOR2_X1 U987 ( .A(n888), .B(G162), .ZN(n892) );
  XOR2_X1 U988 ( .A(KEYINPUT114), .B(KEYINPUT46), .Z(n890) );
  XNOR2_X1 U989 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n889) );
  XNOR2_X1 U990 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U991 ( .A(n892), .B(n891), .Z(n897) );
  XNOR2_X1 U992 ( .A(G160), .B(n893), .ZN(n894) );
  XNOR2_X1 U993 ( .A(n894), .B(n969), .ZN(n895) );
  XNOR2_X1 U994 ( .A(n895), .B(KEYINPUT48), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U996 ( .A(n977), .B(n898), .Z(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U999 ( .A1(G37), .A2(n903), .ZN(G395) );
  XOR2_X1 U1000 ( .A(n904), .B(G286), .Z(n906) );
  XNOR2_X1 U1001 ( .A(G171), .B(n998), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n907), .ZN(G397) );
  XOR2_X1 U1004 ( .A(G2451), .B(G2430), .Z(n909) );
  XNOR2_X1 U1005 ( .A(G2438), .B(G2443), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n909), .B(n908), .ZN(n915) );
  XOR2_X1 U1007 ( .A(G2435), .B(G2454), .Z(n911) );
  XNOR2_X1 U1008 ( .A(G1348), .B(G1341), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(n913) );
  XOR2_X1 U1010 ( .A(G2446), .B(G2427), .Z(n912) );
  XNOR2_X1 U1011 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1012 ( .A(n915), .B(n914), .Z(n916) );
  NAND2_X1 U1013 ( .A1(G14), .A2(n916), .ZN(n922) );
  NAND2_X1 U1014 ( .A1(G319), .A2(n922), .ZN(n919) );
  NOR2_X1 U1015 ( .A1(G227), .A2(G229), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1017 ( .A1(n919), .A2(n918), .ZN(n921) );
  NOR2_X1 U1018 ( .A1(G395), .A2(G397), .ZN(n920) );
  NAND2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1020 ( .A(G225), .ZN(G308) );
  INV_X1 U1021 ( .A(G69), .ZN(G235) );
  INV_X1 U1022 ( .A(n922), .ZN(G401) );
  XNOR2_X1 U1023 ( .A(G20), .B(n1005), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(G1981), .B(G6), .ZN(n924) );
  XNOR2_X1 U1025 ( .A(G1341), .B(G19), .ZN(n923) );
  NOR2_X1 U1026 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n929) );
  XOR2_X1 U1028 ( .A(KEYINPUT59), .B(G1348), .Z(n927) );
  XNOR2_X1 U1029 ( .A(G4), .B(n927), .ZN(n928) );
  NOR2_X1 U1030 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1031 ( .A(KEYINPUT60), .B(n930), .ZN(n934) );
  XNOR2_X1 U1032 ( .A(G1966), .B(G21), .ZN(n932) );
  XNOR2_X1 U1033 ( .A(G5), .B(G1961), .ZN(n931) );
  NOR2_X1 U1034 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1036 ( .A(KEYINPUT124), .B(n935), .ZN(n943) );
  XOR2_X1 U1037 ( .A(G1986), .B(G24), .Z(n939) );
  XNOR2_X1 U1038 ( .A(G1976), .B(G23), .ZN(n937) );
  XNOR2_X1 U1039 ( .A(G1971), .B(G22), .ZN(n936) );
  NOR2_X1 U1040 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1041 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1042 ( .A(KEYINPUT58), .B(n940), .Z(n941) );
  XNOR2_X1 U1043 ( .A(KEYINPUT125), .B(n941), .ZN(n942) );
  NOR2_X1 U1044 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1045 ( .A(KEYINPUT61), .B(n944), .Z(n945) );
  NOR2_X1 U1046 ( .A1(G16), .A2(n945), .ZN(n946) );
  XOR2_X1 U1047 ( .A(KEYINPUT126), .B(n946), .Z(n997) );
  XOR2_X1 U1048 ( .A(G29), .B(KEYINPUT122), .Z(n967) );
  XOR2_X1 U1049 ( .A(G2084), .B(G34), .Z(n947) );
  XNOR2_X1 U1050 ( .A(KEYINPUT54), .B(n947), .ZN(n963) );
  XNOR2_X1 U1051 ( .A(G2090), .B(G35), .ZN(n961) );
  XNOR2_X1 U1052 ( .A(G1996), .B(G32), .ZN(n949) );
  XNOR2_X1 U1053 ( .A(G33), .B(G2072), .ZN(n948) );
  NOR2_X1 U1054 ( .A1(n949), .A2(n948), .ZN(n955) );
  XOR2_X1 U1055 ( .A(G2067), .B(G26), .Z(n950) );
  NAND2_X1 U1056 ( .A1(n950), .A2(G28), .ZN(n953) );
  XNOR2_X1 U1057 ( .A(G25), .B(G1991), .ZN(n951) );
  XNOR2_X1 U1058 ( .A(KEYINPUT120), .B(n951), .ZN(n952) );
  NOR2_X1 U1059 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1060 ( .A1(n955), .A2(n954), .ZN(n958) );
  XNOR2_X1 U1061 ( .A(G27), .B(n956), .ZN(n957) );
  NOR2_X1 U1062 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1063 ( .A(KEYINPUT53), .B(n959), .ZN(n960) );
  NOR2_X1 U1064 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1065 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1066 ( .A(n964), .B(KEYINPUT121), .ZN(n965) );
  XNOR2_X1 U1067 ( .A(n965), .B(KEYINPUT55), .ZN(n966) );
  NAND2_X1 U1068 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1069 ( .A1(G11), .A2(n968), .ZN(n995) );
  XNOR2_X1 U1070 ( .A(G160), .B(G2084), .ZN(n970) );
  NAND2_X1 U1071 ( .A1(n970), .A2(n969), .ZN(n971) );
  NOR2_X1 U1072 ( .A1(n972), .A2(n971), .ZN(n974) );
  NAND2_X1 U1073 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1074 ( .A1(n976), .A2(n975), .ZN(n987) );
  XOR2_X1 U1075 ( .A(G2072), .B(n977), .Z(n979) );
  XOR2_X1 U1076 ( .A(G164), .B(G2078), .Z(n978) );
  NOR2_X1 U1077 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1078 ( .A(KEYINPUT50), .B(n980), .Z(n985) );
  XOR2_X1 U1079 ( .A(G2090), .B(G162), .Z(n981) );
  NOR2_X1 U1080 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1081 ( .A(KEYINPUT51), .B(n983), .ZN(n984) );
  NOR2_X1 U1082 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1083 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n990) );
  XOR2_X1 U1085 ( .A(KEYINPUT52), .B(n990), .Z(n991) );
  NOR2_X1 U1086 ( .A1(KEYINPUT55), .A2(n991), .ZN(n993) );
  INV_X1 U1087 ( .A(G29), .ZN(n992) );
  NOR2_X1 U1088 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1089 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n1026) );
  XOR2_X1 U1091 ( .A(KEYINPUT56), .B(G16), .Z(n1024) );
  XNOR2_X1 U1092 ( .A(G1348), .B(n998), .ZN(n1000) );
  XNOR2_X1 U1093 ( .A(G171), .B(G1961), .ZN(n999) );
  NAND2_X1 U1094 ( .A1(n1000), .A2(n999), .ZN(n1021) );
  XNOR2_X1 U1095 ( .A(G1966), .B(G168), .ZN(n1002) );
  NAND2_X1 U1096 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1097 ( .A(n1003), .B(KEYINPUT57), .ZN(n1019) );
  XNOR2_X1 U1098 ( .A(n1005), .B(n1004), .ZN(n1008) );
  INV_X1 U1099 ( .A(G1971), .ZN(n1006) );
  NOR2_X1 U1100 ( .A1(n1006), .A2(G166), .ZN(n1007) );
  NOR2_X1 U1101 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(G1341), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1109 ( .A(KEYINPUT123), .B(n1022), .Z(n1023) );
  NOR2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1112 ( .A(n1027), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

