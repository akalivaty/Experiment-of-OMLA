//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 0 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961;
  INV_X1    g000(.A(KEYINPUT3), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  NOR3_X1   g002(.A1(new_n188), .A2(KEYINPUT80), .A3(G107), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n187), .B1(new_n189), .B2(KEYINPUT79), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT79), .A3(G104), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n188), .A2(G107), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT81), .B(G101), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT80), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(new_n191), .A3(G104), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT79), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(new_n199), .A3(KEYINPUT3), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n190), .A2(new_n195), .A3(new_n196), .A4(new_n200), .ZN(new_n201));
  AND3_X1   g015(.A1(new_n198), .A2(new_n199), .A3(KEYINPUT3), .ZN(new_n202));
  AOI21_X1  g016(.A(KEYINPUT3), .B1(new_n198), .B2(new_n199), .ZN(new_n203));
  NOR3_X1   g017(.A1(new_n202), .A2(new_n203), .A3(new_n194), .ZN(new_n204));
  INV_X1    g018(.A(G101), .ZN(new_n205));
  OAI211_X1 g019(.A(KEYINPUT4), .B(new_n201), .C1(new_n204), .C2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT2), .ZN(new_n207));
  INV_X1    g021(.A(G113), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT67), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT67), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n210), .B1(KEYINPUT2), .B2(G113), .ZN(new_n211));
  AOI22_X1  g025(.A1(new_n209), .A2(new_n211), .B1(KEYINPUT2), .B2(G113), .ZN(new_n212));
  XNOR2_X1  g026(.A(G116), .B(G119), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G119), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G116), .ZN(new_n216));
  INV_X1    g030(.A(G116), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G119), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT69), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT69), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n213), .A2(new_n221), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n220), .B(new_n222), .C1(new_n212), .C2(KEYINPUT68), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n209), .A2(new_n211), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT2), .A2(G113), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n224), .A2(KEYINPUT68), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n214), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n190), .A2(new_n195), .A3(new_n200), .ZN(new_n228));
  XOR2_X1   g042(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(G101), .A3(new_n229), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n206), .A2(KEYINPUT85), .A3(new_n227), .A4(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT5), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n232), .B1(new_n220), .B2(new_n222), .ZN(new_n233));
  OAI21_X1  g047(.A(G113), .B1(new_n216), .B2(KEYINPUT5), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n214), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n193), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n188), .A2(G107), .ZN(new_n237));
  OAI21_X1  g051(.A(G101), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n201), .A2(new_n238), .ZN(new_n239));
  OR2_X1    g053(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n231), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n224), .A2(new_n225), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n212), .A2(KEYINPUT68), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n244), .A2(new_n245), .A3(new_n220), .A4(new_n222), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n198), .A2(new_n199), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n194), .B1(new_n247), .B2(new_n187), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n205), .B1(new_n248), .B2(new_n200), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n246), .A2(new_n214), .B1(new_n249), .B2(new_n229), .ZN(new_n250));
  AOI21_X1  g064(.A(KEYINPUT85), .B1(new_n250), .B2(new_n206), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT86), .B1(new_n241), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT85), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n227), .A2(new_n230), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n201), .A2(KEYINPUT4), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(new_n249), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n253), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT86), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n257), .A2(new_n258), .A3(new_n231), .A4(new_n240), .ZN(new_n259));
  XNOR2_X1  g073(.A(G110), .B(G122), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n252), .A2(KEYINPUT6), .A3(new_n259), .A4(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n257), .A2(new_n231), .A3(new_n240), .A4(new_n260), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT87), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n231), .A2(new_n240), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT87), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n266), .A2(new_n267), .A3(new_n257), .A4(new_n260), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n263), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n252), .A2(new_n259), .A3(new_n261), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n262), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT1), .ZN(new_n272));
  INV_X1    g086(.A(G146), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n272), .B1(G143), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G128), .ZN(new_n275));
  INV_X1    g089(.A(G143), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(G146), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n273), .A2(G143), .ZN(new_n278));
  OAI22_X1  g092(.A1(new_n274), .A2(new_n275), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n273), .A2(G143), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n276), .A2(G146), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n280), .A2(new_n281), .A3(new_n272), .A4(G128), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(G125), .ZN(new_n284));
  OR2_X1    g098(.A1(new_n284), .A2(KEYINPUT88), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(KEYINPUT88), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT0), .A4(G128), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n277), .A2(new_n278), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT0), .B(G128), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(G125), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G953), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G224), .ZN(new_n295));
  XOR2_X1   g109(.A(new_n293), .B(new_n295), .Z(new_n296));
  NAND2_X1  g110(.A1(new_n271), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n265), .A2(new_n268), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n235), .B1(new_n201), .B2(new_n238), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n260), .B(KEYINPUT8), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT89), .B1(new_n213), .B2(KEYINPUT5), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n301), .A2(new_n234), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n213), .A2(KEYINPUT89), .A3(KEYINPUT5), .ZN(new_n303));
  AOI22_X1  g117(.A1(new_n302), .A2(new_n303), .B1(new_n212), .B2(new_n213), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n300), .B1(new_n304), .B2(new_n239), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n299), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT90), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n287), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n285), .A2(KEYINPUT90), .A3(new_n286), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n295), .A2(KEYINPUT7), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n308), .A2(new_n292), .A3(new_n309), .A4(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n293), .A2(KEYINPUT7), .A3(new_n295), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n306), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n298), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G902), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n297), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(G210), .B1(G237), .B2(G902), .ZN(new_n319));
  XOR2_X1   g133(.A(new_n319), .B(KEYINPUT91), .Z(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n297), .A2(new_n317), .A3(new_n319), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(G214), .B1(G237), .B2(G902), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n324), .B(KEYINPUT84), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT9), .B(G234), .ZN(new_n328));
  INV_X1    g142(.A(G217), .ZN(new_n329));
  NOR3_X1   g143(.A1(new_n328), .A2(new_n329), .A3(G953), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT96), .ZN(new_n331));
  INV_X1    g145(.A(G122), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n331), .B1(new_n332), .B2(G116), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n217), .A2(KEYINPUT96), .A3(G122), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n335), .A2(KEYINPUT14), .B1(G116), .B2(new_n332), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(KEYINPUT14), .B2(new_n335), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G107), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n332), .A2(G116), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n335), .A2(new_n191), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n276), .A2(G128), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n275), .A2(G143), .ZN(new_n342));
  INV_X1    g156(.A(G134), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n341), .A2(new_n342), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G134), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n340), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n338), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT13), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n341), .A2(KEYINPUT97), .A3(new_n349), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n350), .B(new_n342), .C1(new_n349), .C2(new_n341), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT97), .B1(new_n341), .B2(new_n349), .ZN(new_n352));
  OAI21_X1  g166(.A(G134), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n191), .B1(new_n335), .B2(new_n339), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n353), .B(new_n344), .C1(new_n354), .C2(new_n340), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n330), .B1(new_n348), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n348), .A2(new_n355), .A3(new_n330), .ZN(new_n358));
  AOI21_X1  g172(.A(G902), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT98), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n358), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n315), .B1(new_n362), .B2(new_n356), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT98), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT15), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n361), .A2(new_n364), .B1(new_n365), .B2(G478), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n363), .A2(KEYINPUT98), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(G478), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT99), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n359), .A2(new_n360), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n368), .B1(new_n371), .B2(new_n367), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT99), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n361), .A2(new_n365), .A3(G478), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n294), .A2(G952), .ZN(new_n377));
  NAND2_X1  g191(.A1(G234), .A2(G237), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT21), .B(G898), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n378), .A2(G902), .A3(G953), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n379), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT92), .ZN(new_n384));
  INV_X1    g198(.A(G237), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(new_n294), .A3(G214), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(new_n276), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n384), .B1(new_n387), .B2(G131), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n386), .B(G143), .ZN(new_n389));
  INV_X1    g203(.A(G131), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(KEYINPUT92), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n387), .A2(G131), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n388), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  OR2_X1    g207(.A1(new_n393), .A2(KEYINPUT17), .ZN(new_n394));
  XNOR2_X1  g208(.A(G125), .B(G140), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT16), .ZN(new_n396));
  INV_X1    g210(.A(G125), .ZN(new_n397));
  OR3_X1    g211(.A1(new_n397), .A2(KEYINPUT16), .A3(G140), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n273), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n396), .A2(G146), .A3(new_n398), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n387), .A2(KEYINPUT17), .A3(G131), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT94), .ZN(new_n404));
  OR2_X1    g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n404), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n402), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n394), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT18), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n389), .B1(new_n409), .B2(new_n390), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n387), .A2(KEYINPUT18), .A3(G131), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n395), .B(new_n273), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(G113), .B(G122), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n415), .B(new_n188), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT20), .ZN(new_n418));
  INV_X1    g232(.A(new_n413), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n419), .A2(new_n416), .ZN(new_n420));
  NOR2_X1   g234(.A1(KEYINPUT93), .A2(KEYINPUT19), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n395), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(KEYINPUT93), .A2(KEYINPUT19), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n422), .B(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n273), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(new_n393), .A3(new_n401), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(G475), .A2(G902), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n417), .A2(new_n418), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n419), .B1(new_n394), .B2(new_n407), .ZN(new_n430));
  INV_X1    g244(.A(new_n416), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n427), .B(new_n428), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT20), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n416), .A2(KEYINPUT95), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n315), .B1(new_n414), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n430), .A2(new_n435), .ZN(new_n438));
  OAI21_X1  g252(.A(G475), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n376), .A2(new_n383), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n291), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n443), .B(new_n230), .C1(new_n255), .C2(new_n249), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n201), .A2(new_n283), .A3(new_n238), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT10), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n201), .A2(new_n283), .A3(KEYINPUT10), .A4(new_n238), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n444), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT11), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n450), .B1(new_n343), .B2(G137), .ZN(new_n451));
  INV_X1    g265(.A(G137), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(KEYINPUT11), .A3(G134), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n343), .A2(G137), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(KEYINPUT64), .A2(G131), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n451), .A2(new_n453), .A3(new_n456), .A4(new_n454), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n449), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n460), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n444), .A2(new_n462), .A3(new_n447), .A4(new_n448), .ZN(new_n463));
  XNOR2_X1  g277(.A(G110), .B(G140), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n294), .A2(G227), .ZN(new_n465));
  XOR2_X1   g279(.A(new_n464), .B(new_n465), .Z(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n461), .A2(new_n463), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n463), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n283), .B1(new_n201), .B2(new_n238), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n470), .B1(KEYINPUT83), .B2(new_n445), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT83), .ZN(new_n472));
  AOI211_X1 g286(.A(new_n472), .B(new_n283), .C1(new_n201), .C2(new_n238), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n460), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT12), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g290(.A(KEYINPUT12), .B(new_n460), .C1(new_n471), .C2(new_n473), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n469), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n466), .B(KEYINPUT78), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n468), .B(G469), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G469), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n463), .A2(new_n467), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n482), .B1(new_n476), .B2(new_n477), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n467), .B1(new_n461), .B2(new_n463), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n481), .B(new_n315), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n481), .A2(new_n315), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n480), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(G221), .B1(new_n328), .B2(G902), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(KEYINPUT77), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NOR3_X1   g306(.A1(new_n327), .A2(new_n442), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT23), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n494), .A2(new_n215), .A3(G128), .ZN(new_n495));
  AOI21_X1  g309(.A(KEYINPUT23), .B1(new_n275), .B2(G119), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n275), .A2(G119), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G110), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(G119), .B(G128), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(KEYINPUT75), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT24), .B(G110), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n500), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  OR2_X1    g319(.A1(new_n505), .A2(KEYINPUT76), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(KEYINPUT76), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n395), .A2(new_n273), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n506), .A2(new_n507), .A3(new_n401), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n502), .A2(new_n504), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n402), .B(new_n510), .C1(new_n499), .C2(new_n498), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT22), .B(G137), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n294), .A2(G221), .A3(G234), .ZN(new_n514));
  XOR2_X1   g328(.A(new_n513), .B(new_n514), .Z(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n509), .A2(new_n511), .A3(new_n515), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(new_n315), .A3(new_n518), .ZN(new_n519));
  XOR2_X1   g333(.A(new_n519), .B(KEYINPUT25), .Z(new_n520));
  AOI21_X1  g334(.A(new_n329), .B1(G234), .B2(new_n315), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n517), .A2(new_n518), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n521), .A2(G902), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  XOR2_X1   g340(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n527));
  NAND3_X1  g341(.A1(new_n385), .A2(new_n294), .A3(G210), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT26), .B(G101), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n529), .B(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT65), .ZN(new_n532));
  XNOR2_X1  g346(.A(G134), .B(G137), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n532), .B1(new_n533), .B2(new_n390), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n343), .A2(G137), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n452), .A2(G134), .ZN(new_n536));
  OAI211_X1 g350(.A(KEYINPUT65), .B(G131), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n451), .A2(new_n453), .A3(new_n390), .A4(new_n454), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n283), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT66), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n443), .A2(new_n460), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n538), .A2(new_n283), .A3(new_n539), .A4(KEYINPUT66), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n227), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT73), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n543), .A2(new_n540), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n550), .A2(new_n227), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n552), .B1(new_n546), .B2(new_n547), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT28), .B1(new_n549), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n551), .A2(KEYINPUT28), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n531), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n543), .A2(new_n540), .A3(KEYINPUT30), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT70), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n543), .A2(new_n540), .A3(KEYINPUT70), .A4(KEYINPUT30), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT30), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n560), .A2(new_n561), .B1(new_n545), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n551), .B1(new_n563), .B2(new_n227), .ZN(new_n564));
  AOI21_X1  g378(.A(KEYINPUT72), .B1(new_n564), .B2(new_n531), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n560), .A2(new_n561), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n545), .A2(new_n562), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(new_n567), .A3(new_n227), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n568), .A2(KEYINPUT72), .A3(new_n552), .A4(new_n531), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT31), .B1(new_n565), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n568), .A2(new_n552), .A3(new_n531), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT31), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n557), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(G472), .A2(G902), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT74), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT32), .ZN(new_n579));
  INV_X1    g393(.A(new_n531), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT28), .ZN(new_n581));
  INV_X1    g395(.A(new_n553), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n581), .B1(new_n582), .B2(new_n548), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n580), .B1(new_n583), .B2(new_n555), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT72), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n572), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n573), .B1(new_n586), .B2(new_n569), .ZN(new_n587));
  INV_X1    g401(.A(new_n574), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n584), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT74), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(new_n590), .A3(new_n576), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n578), .A2(new_n579), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n550), .B(new_n227), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n555), .B1(new_n593), .B2(KEYINPUT28), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT29), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n580), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(G902), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n583), .A2(new_n555), .A3(new_n580), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n568), .A2(new_n552), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n580), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n595), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n597), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G472), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n589), .A2(KEYINPUT32), .A3(new_n576), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n526), .B1(new_n592), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n493), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(new_n607), .B(new_n196), .Z(G3));
  OAI21_X1  g422(.A(G472), .B1(new_n575), .B2(G902), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n578), .A2(new_n609), .A3(new_n591), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n610), .A2(new_n526), .A3(new_n492), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n297), .A2(new_n319), .A3(new_n317), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n319), .B1(new_n297), .B2(new_n317), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n326), .B(new_n383), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  OR2_X1    g428(.A1(new_n362), .A2(KEYINPUT101), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n362), .A2(KEYINPUT101), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n615), .A2(KEYINPUT33), .A3(new_n357), .A4(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT100), .B(KEYINPUT33), .Z(new_n618));
  OAI21_X1  g432(.A(new_n618), .B1(new_n362), .B2(new_n356), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n315), .A2(G478), .ZN(new_n621));
  OAI22_X1  g435(.A1(new_n620), .A2(new_n621), .B1(G478), .B2(new_n359), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n440), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n614), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n611), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT34), .B(G104), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G6));
  INV_X1    g441(.A(new_n376), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n441), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n614), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n611), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT35), .B(G107), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  NOR2_X1   g447(.A1(new_n516), .A2(KEYINPUT36), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT102), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n512), .B(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n524), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n522), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n610), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n493), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT37), .B(G110), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G12));
  AOI21_X1  g458(.A(new_n316), .B1(new_n296), .B2(new_n271), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(new_n319), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n646), .A2(new_n326), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n592), .A2(new_n605), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n492), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n639), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(new_n379), .B(KEYINPUT103), .Z(new_n652));
  OAI21_X1  g466(.A(new_n652), .B1(G900), .B2(new_n382), .ZN(new_n653));
  XOR2_X1   g467(.A(new_n653), .B(KEYINPUT104), .Z(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n628), .A2(new_n441), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n649), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT105), .B(G128), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G30));
  XOR2_X1   g474(.A(new_n654), .B(KEYINPUT39), .Z(new_n661));
  NAND2_X1  g475(.A1(new_n650), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT107), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT40), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n323), .B(new_n666), .Z(new_n667));
  NOR2_X1   g481(.A1(new_n565), .A2(new_n570), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n593), .A2(new_n580), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g484(.A(G472), .B1(new_n670), .B2(G902), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n671), .A2(new_n604), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n592), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n325), .B1(new_n434), .B2(new_n439), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n674), .A2(new_n370), .A3(new_n375), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n640), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n665), .A2(new_n667), .A3(new_n673), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT108), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G143), .ZN(G45));
  NAND3_X1  g493(.A1(new_n622), .A2(new_n440), .A3(new_n655), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n651), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n649), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G146), .ZN(G48));
  OAI21_X1  g497(.A(new_n315), .B1(new_n483), .B2(new_n484), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(G469), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n489), .A3(new_n485), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n685), .A2(KEYINPUT109), .A3(new_n489), .A4(new_n485), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n606), .A2(new_n624), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT41), .B(G113), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G15));
  NAND3_X1  g507(.A1(new_n606), .A2(new_n630), .A3(new_n690), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G116), .ZN(G18));
  AOI21_X1  g509(.A(new_n442), .B1(new_n592), .B2(new_n605), .ZN(new_n696));
  INV_X1    g510(.A(new_n686), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n326), .B(new_n697), .C1(new_n612), .C2(new_n613), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n640), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G119), .ZN(G21));
  NAND2_X1  g515(.A1(new_n571), .A2(new_n574), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n594), .A2(new_n531), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n577), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n609), .A2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(G472), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n589), .B2(new_n315), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT110), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n705), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n675), .B1(new_n612), .B2(new_n613), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n688), .A2(new_n383), .A3(new_n689), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n526), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n711), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G122), .ZN(G24));
  INV_X1    g531(.A(new_n680), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n699), .A2(new_n711), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  OAI21_X1  g534(.A(new_n579), .B1(new_n575), .B2(new_n577), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n526), .B1(new_n605), .B2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n320), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n322), .B(new_n326), .C1(new_n723), .C2(new_n645), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n488), .A2(new_n489), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n488), .A2(KEYINPUT111), .A3(new_n489), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n724), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n722), .A2(KEYINPUT42), .A3(new_n718), .A4(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n648), .A2(new_n730), .A3(new_n715), .A4(new_n718), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT42), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n733), .B1(new_n732), .B2(new_n734), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n731), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G131), .ZN(G33));
  INV_X1    g552(.A(new_n606), .ZN(new_n739));
  INV_X1    g553(.A(new_n730), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n739), .A2(new_n656), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(new_n343), .ZN(G36));
  INV_X1    g556(.A(new_n489), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n468), .B1(new_n478), .B2(new_n479), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT45), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n744), .A2(new_n745), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n746), .A2(new_n747), .A3(new_n481), .ZN(new_n748));
  OR2_X1    g562(.A1(new_n748), .A2(new_n486), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT46), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n485), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n752), .B1(new_n749), .B2(new_n750), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n743), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n754), .A2(new_n661), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n441), .A2(new_n622), .ZN(new_n756));
  XOR2_X1   g570(.A(new_n756), .B(KEYINPUT43), .Z(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(new_n610), .A3(new_n639), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n724), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n755), .B(new_n760), .C1(new_n759), .C2(new_n758), .ZN(new_n761));
  XOR2_X1   g575(.A(KEYINPUT113), .B(G137), .Z(new_n762));
  XNOR2_X1  g576(.A(new_n761), .B(new_n762), .ZN(G39));
  XNOR2_X1  g577(.A(new_n754), .B(KEYINPUT47), .ZN(new_n764));
  INV_X1    g578(.A(new_n648), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n715), .A2(new_n724), .A3(new_n680), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G140), .ZN(G42));
  NAND2_X1  g582(.A1(new_n732), .A2(new_n734), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(KEYINPUT112), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n741), .B1(new_n772), .B2(new_n731), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n366), .A2(new_n369), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n623), .B1(new_n774), .B2(new_n440), .ZN(new_n775));
  AND4_X1   g589(.A1(new_n326), .A2(new_n323), .A3(new_n383), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n611), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n642), .A2(new_n607), .A3(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n691), .A2(new_n694), .A3(new_n700), .A4(new_n716), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n705), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n709), .A2(KEYINPUT110), .ZN(new_n783));
  AOI211_X1 g597(.A(new_n706), .B(new_n708), .C1(new_n589), .C2(new_n315), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n715), .B(new_n782), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  AOI22_X1  g600(.A1(new_n786), .A2(new_n714), .B1(new_n699), .B2(new_n696), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(KEYINPUT114), .A3(new_n691), .A4(new_n694), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n778), .B1(new_n781), .B2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT115), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n711), .A2(new_n639), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n730), .A2(new_n718), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n441), .A2(new_n774), .A3(new_n655), .ZN(new_n793));
  OR3_X1    g607(.A1(new_n651), .A2(new_n724), .A3(new_n793), .ZN(new_n794));
  OAI22_X1  g608(.A1(new_n791), .A2(new_n792), .B1(new_n794), .B2(new_n765), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n773), .A2(new_n789), .A3(new_n790), .A4(new_n796), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n647), .B(new_n648), .C1(new_n657), .C2(new_n681), .ZN(new_n798));
  INV_X1    g612(.A(new_n712), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n639), .A2(new_n654), .A3(new_n725), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n673), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n798), .A2(new_n719), .A3(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n798), .A2(KEYINPUT52), .A3(new_n719), .A4(new_n801), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n797), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n781), .A2(new_n788), .ZN(new_n809));
  INV_X1    g623(.A(new_n778), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n741), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n737), .A2(new_n812), .A3(new_n796), .ZN(new_n813));
  OAI21_X1  g627(.A(KEYINPUT115), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n807), .A2(new_n808), .A3(KEYINPUT53), .A4(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n814), .A2(KEYINPUT53), .A3(new_n797), .A4(new_n806), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT116), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n814), .A2(new_n797), .A3(new_n806), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n815), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT54), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n779), .B(new_n825), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n778), .A2(new_n795), .A3(new_n819), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n826), .A2(new_n806), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n773), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n824), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n806), .A2(new_n827), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(KEYINPUT118), .A3(new_n773), .A4(new_n826), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n820), .A2(new_n823), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n757), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n836), .A2(new_n652), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n724), .A2(new_n686), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n837), .A2(new_n722), .A3(new_n838), .ZN(new_n839));
  XOR2_X1   g653(.A(new_n839), .B(KEYINPUT48), .Z(new_n840));
  NOR3_X1   g654(.A1(new_n673), .A2(new_n526), .A3(new_n379), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n838), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n837), .A2(new_n786), .ZN(new_n843));
  OAI221_X1 g657(.A(new_n377), .B1(new_n842), .B2(new_n623), .C1(new_n843), .C2(new_n698), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  NOR4_X1   g659(.A1(new_n843), .A2(new_n667), .A3(new_n326), .A4(new_n686), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT50), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n837), .A2(new_n838), .ZN(new_n848));
  OR2_X1    g662(.A1(new_n622), .A2(new_n440), .ZN(new_n849));
  OAI22_X1  g663(.A1(new_n848), .A2(new_n791), .B1(new_n842), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n685), .A2(new_n485), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n851), .A2(new_n491), .ZN(new_n852));
  OR2_X1    g666(.A1(new_n764), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n843), .A2(new_n724), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n850), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n847), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT51), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n845), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(new_n857), .B2(new_n856), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n822), .A2(new_n835), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n860), .B1(G952), .B2(G953), .ZN(new_n861));
  NOR4_X1   g675(.A1(new_n526), .A2(new_n756), .A3(new_n325), .A4(new_n490), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n851), .A2(KEYINPUT49), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n851), .A2(KEYINPUT49), .ZN(new_n865));
  OR4_X1    g679(.A1(new_n667), .A2(new_n864), .A3(new_n673), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n861), .A2(new_n866), .ZN(G75));
  NOR2_X1   g681(.A1(new_n294), .A2(G952), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n315), .B1(new_n820), .B2(new_n833), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT56), .B1(new_n870), .B2(G210), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n271), .B(new_n296), .Z(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT55), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n869), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n820), .A2(new_n833), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n875), .A2(new_n876), .A3(G902), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n818), .A2(new_n819), .B1(new_n830), .B2(new_n832), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT119), .B1(new_n878), .B2(new_n315), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n877), .A2(new_n879), .A3(new_n320), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT56), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n873), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n874), .B1(new_n880), .B2(new_n882), .ZN(G51));
  XNOR2_X1  g697(.A(new_n486), .B(KEYINPUT57), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n823), .B1(new_n820), .B2(new_n833), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n884), .B1(new_n834), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n886), .B1(new_n484), .B2(new_n483), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n877), .A2(new_n879), .A3(new_n748), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n868), .B1(new_n887), .B2(new_n888), .ZN(G54));
  AND2_X1   g703(.A1(KEYINPUT58), .A2(G475), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n877), .A2(new_n879), .A3(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n417), .A2(new_n427), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n877), .A2(new_n879), .A3(new_n892), .A4(new_n890), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n869), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n894), .A2(new_n896), .ZN(G60));
  INV_X1    g711(.A(new_n620), .ZN(new_n898));
  NAND2_X1  g712(.A1(G478), .A2(G902), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT59), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n898), .B(new_n900), .C1(new_n834), .C2(new_n885), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n869), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n822), .A2(new_n835), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n900), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n902), .B1(new_n904), .B2(new_n620), .ZN(G63));
  NAND2_X1  g719(.A1(G217), .A2(G902), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT120), .Z(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT60), .Z(new_n908));
  NAND3_X1  g722(.A1(new_n875), .A2(new_n637), .A3(new_n908), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n523), .B(KEYINPUT121), .ZN(new_n910));
  INV_X1    g724(.A(new_n908), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n910), .B1(new_n878), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n909), .A2(new_n912), .A3(new_n869), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n913), .B(new_n914), .ZN(G66));
  NAND2_X1  g729(.A1(new_n811), .A2(new_n294), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT122), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n294), .B1(new_n381), .B2(G224), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI221_X1 g733(.A(new_n262), .B1(G898), .B2(new_n294), .C1(new_n269), .C2(new_n270), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n919), .B(new_n920), .Z(G69));
  XNOR2_X1  g735(.A(new_n563), .B(new_n424), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT123), .Z(new_n923));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT108), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n677), .B(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n798), .A2(new_n719), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n927), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n678), .A2(KEYINPUT62), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n767), .A2(new_n761), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n775), .A2(new_n321), .A3(new_n326), .A4(new_n322), .ZN(new_n933));
  OR3_X1    g747(.A1(new_n739), .A2(new_n933), .A3(new_n663), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n923), .B1(new_n936), .B2(G953), .ZN(new_n937));
  NAND2_X1  g751(.A1(G900), .A2(G953), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n755), .A2(new_n799), .A3(new_n722), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n932), .A2(new_n773), .A3(new_n929), .A4(new_n939), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n938), .B(new_n922), .C1(new_n940), .C2(G953), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n294), .B1(G227), .B2(G900), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(G72));
  XNOR2_X1  g758(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n708), .A2(new_n315), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n945), .B(new_n946), .Z(new_n947));
  OAI21_X1  g761(.A(new_n947), .B1(new_n940), .B2(new_n811), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n599), .B(KEYINPUT126), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n580), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT127), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n868), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n931), .A2(new_n789), .A3(new_n935), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT125), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n953), .A2(new_n954), .A3(new_n947), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n949), .A2(new_n580), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n954), .B1(new_n953), .B2(new_n947), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n952), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n947), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n668), .B2(new_n600), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n959), .B1(new_n821), .B2(new_n961), .ZN(G57));
endmodule


