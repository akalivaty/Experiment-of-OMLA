

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764;

  AND2_X1 U372 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U373 ( .A(n482), .B(G119), .ZN(n484) );
  XNOR2_X1 U374 ( .A(G116), .B(G113), .ZN(n483) );
  INV_X1 U375 ( .A(KEYINPUT3), .ZN(n482) );
  XNOR2_X2 U376 ( .A(n453), .B(n373), .ZN(n525) );
  NOR2_X1 U377 ( .A1(G953), .A2(G237), .ZN(n500) );
  NAND2_X2 U378 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X2 U379 ( .A(n525), .B(n546), .ZN(n745) );
  XOR2_X2 U380 ( .A(n545), .B(n493), .Z(n752) );
  INV_X2 U381 ( .A(G953), .ZN(n746) );
  INV_X1 U382 ( .A(G146), .ZN(n479) );
  INV_X1 U383 ( .A(G125), .ZN(n380) );
  XNOR2_X1 U384 ( .A(n562), .B(n491), .ZN(n627) );
  XNOR2_X1 U385 ( .A(n479), .B(n380), .ZN(n379) );
  XNOR2_X1 U386 ( .A(n520), .B(KEYINPUT104), .ZN(n590) );
  NAND2_X1 U387 ( .A1(n519), .A2(n688), .ZN(n520) );
  XNOR2_X1 U388 ( .A(n425), .B(n563), .ZN(n582) );
  NOR2_X1 U389 ( .A1(n603), .A2(n601), .ZN(n702) );
  XNOR2_X1 U390 ( .A(n592), .B(n578), .ZN(n437) );
  XNOR2_X1 U391 ( .A(n409), .B(n408), .ZN(n737) );
  XNOR2_X1 U392 ( .A(n379), .B(KEYINPUT10), .ZN(n493) );
  NOR2_X1 U393 ( .A1(n451), .A2(n445), .ZN(n671) );
  OR2_X2 U394 ( .A1(n663), .A2(G902), .ZN(n490) );
  XNOR2_X2 U395 ( .A(n515), .B(n366), .ZN(n751) );
  XNOR2_X1 U396 ( .A(n586), .B(n357), .ZN(n419) );
  INV_X1 U397 ( .A(KEYINPUT6), .ZN(n491) );
  NOR2_X1 U398 ( .A1(n658), .A2(n534), .ZN(n539) );
  XNOR2_X1 U399 ( .A(n506), .B(n505), .ZN(n576) );
  XNOR2_X1 U400 ( .A(n504), .B(G475), .ZN(n505) );
  XNOR2_X1 U401 ( .A(n365), .B(n524), .ZN(n546) );
  XOR2_X1 U402 ( .A(KEYINPUT74), .B(G107), .Z(n524) );
  XNOR2_X1 U403 ( .A(n523), .B(G110), .ZN(n365) );
  INV_X1 U404 ( .A(KEYINPUT0), .ZN(n376) );
  INV_X1 U405 ( .A(KEYINPUT121), .ZN(n401) );
  INV_X1 U406 ( .A(n690), .ZN(n381) );
  AND2_X1 U407 ( .A1(n418), .A2(n595), .ZN(n417) );
  NOR2_X1 U408 ( .A1(n671), .A2(n559), .ZN(n572) );
  XNOR2_X1 U409 ( .A(n467), .B(n466), .ZN(n560) );
  XNOR2_X1 U410 ( .A(n465), .B(KEYINPUT25), .ZN(n466) );
  NOR2_X1 U411 ( .A1(n737), .A2(G902), .ZN(n467) );
  XNOR2_X1 U412 ( .A(n396), .B(n395), .ZN(n510) );
  INV_X1 U413 ( .A(KEYINPUT8), .ZN(n395) );
  NAND2_X1 U414 ( .A1(n746), .A2(G234), .ZN(n396) );
  XNOR2_X1 U415 ( .A(n478), .B(n530), .ZN(n366) );
  XNOR2_X1 U416 ( .A(KEYINPUT67), .B(G137), .ZN(n478) );
  NOR2_X1 U417 ( .A1(n415), .A2(n414), .ZN(n413) );
  XNOR2_X1 U418 ( .A(n367), .B(KEYINPUT33), .ZN(n374) );
  AND2_X1 U419 ( .A1(n703), .A2(n702), .ZN(n633) );
  BUF_X1 U420 ( .A(n627), .Z(n388) );
  XNOR2_X1 U421 ( .A(n480), .B(n444), .ZN(n443) );
  INV_X1 U422 ( .A(KEYINPUT73), .ZN(n444) );
  XNOR2_X1 U423 ( .A(G137), .B(KEYINPUT23), .ZN(n459) );
  XNOR2_X1 U424 ( .A(n462), .B(n458), .ZN(n410) );
  XNOR2_X1 U425 ( .A(KEYINPUT92), .B(KEYINPUT83), .ZN(n458) );
  XNOR2_X1 U426 ( .A(G110), .B(G119), .ZN(n456) );
  XNOR2_X1 U427 ( .A(n751), .B(G146), .ZN(n363) );
  XNOR2_X1 U428 ( .A(n387), .B(n527), .ZN(n532) );
  XNOR2_X1 U429 ( .A(n580), .B(n579), .ZN(n711) );
  NAND2_X1 U430 ( .A1(n448), .A2(KEYINPUT36), .ZN(n447) );
  INV_X1 U431 ( .A(n542), .ZN(n448) );
  AND2_X1 U432 ( .A1(n542), .A2(n543), .ZN(n450) );
  AND2_X1 U433 ( .A1(n577), .A2(n351), .ZN(n424) );
  INV_X1 U434 ( .A(KEYINPUT22), .ZN(n436) );
  AND2_X1 U435 ( .A1(n402), .A2(n399), .ZN(n398) );
  AND2_X1 U436 ( .A1(n400), .A2(n746), .ZN(n399) );
  NAND2_X1 U437 ( .A1(n735), .A2(n401), .ZN(n400) );
  NAND2_X1 U438 ( .A1(n669), .A2(n668), .ZN(n622) );
  INV_X1 U439 ( .A(G237), .ZN(n535) );
  XOR2_X1 U440 ( .A(G140), .B(G128), .Z(n457) );
  XNOR2_X1 U441 ( .A(G113), .B(G143), .ZN(n494) );
  XOR2_X1 U442 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n495) );
  XNOR2_X1 U443 ( .A(G104), .B(G122), .ZN(n497) );
  XNOR2_X1 U444 ( .A(n379), .B(n350), .ZN(n387) );
  OR2_X1 U445 ( .A1(G953), .A2(G952), .ZN(n475) );
  INV_X1 U446 ( .A(G122), .ZN(n521) );
  NAND2_X1 U447 ( .A1(n349), .A2(n534), .ZN(n428) );
  INV_X1 U448 ( .A(KEYINPUT84), .ZN(n427) );
  XNOR2_X1 U449 ( .A(G107), .B(G116), .ZN(n508) );
  NAND2_X1 U450 ( .A1(n711), .A2(n374), .ZN(n731) );
  XNOR2_X1 U451 ( .A(n411), .B(n583), .ZN(n594) );
  INV_X1 U452 ( .A(n637), .ZN(n412) );
  INV_X1 U453 ( .A(KEYINPUT19), .ZN(n377) );
  INV_X1 U454 ( .A(n388), .ZN(n435) );
  XNOR2_X1 U455 ( .A(n441), .B(n363), .ZN(n663) );
  XNOR2_X1 U456 ( .A(n486), .B(n442), .ZN(n441) );
  XNOR2_X1 U457 ( .A(n443), .B(n481), .ZN(n442) );
  NAND2_X1 U458 ( .A1(G953), .A2(G900), .ZN(n757) );
  XNOR2_X1 U459 ( .A(n493), .B(n454), .ZN(n408) );
  XNOR2_X1 U460 ( .A(n461), .B(n410), .ZN(n409) );
  XNOR2_X1 U461 ( .A(n546), .B(n547), .ZN(n364) );
  XNOR2_X1 U462 ( .A(n440), .B(n438), .ZN(n763) );
  XNOR2_X1 U463 ( .A(n439), .B(KEYINPUT42), .ZN(n438) );
  INV_X1 U464 ( .A(KEYINPUT110), .ZN(n439) );
  AND2_X1 U465 ( .A1(n703), .A2(n447), .ZN(n446) );
  XNOR2_X1 U466 ( .A(n636), .B(n635), .ZN(n690) );
  XNOR2_X1 U467 ( .A(n368), .B(KEYINPUT107), .ZN(n762) );
  XNOR2_X1 U468 ( .A(n370), .B(KEYINPUT106), .ZN(n369) );
  NOR2_X1 U469 ( .A1(n564), .A2(n637), .ZN(n370) );
  AND2_X1 U470 ( .A1(n599), .A2(n581), .ZN(n686) );
  INV_X1 U471 ( .A(KEYINPUT56), .ZN(n385) );
  INV_X1 U472 ( .A(KEYINPUT53), .ZN(n405) );
  NAND2_X1 U473 ( .A1(n398), .A2(n397), .ZN(n406) );
  NAND2_X1 U474 ( .A1(n734), .A2(n401), .ZN(n397) );
  AND2_X1 U475 ( .A1(n650), .A2(n753), .ZN(n349) );
  XOR2_X1 U476 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n350) );
  INV_X1 U477 ( .A(n735), .ZN(n407) );
  AND2_X1 U478 ( .A1(n598), .A2(n757), .ZN(n351) );
  NAND2_X1 U479 ( .A1(n640), .A2(n639), .ZN(n352) );
  AND2_X1 U480 ( .A1(n633), .A2(n699), .ZN(n353) );
  NOR2_X1 U481 ( .A1(n637), .A2(n699), .ZN(n354) );
  NOR2_X1 U482 ( .A1(n716), .A2(n601), .ZN(n355) );
  AND2_X1 U483 ( .A1(n612), .A2(n630), .ZN(n356) );
  INV_X1 U484 ( .A(n374), .ZN(n723) );
  XOR2_X1 U485 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n357) );
  XNOR2_X1 U486 ( .A(n745), .B(n533), .ZN(n658) );
  XOR2_X1 U487 ( .A(n674), .B(n673), .Z(n358) );
  XOR2_X1 U488 ( .A(n666), .B(n665), .Z(n359) );
  XOR2_X1 U489 ( .A(n663), .B(n662), .Z(n360) );
  XOR2_X1 U490 ( .A(n658), .B(n660), .Z(n361) );
  INV_X1 U491 ( .A(n740), .ZN(n392) );
  NOR2_X1 U492 ( .A1(n746), .A2(G952), .ZN(n740) );
  XOR2_X1 U493 ( .A(KEYINPUT66), .B(KEYINPUT60), .Z(n362) );
  XNOR2_X1 U494 ( .A(n364), .B(n363), .ZN(n666) );
  XNOR2_X2 U495 ( .A(n526), .B(G134), .ZN(n515) );
  NAND2_X1 U496 ( .A1(n633), .A2(n627), .ZN(n367) );
  NAND2_X1 U497 ( .A1(n369), .A2(n615), .ZN(n368) );
  XNOR2_X1 U498 ( .A(n590), .B(KEYINPUT111), .ZN(n452) );
  NAND2_X1 U499 ( .A1(n433), .A2(n371), .ZN(n432) );
  INV_X1 U500 ( .A(n649), .ZN(n371) );
  XNOR2_X1 U501 ( .A(n649), .B(n372), .ZN(n754) );
  INV_X1 U502 ( .A(n755), .ZN(n372) );
  XNOR2_X2 U503 ( .A(n484), .B(n483), .ZN(n373) );
  XNOR2_X1 U504 ( .A(n373), .B(n485), .ZN(n486) );
  NAND2_X1 U505 ( .A1(n375), .A2(n374), .ZN(n614) );
  NAND2_X1 U506 ( .A1(n375), .A2(n355), .ZN(n602) );
  NAND2_X1 U507 ( .A1(n375), .A2(n353), .ZN(n636) );
  NAND2_X1 U508 ( .A1(n375), .A2(n354), .ZN(n638) );
  XNOR2_X2 U509 ( .A(n600), .B(n376), .ZN(n375) );
  XNOR2_X1 U510 ( .A(n556), .B(n377), .ZN(n599) );
  XNOR2_X2 U511 ( .A(n378), .B(n541), .ZN(n556) );
  NAND2_X1 U512 ( .A1(n577), .A2(n714), .ZN(n378) );
  NAND2_X1 U513 ( .A1(n381), .A2(n638), .ZN(n640) );
  AND2_X2 U514 ( .A1(n650), .A2(KEYINPUT84), .ZN(n433) );
  XNOR2_X1 U515 ( .A(n382), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U516 ( .A1(n389), .A2(n392), .ZN(n382) );
  XNOR2_X1 U517 ( .A(n383), .B(KEYINPUT123), .ZN(G54) );
  NAND2_X1 U518 ( .A1(n390), .A2(n392), .ZN(n383) );
  XNOR2_X1 U519 ( .A(n384), .B(n362), .ZN(G60) );
  NAND2_X1 U520 ( .A1(n391), .A2(n392), .ZN(n384) );
  XNOR2_X1 U521 ( .A(n386), .B(n385), .ZN(G51) );
  NAND2_X1 U522 ( .A1(n393), .A2(n392), .ZN(n386) );
  AND2_X1 U523 ( .A1(n352), .A2(n434), .ZN(n643) );
  NAND2_X1 U524 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X2 U525 ( .A(n602), .B(n436), .ZN(n610) );
  INV_X1 U526 ( .A(n622), .ZN(n625) );
  XNOR2_X1 U527 ( .A(n664), .B(n360), .ZN(n389) );
  XNOR2_X1 U528 ( .A(n667), .B(n359), .ZN(n390) );
  XNOR2_X1 U529 ( .A(n675), .B(n358), .ZN(n391) );
  XNOR2_X1 U530 ( .A(n661), .B(n361), .ZN(n393) );
  NAND2_X1 U531 ( .A1(n394), .A2(n626), .ZN(n645) );
  NAND2_X1 U532 ( .A1(n621), .A2(n622), .ZN(n394) );
  NOR2_X1 U533 ( .A1(n419), .A2(KEYINPUT48), .ZN(n421) );
  NAND2_X1 U534 ( .A1(n404), .A2(n403), .ZN(n402) );
  AND2_X1 U535 ( .A1(n407), .A2(KEYINPUT121), .ZN(n403) );
  INV_X1 U536 ( .A(n734), .ZN(n404) );
  XNOR2_X1 U537 ( .A(n406), .B(n405), .ZN(G75) );
  NAND2_X1 U538 ( .A1(n413), .A2(n412), .ZN(n411) );
  NAND2_X1 U539 ( .A1(n582), .A2(n351), .ZN(n414) );
  INV_X1 U540 ( .A(n437), .ZN(n415) );
  NOR2_X2 U541 ( .A1(n422), .A2(n416), .ZN(n753) );
  NAND2_X1 U542 ( .A1(n420), .A2(n417), .ZN(n416) );
  NAND2_X1 U543 ( .A1(n419), .A2(KEYINPUT48), .ZN(n418) );
  NAND2_X1 U544 ( .A1(n423), .A2(n421), .ZN(n420) );
  NOR2_X1 U545 ( .A1(n423), .A2(n587), .ZN(n422) );
  XNOR2_X1 U546 ( .A(n574), .B(n573), .ZN(n423) );
  NAND2_X1 U547 ( .A1(n582), .A2(n424), .ZN(n564) );
  NAND2_X1 U548 ( .A1(n562), .A2(n714), .ZN(n425) );
  XNOR2_X2 U549 ( .A(n539), .B(n538), .ZN(n577) );
  AND2_X2 U550 ( .A1(n429), .A2(n426), .ZN(n652) );
  NAND2_X1 U551 ( .A1(n428), .A2(n427), .ZN(n426) );
  NAND2_X1 U552 ( .A1(n430), .A2(n534), .ZN(n429) );
  NAND2_X1 U553 ( .A1(n432), .A2(n431), .ZN(n430) );
  INV_X1 U554 ( .A(KEYINPUT2), .ZN(n431) );
  XNOR2_X1 U555 ( .A(n434), .B(G101), .ZN(G3) );
  NAND2_X1 U556 ( .A1(n632), .A2(n631), .ZN(n434) );
  NAND2_X1 U557 ( .A1(n610), .A2(n435), .ZN(n629) );
  NAND2_X1 U558 ( .A1(n610), .A2(n356), .ZN(n668) );
  NAND2_X1 U559 ( .A1(n437), .A2(n714), .ZN(n719) );
  NOR2_X1 U560 ( .A1(n437), .A2(n714), .ZN(n715) );
  NAND2_X1 U561 ( .A1(n711), .A2(n581), .ZN(n440) );
  NAND2_X1 U562 ( .A1(n449), .A2(n446), .ZN(n445) );
  NAND2_X1 U563 ( .A1(n452), .A2(n450), .ZN(n449) );
  NOR2_X1 U564 ( .A1(n452), .A2(n543), .ZN(n451) );
  XOR2_X1 U565 ( .A(n522), .B(n521), .Z(n453) );
  XOR2_X1 U566 ( .A(n460), .B(n459), .Z(n454) );
  AND2_X1 U567 ( .A1(n598), .A2(n597), .ZN(n455) );
  BUF_X1 U568 ( .A(n526), .Z(n527) );
  INV_X1 U569 ( .A(KEYINPUT68), .ZN(n573) );
  INV_X1 U570 ( .A(KEYINPUT98), .ZN(n496) );
  XNOR2_X1 U571 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U572 ( .A(n499), .B(n498), .ZN(n502) );
  XNOR2_X1 U573 ( .A(KEYINPUT108), .B(KEYINPUT28), .ZN(n552) );
  XNOR2_X1 U574 ( .A(n553), .B(n552), .ZN(n555) );
  XNOR2_X1 U575 ( .A(n457), .B(n456), .ZN(n462) );
  NAND2_X1 U576 ( .A1(G221), .A2(n510), .ZN(n461) );
  XOR2_X1 U577 ( .A(KEYINPUT24), .B(KEYINPUT76), .Z(n460) );
  XNOR2_X1 U578 ( .A(G902), .B(KEYINPUT90), .ZN(n463) );
  XNOR2_X1 U579 ( .A(n463), .B(KEYINPUT15), .ZN(n651) );
  NAND2_X1 U580 ( .A1(G234), .A2(n651), .ZN(n464) );
  XNOR2_X1 U581 ( .A(n464), .B(KEYINPUT20), .ZN(n468) );
  NAND2_X1 U582 ( .A1(n468), .A2(G217), .ZN(n465) );
  AND2_X1 U583 ( .A1(n468), .A2(G221), .ZN(n471) );
  INV_X1 U584 ( .A(KEYINPUT93), .ZN(n469) );
  XNOR2_X1 U585 ( .A(n469), .B(KEYINPUT21), .ZN(n470) );
  XNOR2_X1 U586 ( .A(n471), .B(n470), .ZN(n697) );
  NAND2_X1 U587 ( .A1(G234), .A2(G237), .ZN(n473) );
  INV_X1 U588 ( .A(KEYINPUT14), .ZN(n472) );
  XNOR2_X1 U589 ( .A(n473), .B(n472), .ZN(n728) );
  OR2_X1 U590 ( .A1(G902), .A2(n746), .ZN(n474) );
  NAND2_X1 U591 ( .A1(n475), .A2(n474), .ZN(n476) );
  NOR2_X1 U592 ( .A1(n728), .A2(n476), .ZN(n598) );
  NAND2_X1 U593 ( .A1(n697), .A2(n351), .ZN(n477) );
  NOR2_X1 U594 ( .A1(n560), .A2(n477), .ZN(n551) );
  XNOR2_X2 U595 ( .A(G143), .B(G128), .ZN(n526) );
  XNOR2_X2 U596 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n530) );
  XOR2_X1 U597 ( .A(KEYINPUT94), .B(KEYINPUT5), .Z(n481) );
  NAND2_X1 U598 ( .A1(n500), .A2(G210), .ZN(n480) );
  XNOR2_X1 U599 ( .A(G101), .B(G131), .ZN(n485) );
  XNOR2_X1 U600 ( .A(G472), .B(KEYINPUT95), .ZN(n488) );
  INV_X1 U601 ( .A(KEYINPUT70), .ZN(n487) );
  XNOR2_X1 U602 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X2 U603 ( .A(n490), .B(n489), .ZN(n562) );
  NAND2_X1 U604 ( .A1(n551), .A2(n627), .ZN(n492) );
  XNOR2_X1 U605 ( .A(n492), .B(KEYINPUT103), .ZN(n519) );
  XOR2_X1 U606 ( .A(G131), .B(G140), .Z(n545) );
  XNOR2_X1 U607 ( .A(n495), .B(n494), .ZN(n499) );
  NAND2_X1 U608 ( .A1(G214), .A2(n500), .ZN(n501) );
  XNOR2_X1 U609 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U610 ( .A(n752), .B(n503), .Z(n674) );
  NOR2_X1 U611 ( .A1(G902), .A2(n674), .ZN(n506) );
  XNOR2_X1 U612 ( .A(KEYINPUT13), .B(KEYINPUT99), .ZN(n504) );
  INV_X1 U613 ( .A(KEYINPUT100), .ZN(n507) );
  XNOR2_X1 U614 ( .A(n576), .B(n507), .ZN(n557) );
  XOR2_X1 U615 ( .A(KEYINPUT7), .B(G122), .Z(n509) );
  XNOR2_X1 U616 ( .A(n509), .B(n508), .ZN(n514) );
  XOR2_X1 U617 ( .A(KEYINPUT9), .B(KEYINPUT101), .Z(n512) );
  NAND2_X1 U618 ( .A1(G217), .A2(n510), .ZN(n511) );
  XNOR2_X1 U619 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U620 ( .A(n514), .B(n513), .ZN(n516) );
  XNOR2_X1 U621 ( .A(n515), .B(n516), .ZN(n653) );
  INV_X1 U622 ( .A(G902), .ZN(n548) );
  NAND2_X1 U623 ( .A1(n653), .A2(n548), .ZN(n518) );
  INV_X1 U624 ( .A(G478), .ZN(n517) );
  XNOR2_X1 U625 ( .A(n518), .B(n517), .ZN(n575) );
  AND2_X2 U626 ( .A1(n557), .A2(n575), .ZN(n688) );
  XNOR2_X1 U627 ( .A(KEYINPUT71), .B(KEYINPUT16), .ZN(n522) );
  XNOR2_X1 U628 ( .A(G104), .B(G101), .ZN(n523) );
  NAND2_X1 U629 ( .A1(n746), .A2(G224), .ZN(n528) );
  XNOR2_X1 U630 ( .A(n528), .B(KEYINPUT77), .ZN(n529) );
  XNOR2_X1 U631 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U632 ( .A(n532), .B(n531), .ZN(n533) );
  INV_X1 U633 ( .A(n651), .ZN(n534) );
  NAND2_X1 U634 ( .A1(n548), .A2(n535), .ZN(n540) );
  NAND2_X1 U635 ( .A1(n540), .A2(G210), .ZN(n537) );
  INV_X1 U636 ( .A(KEYINPUT91), .ZN(n536) );
  XNOR2_X1 U637 ( .A(n537), .B(n536), .ZN(n538) );
  NAND2_X1 U638 ( .A1(n540), .A2(G214), .ZN(n714) );
  INV_X1 U639 ( .A(KEYINPUT88), .ZN(n541) );
  BUF_X1 U640 ( .A(n556), .Z(n542) );
  INV_X1 U641 ( .A(KEYINPUT36), .ZN(n543) );
  NAND2_X1 U642 ( .A1(G227), .A2(n746), .ZN(n544) );
  XNOR2_X1 U643 ( .A(n545), .B(n544), .ZN(n547) );
  NAND2_X1 U644 ( .A1(n666), .A2(n548), .ZN(n550) );
  XOR2_X1 U645 ( .A(KEYINPUT69), .B(G469), .Z(n549) );
  XNOR2_X2 U646 ( .A(n550), .B(n549), .ZN(n561) );
  XNOR2_X2 U647 ( .A(n561), .B(KEYINPUT1), .ZN(n703) );
  BUF_X2 U648 ( .A(n562), .Z(n699) );
  NAND2_X1 U649 ( .A1(n551), .A2(n699), .ZN(n553) );
  INV_X1 U650 ( .A(n561), .ZN(n554) );
  NOR2_X1 U651 ( .A1(n555), .A2(n554), .ZN(n581) );
  INV_X1 U652 ( .A(n688), .ZN(n584) );
  OR2_X1 U653 ( .A1(n557), .A2(n575), .ZN(n678) );
  AND2_X1 U654 ( .A1(n584), .A2(n678), .ZN(n718) );
  NOR2_X1 U655 ( .A1(n718), .A2(KEYINPUT47), .ZN(n558) );
  AND2_X1 U656 ( .A1(n686), .A2(n558), .ZN(n559) );
  INV_X1 U657 ( .A(n560), .ZN(n603) );
  INV_X1 U658 ( .A(n697), .ZN(n601) );
  NAND2_X1 U659 ( .A1(n561), .A2(n702), .ZN(n637) );
  XNOR2_X1 U660 ( .A(KEYINPUT105), .B(KEYINPUT30), .ZN(n563) );
  NOR2_X1 U661 ( .A1(n576), .A2(n575), .ZN(n615) );
  AND2_X1 U662 ( .A1(n718), .A2(KEYINPUT47), .ZN(n565) );
  NOR2_X1 U663 ( .A1(n762), .A2(n565), .ZN(n569) );
  INV_X1 U664 ( .A(n686), .ZN(n566) );
  NAND2_X1 U665 ( .A1(n566), .A2(KEYINPUT47), .ZN(n567) );
  XNOR2_X1 U666 ( .A(n567), .B(KEYINPUT82), .ZN(n568) );
  NAND2_X1 U667 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U668 ( .A(n570), .B(KEYINPUT81), .ZN(n571) );
  NAND2_X1 U669 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U670 ( .A1(n576), .A2(n575), .ZN(n716) );
  INV_X1 U671 ( .A(n577), .ZN(n592) );
  XNOR2_X1 U672 ( .A(KEYINPUT72), .B(KEYINPUT38), .ZN(n578) );
  NOR2_X1 U673 ( .A1(n716), .A2(n719), .ZN(n580) );
  XNOR2_X1 U674 ( .A(KEYINPUT41), .B(KEYINPUT109), .ZN(n579) );
  INV_X1 U675 ( .A(KEYINPUT39), .ZN(n583) );
  NOR2_X1 U676 ( .A1(n594), .A2(n584), .ZN(n585) );
  XNOR2_X1 U677 ( .A(n585), .B(KEYINPUT40), .ZN(n764) );
  NOR2_X1 U678 ( .A1(n763), .A2(n764), .ZN(n586) );
  INV_X1 U679 ( .A(KEYINPUT48), .ZN(n587) );
  INV_X1 U680 ( .A(n714), .ZN(n588) );
  OR2_X1 U681 ( .A1(n703), .A2(n588), .ZN(n589) );
  OR2_X1 U682 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U683 ( .A(n591), .B(KEYINPUT43), .ZN(n593) );
  NAND2_X1 U684 ( .A1(n593), .A2(n592), .ZN(n670) );
  OR2_X1 U685 ( .A1(n678), .A2(n594), .ZN(n694) );
  AND2_X1 U686 ( .A1(n670), .A2(n694), .ZN(n595) );
  NAND2_X1 U687 ( .A1(n753), .A2(KEYINPUT2), .ZN(n596) );
  XNOR2_X1 U688 ( .A(n596), .B(KEYINPUT85), .ZN(n647) );
  NAND2_X1 U689 ( .A1(G953), .A2(G898), .ZN(n597) );
  NAND2_X1 U690 ( .A1(n599), .A2(n455), .ZN(n600) );
  INV_X1 U691 ( .A(n703), .ZN(n630) );
  INV_X1 U692 ( .A(n603), .ZN(n696) );
  NOR2_X1 U693 ( .A1(n630), .A2(n696), .ZN(n604) );
  XOR2_X1 U694 ( .A(KEYINPUT102), .B(n604), .Z(n606) );
  XNOR2_X1 U695 ( .A(n388), .B(KEYINPUT80), .ZN(n605) );
  NOR2_X1 U696 ( .A1(n606), .A2(n605), .ZN(n608) );
  INV_X1 U697 ( .A(KEYINPUT79), .ZN(n607) );
  XNOR2_X1 U698 ( .A(n608), .B(n607), .ZN(n609) );
  XNOR2_X2 U699 ( .A(n611), .B(KEYINPUT32), .ZN(n669) );
  NOR2_X1 U700 ( .A1(n696), .A2(n699), .ZN(n612) );
  INV_X1 U701 ( .A(KEYINPUT34), .ZN(n613) );
  XNOR2_X1 U702 ( .A(n614), .B(n613), .ZN(n617) );
  XNOR2_X1 U703 ( .A(n615), .B(KEYINPUT78), .ZN(n616) );
  NAND2_X1 U704 ( .A1(n617), .A2(n616), .ZN(n619) );
  INV_X1 U705 ( .A(KEYINPUT35), .ZN(n618) );
  XNOR2_X2 U706 ( .A(n619), .B(n618), .ZN(n761) );
  NAND2_X1 U707 ( .A1(n761), .A2(KEYINPUT87), .ZN(n620) );
  INV_X1 U708 ( .A(KEYINPUT44), .ZN(n641) );
  AND2_X1 U709 ( .A1(n620), .A2(n641), .ZN(n621) );
  NOR2_X1 U710 ( .A1(KEYINPUT44), .A2(KEYINPUT87), .ZN(n623) );
  NAND2_X1 U711 ( .A1(n761), .A2(n623), .ZN(n624) );
  NAND2_X1 U712 ( .A1(n625), .A2(n624), .ZN(n626) );
  INV_X1 U713 ( .A(KEYINPUT86), .ZN(n628) );
  XNOR2_X1 U714 ( .A(n629), .B(n628), .ZN(n632) );
  AND2_X1 U715 ( .A1(n696), .A2(n630), .ZN(n631) );
  XNOR2_X1 U716 ( .A(KEYINPUT96), .B(KEYINPUT97), .ZN(n634) );
  XOR2_X1 U717 ( .A(n634), .B(KEYINPUT31), .Z(n635) );
  INV_X1 U718 ( .A(n638), .ZN(n679) );
  INV_X1 U719 ( .A(n718), .ZN(n639) );
  OR2_X1 U720 ( .A1(n761), .A2(n641), .ZN(n642) );
  XNOR2_X2 U721 ( .A(n646), .B(KEYINPUT45), .ZN(n650) );
  NAND2_X1 U722 ( .A1(n647), .A2(n650), .ZN(n648) );
  XNOR2_X2 U723 ( .A(n648), .B(KEYINPUT75), .ZN(n733) );
  INV_X1 U724 ( .A(n753), .ZN(n649) );
  NOR2_X4 U725 ( .A1(n733), .A2(n652), .ZN(n736) );
  NAND2_X1 U726 ( .A1(n736), .A2(G478), .ZN(n654) );
  XNOR2_X1 U727 ( .A(n654), .B(n653), .ZN(n655) );
  NAND2_X1 U728 ( .A1(n655), .A2(n392), .ZN(n657) );
  INV_X1 U729 ( .A(KEYINPUT124), .ZN(n656) );
  XNOR2_X1 U730 ( .A(n657), .B(n656), .ZN(G63) );
  NAND2_X1 U731 ( .A1(n736), .A2(G210), .ZN(n661) );
  XOR2_X1 U732 ( .A(KEYINPUT122), .B(KEYINPUT54), .Z(n659) );
  XNOR2_X1 U733 ( .A(n659), .B(KEYINPUT55), .ZN(n660) );
  NAND2_X1 U734 ( .A1(n736), .A2(G472), .ZN(n664) );
  XNOR2_X1 U735 ( .A(KEYINPUT112), .B(KEYINPUT62), .ZN(n662) );
  NAND2_X1 U736 ( .A1(n736), .A2(G469), .ZN(n667) );
  XNOR2_X1 U737 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n665) );
  XNOR2_X1 U738 ( .A(n668), .B(G110), .ZN(G12) );
  XNOR2_X1 U739 ( .A(n669), .B(G119), .ZN(G21) );
  XNOR2_X1 U740 ( .A(n670), .B(G140), .ZN(G42) );
  XOR2_X1 U741 ( .A(G125), .B(KEYINPUT37), .Z(n672) );
  XOR2_X1 U742 ( .A(n672), .B(n671), .Z(G27) );
  NAND2_X1 U743 ( .A1(n736), .A2(G475), .ZN(n675) );
  XNOR2_X1 U744 ( .A(KEYINPUT89), .B(KEYINPUT59), .ZN(n673) );
  XOR2_X1 U745 ( .A(G104), .B(KEYINPUT113), .Z(n677) );
  NAND2_X1 U746 ( .A1(n679), .A2(n688), .ZN(n676) );
  XNOR2_X1 U747 ( .A(n677), .B(n676), .ZN(G6) );
  XNOR2_X1 U748 ( .A(G107), .B(KEYINPUT27), .ZN(n683) );
  XOR2_X1 U749 ( .A(KEYINPUT114), .B(KEYINPUT26), .Z(n681) );
  INV_X1 U750 ( .A(n678), .ZN(n691) );
  NAND2_X1 U751 ( .A1(n679), .A2(n691), .ZN(n680) );
  XNOR2_X1 U752 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U753 ( .A(n683), .B(n682), .ZN(G9) );
  XOR2_X1 U754 ( .A(G128), .B(KEYINPUT29), .Z(n685) );
  NAND2_X1 U755 ( .A1(n686), .A2(n691), .ZN(n684) );
  XNOR2_X1 U756 ( .A(n685), .B(n684), .ZN(G30) );
  NAND2_X1 U757 ( .A1(n686), .A2(n688), .ZN(n687) );
  XNOR2_X1 U758 ( .A(n687), .B(G146), .ZN(G48) );
  NAND2_X1 U759 ( .A1(n690), .A2(n688), .ZN(n689) );
  XNOR2_X1 U760 ( .A(n689), .B(G113), .ZN(G15) );
  XOR2_X1 U761 ( .A(G116), .B(KEYINPUT115), .Z(n693) );
  NAND2_X1 U762 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U763 ( .A(n693), .B(n692), .ZN(G18) );
  INV_X1 U764 ( .A(n694), .ZN(n695) );
  XOR2_X1 U765 ( .A(G134), .B(n695), .Z(G36) );
  NOR2_X1 U766 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U767 ( .A(KEYINPUT49), .B(n698), .Z(n700) );
  NOR2_X1 U768 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U769 ( .A(n701), .B(KEYINPUT116), .Z(n707) );
  NOR2_X1 U770 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U771 ( .A(KEYINPUT117), .B(n704), .Z(n705) );
  XNOR2_X1 U772 ( .A(KEYINPUT50), .B(n705), .ZN(n706) );
  NOR2_X1 U773 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U774 ( .A(n708), .B(KEYINPUT118), .ZN(n709) );
  NOR2_X1 U775 ( .A1(n709), .A2(n353), .ZN(n710) );
  XNOR2_X1 U776 ( .A(KEYINPUT51), .B(n710), .ZN(n712) );
  NAND2_X1 U777 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U778 ( .A(n713), .B(KEYINPUT119), .ZN(n725) );
  NOR2_X1 U779 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U780 ( .A(n717), .B(KEYINPUT120), .ZN(n721) );
  NOR2_X1 U781 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U782 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U783 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U784 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U785 ( .A(n726), .B(KEYINPUT52), .ZN(n727) );
  NOR2_X1 U786 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U787 ( .A1(n729), .A2(G952), .ZN(n730) );
  NAND2_X1 U788 ( .A1(n731), .A2(n730), .ZN(n735) );
  NOR2_X1 U789 ( .A1(n349), .A2(KEYINPUT2), .ZN(n732) );
  NOR2_X1 U790 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U791 ( .A1(n736), .A2(G217), .ZN(n738) );
  XNOR2_X1 U792 ( .A(n738), .B(n737), .ZN(n739) );
  NOR2_X1 U793 ( .A1(n740), .A2(n739), .ZN(G66) );
  NAND2_X1 U794 ( .A1(n650), .A2(n746), .ZN(n744) );
  NAND2_X1 U795 ( .A1(G953), .A2(G224), .ZN(n741) );
  XNOR2_X1 U796 ( .A(KEYINPUT61), .B(n741), .ZN(n742) );
  NAND2_X1 U797 ( .A1(n742), .A2(G898), .ZN(n743) );
  NAND2_X1 U798 ( .A1(n744), .A2(n743), .ZN(n750) );
  XNOR2_X1 U799 ( .A(n745), .B(KEYINPUT125), .ZN(n748) );
  NOR2_X1 U800 ( .A1(G898), .A2(n746), .ZN(n747) );
  NOR2_X1 U801 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U802 ( .A(n750), .B(n749), .ZN(G69) );
  XNOR2_X1 U803 ( .A(n751), .B(n752), .ZN(n755) );
  NOR2_X1 U804 ( .A1(n754), .A2(G953), .ZN(n759) );
  XNOR2_X1 U805 ( .A(n755), .B(G227), .ZN(n756) );
  NOR2_X1 U806 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X1 U807 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U808 ( .A(KEYINPUT126), .B(n760), .ZN(G72) );
  XNOR2_X1 U809 ( .A(n761), .B(G122), .ZN(G24) );
  XOR2_X1 U810 ( .A(G143), .B(n762), .Z(G45) );
  XOR2_X1 U811 ( .A(G137), .B(n763), .Z(G39) );
  XOR2_X1 U812 ( .A(G131), .B(n764), .Z(G33) );
endmodule

