//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n851, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944;
  XNOR2_X1  g000(.A(KEYINPUT76), .B(KEYINPUT34), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT73), .ZN(new_n203));
  INV_X1    g002(.A(G134gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT72), .ZN(new_n205));
  INV_X1    g004(.A(G127gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(KEYINPUT72), .A2(G127gat), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n204), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(G127gat), .A2(G134gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n203), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n208), .ZN(new_n212));
  NOR2_X1   g011(.A1(KEYINPUT72), .A2(G127gat), .ZN(new_n213));
  OAI21_X1  g012(.A(G134gat), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n210), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n214), .A2(KEYINPUT73), .A3(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G120gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G113gat), .ZN(new_n218));
  INV_X1    g017(.A(G113gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G120gat), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT1), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n211), .A2(new_n216), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n218), .A2(KEYINPUT74), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT74), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(new_n217), .A3(G113gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n220), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G127gat), .A2(G134gat), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT1), .B1(new_n215), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  AND2_X1   g029(.A1(new_n223), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(KEYINPUT27), .B(G183gat), .ZN(new_n232));
  INV_X1    g031(.A(G190gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(KEYINPUT70), .A2(KEYINPUT28), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n234), .B1(new_n232), .B2(new_n233), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT26), .ZN(new_n239));
  INV_X1    g038(.A(G169gat), .ZN(new_n240));
  INV_X1    g039(.A(G176gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n243));
  AND3_X1   g042(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n242), .B(new_n243), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G183gat), .A2(G190gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(KEYINPUT71), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT71), .B1(new_n246), .B2(new_n247), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n238), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT64), .ZN(new_n252));
  NAND3_X1  g051(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n253), .B1(G183gat), .B2(G190gat), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n252), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n255), .ZN(new_n257));
  OR2_X1    g056(.A1(G183gat), .A2(G190gat), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n257), .A2(new_n258), .A3(KEYINPUT64), .A4(new_n253), .ZN(new_n259));
  NAND2_X1  g058(.A1(G169gat), .A2(G176gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT66), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n240), .A2(new_n241), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT23), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n262), .A2(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OR2_X1    g065(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n267), .A2(KEYINPUT23), .A3(new_n241), .A4(new_n268), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n256), .A2(new_n259), .A3(new_n266), .A4(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT25), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT24), .B1(new_n247), .B2(KEYINPUT67), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT67), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n273), .A2(G183gat), .A3(G190gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n253), .A2(KEYINPUT68), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n253), .A2(KEYINPUT68), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n275), .B(new_n258), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  OAI22_X1  g078(.A1(new_n244), .A2(new_n245), .B1(KEYINPUT23), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT25), .B1(new_n264), .B2(new_n265), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI22_X1  g081(.A1(new_n270), .A2(new_n271), .B1(new_n278), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n251), .B1(new_n283), .B2(KEYINPUT69), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n270), .A2(new_n271), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n278), .A2(new_n282), .ZN(new_n286));
  AND3_X1   g085(.A1(new_n285), .A2(KEYINPUT69), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n231), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n285), .A2(new_n286), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT69), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n223), .A2(new_n230), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n283), .A2(KEYINPUT69), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n291), .A2(new_n292), .A3(new_n251), .A4(new_n293), .ZN(new_n294));
  AND2_X1   g093(.A1(new_n288), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G227gat), .ZN(new_n296));
  INV_X1    g095(.A(G233gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n202), .B1(new_n295), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT77), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n288), .A2(new_n294), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n298), .A2(KEYINPUT34), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n302), .ZN(new_n304));
  AOI211_X1 g103(.A(KEYINPUT77), .B(new_n304), .C1(new_n288), .C2(new_n294), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n299), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n288), .A2(new_n294), .A3(new_n298), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT32), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT33), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G15gat), .B(G43gat), .ZN(new_n311));
  INV_X1    g110(.A(G71gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n313), .B(KEYINPUT75), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n314), .B(G99gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n310), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n308), .B1(new_n315), .B2(KEYINPUT33), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(new_n307), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n306), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT77), .B1(new_n295), .B2(new_n304), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n301), .A2(new_n300), .A3(new_n302), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n310), .A2(new_n315), .B1(new_n307), .B2(new_n317), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(new_n324), .A3(new_n299), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT79), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n320), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT79), .A4(new_n299), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G226gat), .A2(G233gat), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n291), .A2(new_n331), .A3(new_n251), .A4(new_n293), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n289), .A2(new_n251), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n331), .A2(KEYINPUT29), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT22), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT80), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT80), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT22), .ZN(new_n340));
  NAND2_X1  g139(.A1(G211gat), .A2(G218gat), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n338), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT81), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT81), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n338), .A2(new_n340), .A3(new_n344), .A4(new_n341), .ZN(new_n345));
  AND2_X1   g144(.A1(G197gat), .A2(G204gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(G197gat), .A2(G204gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n343), .A2(new_n345), .A3(new_n349), .ZN(new_n350));
  XOR2_X1   g149(.A(G211gat), .B(G218gat), .Z(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n348), .B1(new_n342), .B2(KEYINPUT81), .ZN(new_n353));
  INV_X1    g152(.A(new_n351), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n353), .A2(new_n354), .A3(new_n345), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n336), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G8gat), .B(G36gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(G64gat), .ZN(new_n359));
  INV_X1    g158(.A(G92gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n334), .B1(new_n284), .B2(new_n287), .ZN(new_n362));
  AND4_X1   g161(.A1(new_n354), .A2(new_n343), .A3(new_n345), .A4(new_n349), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n354), .B1(new_n353), .B2(new_n345), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n289), .A2(new_n251), .A3(new_n331), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n362), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n357), .A2(new_n361), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT30), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n357), .A2(KEYINPUT30), .A3(new_n361), .A4(new_n367), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT82), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n362), .A2(new_n365), .A3(new_n366), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n365), .B1(new_n332), .B2(new_n335), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n357), .A2(KEYINPUT82), .A3(new_n367), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n361), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NOR3_X1   g177(.A1(new_n372), .A2(new_n378), .A3(KEYINPUT35), .ZN(new_n379));
  NAND2_X1  g178(.A1(G155gat), .A2(G162gat), .ZN(new_n380));
  INV_X1    g179(.A(G155gat), .ZN(new_n381));
  INV_X1    g180(.A(G162gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n380), .B1(new_n383), .B2(KEYINPUT2), .ZN(new_n384));
  INV_X1    g183(.A(G148gat), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n385), .A2(KEYINPUT84), .A3(G141gat), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n386), .B1(G141gat), .B2(new_n385), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT84), .B1(new_n385), .B2(G141gat), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n384), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AND2_X1   g188(.A1(G155gat), .A2(G162gat), .ZN(new_n390));
  NOR2_X1   g189(.A1(G155gat), .A2(G162gat), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT83), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT83), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n383), .A2(new_n393), .A3(new_n380), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n380), .A2(KEYINPUT2), .ZN(new_n395));
  XNOR2_X1  g194(.A(G141gat), .B(G148gat), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n392), .B(new_n394), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n389), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n398), .A2(new_n223), .A3(new_n230), .ZN(new_n399));
  NAND2_X1  g198(.A1(G225gat), .A2(G233gat), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n389), .A2(new_n397), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n403), .B1(new_n389), .B2(new_n397), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n292), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n408), .B1(new_n231), .B2(new_n398), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n398), .A2(new_n223), .A3(new_n408), .A4(new_n230), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n402), .B(new_n407), .C1(new_n409), .C2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT5), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n389), .A2(new_n397), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n292), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n399), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n413), .B1(new_n416), .B2(new_n401), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n399), .A2(KEYINPUT4), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n418), .A2(new_n410), .B1(new_n292), .B2(new_n406), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n401), .A2(KEYINPUT5), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n412), .A2(new_n417), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(G1gat), .B(G29gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(KEYINPUT0), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(G57gat), .ZN(new_n424));
  INV_X1    g223(.A(G85gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n421), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT6), .ZN(new_n428));
  INV_X1    g227(.A(new_n426), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n412), .A2(new_n417), .ZN(new_n430));
  AND2_X1   g229(.A1(new_n419), .A2(new_n420), .ZN(new_n431));
  OAI211_X1 g230(.A(KEYINPUT89), .B(new_n429), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT89), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n433), .B1(new_n421), .B2(new_n426), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT6), .B1(new_n421), .B2(new_n426), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n432), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT29), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n437), .B1(new_n414), .B2(KEYINPUT3), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n365), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n439), .A2(G228gat), .A3(G233gat), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n437), .B1(new_n363), .B2(new_n364), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT85), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g242(.A(KEYINPUT85), .B(new_n437), .C1(new_n363), .C2(new_n364), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n403), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n440), .B1(new_n445), .B2(new_n414), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n405), .B1(new_n365), .B2(new_n438), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT29), .B1(new_n352), .B2(new_n355), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n414), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n447), .A2(new_n449), .B1(G228gat), .B2(G233gat), .ZN(new_n450));
  OAI21_X1  g249(.A(G22gat), .B1(new_n446), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n447), .A2(new_n449), .ZN(new_n452));
  NAND2_X1  g251(.A1(G228gat), .A2(G233gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(G22gat), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT3), .B1(new_n448), .B2(KEYINPUT85), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n398), .B1(new_n456), .B2(new_n443), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n454), .B(new_n455), .C1(new_n457), .C2(new_n440), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n451), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n454), .B1(new_n457), .B2(new_n440), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT86), .B1(new_n460), .B2(G22gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(G78gat), .B(G106gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(KEYINPUT31), .B(G50gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n462), .B(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n459), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n451), .A2(KEYINPUT86), .A3(new_n458), .A4(new_n464), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n428), .A2(new_n436), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n329), .A2(new_n379), .A3(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n372), .A2(new_n378), .ZN(new_n470));
  INV_X1    g269(.A(new_n435), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n428), .B1(new_n471), .B2(new_n427), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  AND4_X1   g272(.A1(KEYINPUT86), .A2(new_n451), .A3(new_n458), .A4(new_n464), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT86), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n444), .A2(new_n403), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT85), .B1(new_n356), .B2(new_n437), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n414), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n453), .B1(new_n365), .B2(new_n438), .ZN(new_n479));
  AOI22_X1  g278(.A1(new_n478), .A2(new_n479), .B1(new_n452), .B2(new_n453), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n475), .B1(new_n480), .B2(new_n455), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n481), .A2(new_n464), .B1(new_n458), .B2(new_n451), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n320), .B(new_n325), .C1(new_n474), .C2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT35), .B1(new_n473), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n407), .B1(new_n409), .B2(new_n411), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(new_n401), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n415), .A2(new_n400), .A3(new_n399), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n488), .A2(KEYINPUT39), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n429), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT39), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n486), .A2(new_n491), .A3(new_n401), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT40), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n489), .B1(new_n400), .B2(new_n419), .ZN(new_n494));
  AND4_X1   g293(.A1(KEYINPUT40), .A2(new_n494), .A3(new_n426), .A4(new_n492), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n432), .A2(new_n434), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n496), .B(new_n497), .C1(new_n378), .C2(new_n372), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n466), .A2(new_n467), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT38), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT37), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT37), .B1(new_n357), .B2(new_n367), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n361), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n500), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n332), .A2(new_n365), .A3(new_n335), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n365), .B1(new_n362), .B2(new_n366), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT37), .ZN(new_n509));
  NOR3_X1   g308(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n500), .B(new_n505), .C1(new_n510), .C2(new_n502), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n511), .A2(new_n436), .A3(new_n428), .A4(new_n368), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n498), .B(new_n499), .C1(new_n506), .C2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT78), .B(KEYINPUT36), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n327), .A2(new_n328), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n320), .A2(new_n325), .A3(KEYINPUT36), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT87), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n517), .B1(new_n482), .B2(new_n474), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n466), .A2(KEYINPUT87), .A3(new_n467), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n515), .A2(new_n516), .B1(new_n520), .B2(new_n473), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n513), .B1(new_n521), .B2(KEYINPUT88), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n515), .A2(new_n516), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n520), .A2(new_n473), .ZN(new_n524));
  AND3_X1   g323(.A1(new_n523), .A2(KEYINPUT88), .A3(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n485), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(G8gat), .ZN(new_n527));
  INV_X1    g326(.A(G1gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT16), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT92), .ZN(new_n530));
  XNOR2_X1  g329(.A(G15gat), .B(G22gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT93), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n527), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n532), .B1(G1gat), .B2(new_n531), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI221_X1 g335(.A(new_n532), .B1(new_n533), .B2(new_n527), .C1(G1gat), .C2(new_n531), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G43gat), .B(G50gat), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n540), .A2(KEYINPUT15), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(KEYINPUT15), .ZN(new_n542));
  NAND2_X1  g341(.A1(G29gat), .A2(G36gat), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT14), .ZN(new_n544));
  INV_X1    g343(.A(G29gat), .ZN(new_n545));
  INV_X1    g344(.A(G36gat), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n541), .A2(new_n542), .A3(new_n543), .A4(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n548), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT91), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n551), .B1(new_n547), .B2(new_n552), .ZN(new_n553));
  OR2_X1    g352(.A1(new_n547), .A2(new_n552), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n553), .A2(new_n554), .B1(G29gat), .B2(G36gat), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n550), .B1(new_n555), .B2(new_n542), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT17), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n557), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n539), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G229gat), .A2(G233gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n538), .A2(new_n556), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT18), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n538), .B(new_n556), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n561), .B(KEYINPUT13), .Z(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AND2_X1   g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n560), .A2(new_n562), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n570), .A2(KEYINPUT18), .A3(new_n561), .ZN(new_n571));
  AOI21_X1  g370(.A(KEYINPUT94), .B1(new_n563), .B2(new_n564), .ZN(new_n572));
  XOR2_X1   g371(.A(KEYINPUT90), .B(KEYINPUT11), .Z(new_n573));
  XNOR2_X1  g372(.A(G113gat), .B(G141gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G169gat), .B(G197gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT12), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n569), .B(new_n571), .C1(new_n572), .C2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n571), .A2(new_n565), .A3(new_n568), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n572), .A2(new_n578), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n526), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(G64gat), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n585), .A2(G57gat), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n585), .A2(G57gat), .ZN(new_n587));
  INV_X1    g386(.A(G78gat), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n312), .A2(new_n588), .ZN(new_n589));
  OAI22_X1  g388(.A1(new_n586), .A2(new_n587), .B1(new_n589), .B2(KEYINPUT9), .ZN(new_n590));
  XNOR2_X1  g389(.A(G71gat), .B(G78gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT21), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G127gat), .B(G155gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT95), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n597), .B(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n539), .B1(new_n594), .B2(new_n593), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT96), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n600), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G183gat), .B(G211gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n600), .A2(new_n602), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n600), .A2(new_n602), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n609), .A2(new_n606), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G85gat), .A2(G92gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT7), .ZN(new_n615));
  NAND2_X1  g414(.A1(G99gat), .A2(G106gat), .ZN(new_n616));
  AOI22_X1  g415(.A1(KEYINPUT8), .A2(new_n616), .B1(new_n425), .B2(new_n360), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G99gat), .B(G106gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n558), .A2(new_n559), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n620), .ZN(new_n622));
  AND2_X1   g421(.A1(G232gat), .A2(G233gat), .ZN(new_n623));
  AOI22_X1  g422(.A1(new_n622), .A2(new_n556), .B1(KEYINPUT41), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G190gat), .B(G218gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(G134gat), .B(G162gat), .Z(new_n628));
  NOR2_X1   g427(.A1(new_n623), .A2(KEYINPUT41), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n631), .A2(KEYINPUT97), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(KEYINPUT97), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n627), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(G230gat), .A2(G233gat), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n638), .B(KEYINPUT100), .Z(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n618), .A2(KEYINPUT98), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT99), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n619), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n619), .A2(new_n642), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n618), .B1(KEYINPUT98), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n592), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n620), .A2(new_n593), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n640), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n648), .B(KEYINPUT101), .Z(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n646), .A2(new_n650), .A3(new_n647), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n622), .A2(KEYINPUT10), .A3(new_n592), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n639), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G120gat), .B(G148gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G176gat), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n657), .B(G204gat), .Z(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n649), .A2(new_n658), .A3(new_n654), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n613), .A2(new_n637), .A3(new_n662), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n584), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n472), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT102), .B(G1gat), .Z(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(G1324gat));
  INV_X1    g467(.A(new_n470), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT16), .B(G8gat), .Z(new_n670));
  NAND4_X1  g469(.A1(new_n664), .A2(KEYINPUT42), .A3(new_n669), .A4(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT42), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT103), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n664), .A2(new_n673), .A3(new_n669), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n584), .A2(new_n669), .A3(new_n663), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT103), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n670), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n672), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(KEYINPUT104), .B1(new_n677), .B2(G8gat), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n681));
  AOI211_X1 g480(.A(new_n681), .B(new_n527), .C1(new_n674), .C2(new_n676), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n671), .B(new_n679), .C1(new_n680), .C2(new_n682), .ZN(G1325gat));
  INV_X1    g482(.A(new_n664), .ZN(new_n684));
  OAI21_X1  g483(.A(G15gat), .B1(new_n684), .B2(new_n523), .ZN(new_n685));
  INV_X1    g484(.A(new_n329), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n686), .A2(G15gat), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n685), .B1(new_n684), .B2(new_n687), .ZN(G1326gat));
  NAND2_X1  g487(.A1(new_n664), .A2(new_n520), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT43), .B(G22gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1327gat));
  NOR2_X1   g490(.A1(new_n612), .A2(new_n662), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n637), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n584), .A2(new_n545), .A3(new_n665), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT45), .ZN(new_n696));
  INV_X1    g495(.A(new_n692), .ZN(new_n697));
  INV_X1    g496(.A(new_n583), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AOI22_X1  g498(.A1(new_n521), .A2(new_n513), .B1(new_n484), .B2(new_n469), .ZN(new_n700));
  XOR2_X1   g499(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n701));
  NOR4_X1   g500(.A1(new_n700), .A2(KEYINPUT106), .A3(new_n636), .A4(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n523), .A2(new_n513), .A3(new_n524), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n636), .B1(new_n704), .B2(new_n485), .ZN(new_n705));
  INV_X1    g504(.A(new_n701), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n703), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n709), .B1(new_n526), .B2(new_n637), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n699), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(G29gat), .B1(new_n711), .B2(new_n472), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n712), .ZN(G1328gat));
  NAND4_X1  g512(.A1(new_n584), .A2(new_n546), .A3(new_n669), .A4(new_n694), .ZN(new_n714));
  XOR2_X1   g513(.A(KEYINPUT107), .B(KEYINPUT46), .Z(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(G36gat), .B1(new_n711), .B2(new_n470), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(G1329gat));
  OAI21_X1  g517(.A(G43gat), .B1(new_n711), .B2(new_n523), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n693), .A2(G43gat), .A3(new_n686), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n584), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT47), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1330gat));
  OAI21_X1  g523(.A(G50gat), .B1(new_n711), .B2(new_n499), .ZN(new_n725));
  INV_X1    g524(.A(new_n520), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n693), .A2(new_n726), .A3(G50gat), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n584), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n725), .A2(KEYINPUT48), .A3(new_n728), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n520), .B(new_n699), .C1(new_n708), .C2(new_n710), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n730), .A2(KEYINPUT108), .A3(G50gat), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT108), .B1(new_n730), .B2(G50gat), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n728), .A2(KEYINPUT109), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT109), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n584), .A2(new_n734), .A3(new_n727), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n731), .A2(new_n732), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n729), .B1(new_n737), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g537(.A1(new_n612), .A2(new_n698), .A3(new_n636), .A4(new_n662), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT110), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n704), .A2(new_n485), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OR2_X1    g541(.A1(new_n742), .A2(KEYINPUT111), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(KEYINPUT111), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n745), .A2(new_n472), .ZN(new_n746));
  XOR2_X1   g545(.A(KEYINPUT112), .B(G57gat), .Z(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1332gat));
  AND2_X1   g547(.A1(new_n743), .A2(new_n744), .ZN(new_n749));
  NOR2_X1   g548(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n749), .A2(new_n669), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(KEYINPUT113), .B(KEYINPUT114), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n669), .A2(new_n752), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n750), .B1(new_n745), .B2(new_n755), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n753), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n754), .B1(new_n753), .B2(new_n756), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(G1333gat));
  INV_X1    g558(.A(new_n523), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n749), .A2(G71gat), .A3(new_n760), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n329), .B(KEYINPUT115), .Z(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n312), .B1(new_n745), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT50), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n761), .A2(new_n767), .A3(new_n764), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(G1334gat));
  NOR2_X1   g568(.A1(new_n745), .A2(new_n726), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(new_n588), .ZN(G1335gat));
  NOR2_X1   g570(.A1(new_n612), .A2(new_n583), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n705), .A2(new_n772), .ZN(new_n773));
  OR2_X1    g572(.A1(new_n773), .A2(KEYINPUT51), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(KEYINPUT51), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n774), .A2(new_n662), .A3(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n776), .A2(new_n425), .A3(new_n665), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n708), .A2(new_n710), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n772), .A2(new_n662), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n778), .A2(new_n472), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n777), .B1(new_n780), .B2(new_n425), .ZN(G1336gat));
  INV_X1    g580(.A(new_n779), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n669), .B(new_n782), .C1(new_n708), .C2(new_n710), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G92gat), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n470), .A2(G92gat), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n776), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT116), .ZN(new_n788));
  OR2_X1    g587(.A1(new_n788), .A2(KEYINPUT52), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(KEYINPUT52), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n787), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n784), .A2(new_n786), .A3(new_n788), .A4(KEYINPUT52), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(G1337gat));
  AOI21_X1  g592(.A(G99gat), .B1(new_n776), .B2(new_n329), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n760), .A2(G99gat), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(G1338gat));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n520), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n499), .A2(G106gat), .ZN(new_n799));
  AOI22_X1  g598(.A1(new_n798), .A2(G106gat), .B1(new_n776), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n776), .A2(new_n799), .ZN(new_n802));
  XNOR2_X1  g601(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(G106gat), .ZN(new_n805));
  INV_X1    g604(.A(new_n499), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n805), .B1(new_n795), .B2(new_n806), .ZN(new_n807));
  OAI22_X1  g606(.A1(new_n800), .A2(new_n801), .B1(new_n804), .B2(new_n807), .ZN(G1339gat));
  NAND3_X1  g607(.A1(new_n651), .A2(new_n639), .A3(new_n652), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n654), .A2(KEYINPUT54), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n658), .B1(new_n653), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n812), .A2(KEYINPUT118), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n812), .A2(KEYINPUT118), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n810), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g616(.A(KEYINPUT55), .B(new_n810), .C1(new_n813), .C2(new_n814), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n817), .A2(new_n583), .A3(new_n661), .A4(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n570), .A2(new_n561), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n566), .A2(new_n567), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n577), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n569), .A2(new_n578), .A3(new_n571), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n662), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n637), .B1(new_n819), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n817), .A2(new_n661), .A3(new_n818), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n637), .A2(new_n822), .A3(new_n823), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n613), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n663), .A2(new_n698), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n472), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n483), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT119), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT119), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n831), .A2(new_n835), .A3(new_n832), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n669), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n837), .A2(KEYINPUT120), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n837), .A2(KEYINPUT120), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n219), .B(new_n583), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n520), .B1(new_n829), .B2(new_n830), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n841), .A2(new_n665), .A3(new_n470), .A4(new_n329), .ZN(new_n842));
  OAI21_X1  g641(.A(G113gat), .B1(new_n842), .B2(new_n698), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n840), .A2(new_n843), .ZN(G1340gat));
  NAND2_X1  g643(.A1(new_n662), .A2(new_n217), .ZN(new_n845));
  XOR2_X1   g644(.A(new_n845), .B(KEYINPUT121), .Z(new_n846));
  OAI21_X1  g645(.A(new_n846), .B1(new_n838), .B2(new_n839), .ZN(new_n847));
  INV_X1    g646(.A(new_n662), .ZN(new_n848));
  OAI21_X1  g647(.A(G120gat), .B1(new_n842), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(G1341gat));
  NAND4_X1  g649(.A1(new_n837), .A2(new_n207), .A3(new_n208), .A4(new_n612), .ZN(new_n851));
  OAI22_X1  g650(.A1(new_n842), .A2(new_n613), .B1(new_n213), .B2(new_n212), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(G1342gat));
  NAND3_X1  g652(.A1(new_n837), .A2(new_n204), .A3(new_n637), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n854), .A2(KEYINPUT56), .ZN(new_n855));
  OAI21_X1  g654(.A(G134gat), .B1(new_n842), .B2(new_n636), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(KEYINPUT56), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(G1343gat));
  NOR3_X1   g657(.A1(new_n760), .A2(new_n472), .A3(new_n669), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n726), .B1(new_n829), .B2(new_n830), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(KEYINPUT57), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n829), .A2(new_n830), .ZN(new_n862));
  AOI21_X1  g661(.A(KEYINPUT57), .B1(new_n862), .B2(new_n806), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI211_X1 g664(.A(KEYINPUT122), .B(KEYINPUT57), .C1(new_n862), .C2(new_n806), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n583), .B(new_n859), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(G141gat), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT123), .ZN(new_n869));
  AND4_X1   g668(.A1(new_n470), .A2(new_n831), .A3(new_n806), .A4(new_n523), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n698), .A2(G141gat), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT58), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT58), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n868), .A2(new_n875), .A3(new_n872), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(G1344gat));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n859), .B1(new_n865), .B2(new_n866), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n878), .B(G148gat), .C1(new_n879), .C2(new_n848), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n860), .A2(KEYINPUT57), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n862), .A2(KEYINPUT57), .A3(new_n806), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n859), .A2(new_n662), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n385), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n880), .B1(new_n878), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n870), .A2(new_n385), .A3(new_n662), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1345gat));
  OAI21_X1  g687(.A(G155gat), .B1(new_n879), .B2(new_n613), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n870), .A2(new_n381), .A3(new_n612), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(G1346gat));
  OAI21_X1  g690(.A(G162gat), .B1(new_n879), .B2(new_n636), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n870), .A2(new_n382), .A3(new_n637), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(G1347gat));
  AOI21_X1  g693(.A(new_n665), .B1(new_n829), .B2(new_n830), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n895), .A2(new_n669), .A3(new_n832), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n896), .A2(new_n583), .A3(new_n267), .A4(new_n268), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n665), .A2(new_n470), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n841), .A2(new_n762), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(G169gat), .B1(new_n899), .B2(new_n698), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  XOR2_X1   g700(.A(new_n901), .B(KEYINPUT124), .Z(G1348gat));
  NAND3_X1  g701(.A1(new_n896), .A2(new_n241), .A3(new_n662), .ZN(new_n903));
  OAI21_X1  g702(.A(G176gat), .B1(new_n899), .B2(new_n848), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1349gat));
  NAND3_X1  g704(.A1(new_n896), .A2(new_n232), .A3(new_n612), .ZN(new_n906));
  OAI21_X1  g705(.A(G183gat), .B1(new_n899), .B2(new_n613), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g708(.A(G190gat), .B1(new_n899), .B2(new_n636), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(KEYINPUT61), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n896), .A2(new_n233), .A3(new_n637), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1351gat));
  NOR3_X1   g712(.A1(new_n760), .A2(new_n470), .A3(new_n499), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n895), .A2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(G197gat), .B1(new_n916), .B2(new_n583), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT125), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n883), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n881), .A2(KEYINPUT125), .A3(new_n882), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n898), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n760), .A2(new_n922), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n923), .A2(G197gat), .A3(new_n583), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n917), .B1(new_n921), .B2(new_n924), .ZN(G1352gat));
  NAND4_X1  g724(.A1(new_n919), .A2(new_n662), .A3(new_n920), .A4(new_n923), .ZN(new_n926));
  XNOR2_X1  g725(.A(KEYINPUT126), .B(G204gat), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n915), .A2(new_n848), .A3(new_n927), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT62), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1353gat));
  NAND3_X1  g730(.A1(new_n883), .A2(new_n612), .A3(new_n923), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(G211gat), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT63), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n932), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n935), .A2(KEYINPUT127), .A3(new_n936), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n915), .A2(G211gat), .A3(new_n613), .ZN(new_n938));
  AOI21_X1  g737(.A(KEYINPUT63), .B1(new_n932), .B2(G211gat), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n937), .A2(new_n941), .ZN(G1354gat));
  AOI21_X1  g741(.A(G218gat), .B1(new_n916), .B2(new_n637), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n923), .A2(G218gat), .A3(new_n637), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n943), .B1(new_n921), .B2(new_n944), .ZN(G1355gat));
endmodule


