//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 1 1 1 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n795, new_n796, new_n797, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n864, new_n865, new_n866, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904;
  INV_X1    g000(.A(G50gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  INV_X1    g002(.A(G211gat), .ZN(new_n204));
  INV_X1    g003(.A(G218gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(KEYINPUT22), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  XOR2_X1   g008(.A(new_n209), .B(KEYINPUT75), .Z(new_n210));
  OR3_X1    g009(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212));
  INV_X1    g011(.A(G148gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G141gat), .ZN(new_n214));
  INV_X1    g013(.A(G141gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G148gat), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n211), .A2(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n215), .A2(G148gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n213), .A2(G141gat), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT79), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT79), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n214), .A2(new_n216), .A3(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n220), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(G155gat), .B(G162gat), .Z(new_n225));
  AOI21_X1  g024(.A(new_n217), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  XOR2_X1   g025(.A(KEYINPUT80), .B(KEYINPUT3), .Z(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT81), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT29), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n210), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n209), .A2(KEYINPUT29), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(KEYINPUT3), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n234), .A2(new_n226), .ZN(new_n235));
  OAI211_X1 g034(.A(G228gat), .B(G233gat), .C1(new_n232), .C2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G228gat), .A2(G233gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n224), .A2(new_n225), .ZN(new_n238));
  INV_X1    g037(.A(new_n217), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(new_n233), .B2(new_n227), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n230), .A2(new_n231), .ZN(new_n242));
  INV_X1    g041(.A(new_n209), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n237), .B(new_n241), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n202), .B1(new_n236), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n236), .A2(new_n244), .A3(new_n202), .ZN(new_n247));
  XOR2_X1   g046(.A(G78gat), .B(G106gat), .Z(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(G22gat), .ZN(new_n249));
  XOR2_X1   g048(.A(KEYINPUT85), .B(KEYINPUT31), .Z(new_n250));
  XOR2_X1   g049(.A(new_n249), .B(new_n250), .Z(new_n251));
  NAND3_X1  g050(.A1(new_n246), .A2(new_n247), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n251), .ZN(new_n253));
  INV_X1    g052(.A(new_n247), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n253), .B1(new_n254), .B2(new_n245), .ZN(new_n255));
  AND2_X1   g054(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  AND2_X1   g055(.A1(KEYINPUT71), .A2(G134gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(G113gat), .B(G120gat), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n257), .B1(new_n258), .B2(KEYINPUT1), .ZN(new_n259));
  INV_X1    g058(.A(G127gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n261));
  INV_X1    g060(.A(G134gat), .ZN(new_n262));
  INV_X1    g061(.A(G113gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n263), .A2(G120gat), .ZN(new_n264));
  INV_X1    g063(.A(G120gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n265), .A2(G113gat), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n261), .B(new_n262), .C1(new_n264), .C2(new_n266), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n259), .A2(new_n260), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n260), .B1(new_n259), .B2(new_n267), .ZN(new_n269));
  OR2_X1    g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n271));
  NAND3_X1  g070(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT67), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(G183gat), .A2(G190gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT24), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g076(.A1(KEYINPUT67), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n278));
  INV_X1    g077(.A(G183gat), .ZN(new_n279));
  INV_X1    g078(.A(G190gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AND4_X1   g080(.A1(new_n274), .A2(new_n277), .A3(new_n278), .A4(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT68), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT25), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G169gat), .ZN(new_n285));
  INV_X1    g084(.A(G176gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n286), .A3(KEYINPUT23), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT23), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n288), .B1(G169gat), .B2(G176gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n274), .A2(new_n277), .A3(new_n278), .A4(new_n281), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n292), .B1(new_n293), .B2(KEYINPUT68), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n271), .B1(new_n284), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n291), .B1(new_n282), .B2(new_n283), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT25), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n297), .B1(new_n293), .B2(KEYINPUT68), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n296), .A2(KEYINPUT69), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n300), .A2(KEYINPUT65), .B1(new_n279), .B2(new_n280), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT65), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n277), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n301), .A2(new_n272), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT66), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n301), .A2(new_n303), .A3(KEYINPUT66), .A4(new_n272), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n306), .A2(new_n292), .A3(new_n307), .ZN(new_n308));
  AOI22_X1  g107(.A1(new_n295), .A2(new_n299), .B1(new_n297), .B2(new_n308), .ZN(new_n309));
  AND2_X1   g108(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n280), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT28), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT27), .B(G183gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n315), .A2(KEYINPUT28), .A3(new_n280), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n314), .A2(new_n316), .B1(G183gat), .B2(G190gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT70), .ZN(new_n318));
  OR3_X1    g117(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(new_n290), .A3(new_n320), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n317), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n318), .B1(new_n317), .B2(new_n321), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n270), .B1(new_n309), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n297), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n284), .A2(new_n294), .A3(new_n271), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT69), .B1(new_n296), .B2(new_n298), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n268), .A2(new_n269), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n317), .A2(new_n321), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT70), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n317), .A2(new_n318), .A3(new_n321), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n329), .A2(new_n330), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G227gat), .A2(G233gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n336), .B(KEYINPUT64), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n325), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT72), .B(KEYINPUT33), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT73), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G15gat), .B(G43gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(G71gat), .ZN(new_n343));
  XOR2_X1   g142(.A(new_n343), .B(G99gat), .Z(new_n344));
  NAND2_X1  g143(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n339), .A2(KEYINPUT32), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(new_n341), .A3(new_n344), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n325), .A2(new_n335), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n336), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT34), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT34), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n350), .A2(new_n353), .A3(new_n337), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n348), .A2(new_n349), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n355), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n346), .A2(new_n341), .A3(new_n344), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n346), .B1(new_n341), .B2(new_n344), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n256), .A2(new_n357), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(G225gat), .A2(G233gat), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n226), .B1(new_n268), .B2(new_n269), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NOR3_X1   g167(.A1(new_n226), .A2(new_n268), .A3(new_n269), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n366), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT82), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI211_X1 g171(.A(KEYINPUT82), .B(new_n366), .C1(new_n368), .C2(new_n369), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(KEYINPUT5), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT83), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n240), .A2(KEYINPUT3), .ZN(new_n377));
  AND2_X1   g176(.A1(new_n229), .A2(KEYINPUT81), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n229), .A2(KEYINPUT81), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n330), .B(new_n377), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n367), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n270), .A2(KEYINPUT4), .A3(new_n226), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n380), .A2(new_n382), .A3(new_n383), .A4(new_n365), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n372), .A2(KEYINPUT83), .A3(KEYINPUT5), .A4(new_n373), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n376), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G1gat), .B(G29gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(G85gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(KEYINPUT0), .B(G57gat), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n388), .B(new_n389), .Z(new_n390));
  AND3_X1   g189(.A1(new_n383), .A2(KEYINPUT84), .A3(new_n382), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT84), .B1(new_n383), .B2(new_n382), .ZN(new_n392));
  OR2_X1    g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT5), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n393), .A2(new_n394), .A3(new_n365), .A4(new_n380), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n386), .A2(new_n390), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT6), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n390), .B1(new_n386), .B2(new_n395), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n210), .ZN(new_n401));
  AND2_X1   g200(.A1(G226gat), .A2(G233gat), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n329), .A2(new_n402), .A3(new_n331), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT76), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n405), .B1(new_n309), .B2(new_n324), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n329), .A2(KEYINPUT76), .A3(new_n334), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n402), .A2(KEYINPUT29), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n404), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n406), .A2(new_n407), .A3(new_n402), .ZN(new_n411));
  INV_X1    g210(.A(new_n331), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n409), .B1(new_n309), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n401), .A2(new_n410), .B1(new_n414), .B2(new_n243), .ZN(new_n415));
  XNOR2_X1  g214(.A(G8gat), .B(G36gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(G64gat), .B(G92gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  XOR2_X1   g217(.A(new_n418), .B(KEYINPUT77), .Z(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT78), .B1(new_n415), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n414), .A2(new_n243), .ZN(new_n422));
  NOR3_X1   g221(.A1(new_n309), .A2(new_n324), .A3(new_n405), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT76), .B1(new_n329), .B2(new_n334), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n409), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n425), .A2(new_n401), .A3(new_n403), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT78), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n428), .A3(new_n419), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n421), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n418), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT30), .B1(new_n415), .B2(new_n431), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n422), .A2(new_n426), .A3(KEYINPUT30), .A4(new_n431), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n400), .A2(new_n430), .A3(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT35), .B1(new_n364), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n256), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n428), .B1(new_n427), .B2(new_n419), .ZN(new_n439));
  AOI211_X1 g238(.A(KEYINPUT78), .B(new_n420), .C1(new_n422), .C2(new_n426), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT86), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n422), .A2(new_n426), .A3(new_n431), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT30), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n433), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n441), .A2(new_n442), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT86), .B1(new_n435), .B2(new_n430), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n438), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT91), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n386), .A2(new_n395), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n390), .B(KEYINPUT87), .Z(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n454), .A2(new_n397), .A3(new_n396), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n399), .A2(KEYINPUT6), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT35), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT74), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n361), .A2(new_n458), .A3(new_n356), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n348), .A2(KEYINPUT74), .A3(new_n349), .A4(new_n355), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NOR3_X1   g261(.A1(new_n449), .A2(new_n450), .A3(new_n462), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n457), .A2(new_n461), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n442), .B1(new_n441), .B2(new_n446), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n435), .A2(KEYINPUT86), .A3(new_n430), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n256), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT91), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n437), .B1(new_n463), .B2(new_n468), .ZN(new_n469));
  NOR3_X1   g268(.A1(new_n368), .A2(new_n369), .A3(new_n366), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT88), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT88), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n380), .B1(new_n391), .B2(new_n392), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n472), .B1(new_n473), .B2(new_n366), .ZN(new_n474));
  OAI211_X1 g273(.A(KEYINPUT39), .B(new_n471), .C1(new_n474), .C2(new_n470), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT39), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n473), .A2(new_n476), .A3(new_n366), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n452), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT89), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT40), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n481), .A2(new_n454), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n478), .A2(new_n479), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT40), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n482), .A2(new_n465), .A3(new_n466), .A4(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(KEYINPUT90), .B(KEYINPUT37), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n415), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n410), .A2(new_n401), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n414), .A2(new_n243), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT37), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n487), .A2(new_n490), .A3(new_n419), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT38), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n492), .A3(new_n443), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n431), .B1(new_n427), .B2(KEYINPUT37), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n494), .A2(KEYINPUT38), .A3(new_n487), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n496), .A2(new_n456), .A3(new_n455), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n485), .A2(new_n438), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n436), .A2(new_n256), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n362), .A2(new_n357), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT36), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n502), .B1(new_n461), .B2(new_n501), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n498), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n469), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(G29gat), .ZN(new_n506));
  INV_X1    g305(.A(G36gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(KEYINPUT14), .ZN(new_n509));
  XNOR2_X1  g308(.A(G43gat), .B(G50gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT15), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n511), .A2(KEYINPUT92), .ZN(new_n512));
  OAI221_X1 g311(.A(new_n509), .B1(new_n506), .B2(new_n507), .C1(new_n512), .C2(KEYINPUT93), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT92), .B1(G29gat), .B2(G36gat), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n514), .B1(new_n509), .B2(KEYINPUT93), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n511), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n513), .B(new_n516), .C1(KEYINPUT15), .C2(new_n510), .ZN(new_n517));
  XOR2_X1   g316(.A(new_n517), .B(KEYINPUT94), .Z(new_n518));
  XNOR2_X1  g317(.A(G15gat), .B(G22gat), .ZN(new_n519));
  INV_X1    g318(.A(G1gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(KEYINPUT16), .A3(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(new_n520), .B2(new_n519), .ZN(new_n522));
  INV_X1    g321(.A(G8gat), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n522), .B1(KEYINPUT95), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(KEYINPUT95), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n518), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n526), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n517), .A2(KEYINPUT17), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT17), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n529), .B1(new_n518), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n527), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G229gat), .A2(G233gat), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OR3_X1    g333(.A1(new_n534), .A2(KEYINPUT96), .A3(KEYINPUT18), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n534), .B1(KEYINPUT96), .B2(KEYINPUT18), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n518), .B(new_n526), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n533), .B(KEYINPUT13), .Z(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n535), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G113gat), .B(G141gat), .ZN(new_n541));
  INV_X1    g340(.A(G197gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(KEYINPUT11), .B(G169gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT12), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n540), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n540), .A2(new_n547), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G120gat), .B(G148gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(G176gat), .B(G204gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT97), .ZN(new_n556));
  XNOR2_X1  g355(.A(G71gat), .B(G78gat), .ZN(new_n557));
  INV_X1    g356(.A(G57gat), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n558), .A2(G64gat), .ZN(new_n559));
  INV_X1    g358(.A(G64gat), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n560), .A2(G57gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT98), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT98), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n563), .B1(new_n560), .B2(G57gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n556), .B(new_n557), .C1(new_n559), .C2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT99), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n556), .B1(new_n561), .B2(new_n559), .ZN(new_n569));
  INV_X1    g368(.A(new_n557), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n566), .A2(new_n567), .ZN(new_n572));
  NOR3_X1   g371(.A1(new_n568), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT102), .B(G85gat), .ZN(new_n574));
  INV_X1    g373(.A(G92gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(G99gat), .A2(G106gat), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n574), .A2(new_n575), .B1(KEYINPUT8), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G85gat), .A2(G92gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT7), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT100), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT101), .ZN(new_n581));
  OR3_X1    g380(.A1(new_n578), .A2(new_n581), .A3(KEYINPUT7), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n581), .B1(new_n578), .B2(KEYINPUT7), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n577), .B1(new_n580), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G99gat), .B(G106gat), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n585), .B(new_n586), .Z(new_n587));
  XNOR2_X1  g386(.A(new_n573), .B(new_n587), .ZN(new_n588));
  AND2_X1   g387(.A1(G230gat), .A2(G233gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n587), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n591), .A2(KEYINPUT10), .A3(new_n573), .ZN(new_n592));
  INV_X1    g391(.A(new_n588), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n592), .B1(new_n593), .B2(KEYINPUT10), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n594), .A2(new_n590), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n595), .A2(KEYINPUT106), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n594), .A2(KEYINPUT106), .A3(new_n590), .ZN(new_n597));
  OAI221_X1 g396(.A(new_n554), .B1(new_n588), .B2(new_n590), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n588), .A2(new_n590), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n553), .B1(new_n595), .B2(new_n599), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n550), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n526), .B1(KEYINPUT21), .B2(new_n573), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(new_n279), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n573), .A2(KEYINPUT21), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G127gat), .B(G155gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(G211gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n609), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G232gat), .A2(G233gat), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT41), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n619), .B1(new_n518), .B2(new_n591), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n620), .B(KEYINPUT103), .Z(new_n621));
  NAND2_X1  g420(.A1(new_n531), .A2(new_n587), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT104), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n625), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n621), .A2(new_n627), .A3(new_n622), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G134gat), .B(G162gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n617), .A2(new_n618), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n629), .A2(KEYINPUT105), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(KEYINPUT105), .ZN(new_n634));
  OAI211_X1 g433(.A(new_n634), .B(new_n628), .C1(new_n626), .C2(new_n632), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n505), .A2(new_n603), .A3(new_n616), .A4(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(new_n400), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(new_n520), .ZN(G1324gat));
  NOR2_X1   g439(.A1(new_n447), .A2(new_n448), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n643), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n644), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n645), .B(KEYINPUT42), .Z(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(new_n523), .B2(new_n643), .ZN(G1325gat));
  INV_X1    g446(.A(G15gat), .ZN(new_n648));
  INV_X1    g447(.A(new_n461), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n648), .B1(new_n638), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT107), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n638), .A2(new_n648), .A3(new_n503), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(G1326gat));
  NOR2_X1   g452(.A1(new_n638), .A2(new_n438), .ZN(new_n654));
  XOR2_X1   g453(.A(KEYINPUT43), .B(G22gat), .Z(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(G1327gat));
  NOR2_X1   g455(.A1(new_n637), .A2(KEYINPUT44), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n469), .A2(KEYINPUT108), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT108), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n659), .B(new_n437), .C1(new_n463), .C2(new_n468), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT109), .B1(new_n661), .B2(new_n504), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT109), .ZN(new_n663));
  INV_X1    g462(.A(new_n504), .ZN(new_n664));
  AOI211_X1 g463(.A(new_n663), .B(new_n664), .C1(new_n658), .C2(new_n660), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n657), .B1(new_n662), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(KEYINPUT110), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n637), .B1(new_n469), .B2(new_n504), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n669));
  OR2_X1    g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT110), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n671), .B(new_n657), .C1(new_n662), .C2(new_n665), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n667), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n400), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n616), .A2(new_n602), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n676), .A2(KEYINPUT111), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(KEYINPUT111), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n677), .A2(G29gat), .A3(new_n678), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n675), .A2(new_n668), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n680), .A2(new_n506), .A3(new_n674), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT45), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n679), .A2(new_n682), .ZN(G1328gat));
  NAND3_X1  g482(.A1(new_n680), .A2(new_n507), .A3(new_n641), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT112), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT113), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n685), .B1(new_n686), .B2(KEYINPUT46), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(KEYINPUT46), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n687), .B(new_n688), .Z(new_n689));
  AND3_X1   g488(.A1(new_n673), .A2(new_n641), .A3(new_n675), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n689), .B1(new_n507), .B2(new_n690), .ZN(G1329gat));
  INV_X1    g490(.A(new_n503), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n673), .A2(new_n692), .A3(new_n675), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(G43gat), .ZN(new_n694));
  INV_X1    g493(.A(new_n680), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n695), .A2(G43gat), .A3(new_n649), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT114), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT47), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n696), .B1(new_n693), .B2(G43gat), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT47), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n701), .A2(KEYINPUT114), .A3(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n700), .A2(new_n703), .ZN(G1330gat));
  NAND4_X1  g503(.A1(new_n673), .A2(G50gat), .A3(new_n256), .A4(new_n675), .ZN(new_n705));
  NAND2_X1  g504(.A1(KEYINPUT115), .A2(KEYINPUT48), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n202), .B1(new_n695), .B2(new_n438), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(KEYINPUT115), .A2(KEYINPUT48), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n708), .B(new_n709), .Z(G1331gat));
  INV_X1    g509(.A(new_n601), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n614), .A2(new_n615), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n712), .A2(new_n550), .A3(new_n636), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n711), .B(new_n713), .C1(new_n662), .C2(new_n665), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n714), .A2(new_n400), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(new_n558), .ZN(G1332gat));
  NOR2_X1   g515(.A1(new_n714), .A2(new_n642), .ZN(new_n717));
  NOR2_X1   g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  AND2_X1   g517(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n720), .B1(new_n717), .B2(new_n718), .ZN(G1333gat));
  OR3_X1    g520(.A1(new_n714), .A2(G71gat), .A3(new_n649), .ZN(new_n722));
  OAI21_X1  g521(.A(G71gat), .B1(new_n714), .B2(new_n503), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XOR2_X1   g523(.A(new_n724), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g524(.A1(new_n714), .A2(new_n438), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT116), .B(G78gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1335gat));
  NOR2_X1   g527(.A1(new_n616), .A2(new_n550), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n673), .A2(new_n711), .A3(new_n729), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n730), .A2(new_n400), .A3(new_n574), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n661), .A2(new_n504), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n732), .A2(new_n636), .A3(new_n729), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n733), .A2(KEYINPUT51), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(KEYINPUT51), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n736), .A2(new_n674), .A3(new_n711), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n731), .B1(new_n574), .B2(new_n737), .ZN(G1336gat));
  NAND4_X1  g537(.A1(new_n734), .A2(new_n711), .A3(new_n641), .A4(new_n735), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n575), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n641), .A2(G92gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n730), .B2(new_n741), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n742), .B(KEYINPUT52), .Z(G1337gat));
  OAI21_X1  g542(.A(G99gat), .B1(new_n730), .B2(new_n503), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n736), .A2(new_n711), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n649), .A2(G99gat), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(G1338gat));
  OAI21_X1  g546(.A(G106gat), .B1(new_n730), .B2(new_n438), .ZN(new_n748));
  INV_X1    g547(.A(G106gat), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n736), .A2(new_n749), .A3(new_n711), .A4(new_n256), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n748), .A2(new_n752), .A3(new_n750), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(G1339gat));
  OAI221_X1 g555(.A(KEYINPUT54), .B1(new_n590), .B2(new_n594), .C1(new_n596), .C2(new_n597), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT54), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n554), .B1(new_n595), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT55), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n757), .A2(KEYINPUT55), .A3(new_n759), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n762), .A2(new_n598), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT118), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n762), .A2(KEYINPUT118), .A3(new_n598), .A4(new_n763), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n766), .A2(new_n550), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n532), .A2(new_n533), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n537), .A2(new_n538), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n545), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n548), .A2(new_n711), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n636), .B1(new_n768), .B2(new_n772), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n548), .A2(new_n636), .A3(new_n771), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n774), .A2(new_n766), .A3(new_n767), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n712), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n713), .A2(new_n601), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT119), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT119), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n776), .A2(new_n780), .A3(new_n777), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n779), .A2(new_n674), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n467), .ZN(new_n783));
  INV_X1    g582(.A(new_n500), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT120), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT120), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n782), .A2(new_n786), .A3(new_n500), .A4(new_n467), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n785), .A2(new_n787), .A3(new_n263), .A4(new_n550), .ZN(new_n788));
  INV_X1    g587(.A(new_n550), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n783), .A2(new_n789), .A3(new_n649), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n788), .B1(new_n263), .B2(new_n790), .ZN(G1340gat));
  NAND4_X1  g590(.A1(new_n785), .A2(new_n787), .A3(new_n265), .A4(new_n711), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n783), .A2(new_n601), .A3(new_n649), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n792), .B1(new_n265), .B2(new_n793), .ZN(G1341gat));
  NOR2_X1   g593(.A1(new_n783), .A2(new_n649), .ZN(new_n795));
  XOR2_X1   g594(.A(KEYINPUT71), .B(G127gat), .Z(new_n796));
  NOR2_X1   g595(.A1(new_n712), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n782), .A2(new_n500), .A3(new_n467), .A4(new_n616), .ZN(new_n798));
  AOI22_X1  g597(.A1(new_n795), .A2(new_n797), .B1(new_n796), .B2(new_n798), .ZN(G1342gat));
  NAND4_X1  g598(.A1(new_n782), .A2(new_n262), .A3(new_n500), .A4(new_n467), .ZN(new_n800));
  OR3_X1    g599(.A1(new_n800), .A2(KEYINPUT56), .A3(new_n637), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT56), .B1(new_n800), .B2(new_n637), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n783), .A2(new_n649), .A3(new_n637), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n801), .B(new_n802), .C1(new_n262), .C2(new_n803), .ZN(G1343gat));
  NAND3_X1  g603(.A1(new_n779), .A2(new_n256), .A3(new_n781), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n692), .A2(new_n400), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  OR3_X1    g606(.A1(new_n805), .A2(KEYINPUT121), .A3(new_n807), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n789), .A2(G141gat), .A3(new_n641), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT121), .B1(new_n805), .B2(new_n807), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n807), .A2(new_n641), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n772), .B1(new_n789), .B2(new_n764), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n775), .B1(new_n637), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n777), .B1(new_n815), .B2(new_n616), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n256), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n813), .B1(new_n817), .B2(KEYINPUT57), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n779), .A2(new_n819), .A3(new_n256), .A4(new_n781), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n818), .A2(new_n820), .A3(new_n550), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(G141gat), .ZN(new_n822));
  XOR2_X1   g621(.A(KEYINPUT122), .B(KEYINPUT58), .Z(new_n823));
  NAND3_X1  g622(.A1(new_n811), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT58), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n805), .A2(new_n807), .ZN(new_n826));
  AOI22_X1  g625(.A1(new_n821), .A2(G141gat), .B1(new_n826), .B2(new_n809), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n824), .B1(new_n825), .B2(new_n827), .ZN(G1344gat));
  NOR2_X1   g627(.A1(new_n601), .A2(G148gat), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n808), .A2(new_n642), .A3(new_n810), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n818), .A2(new_n820), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(new_n601), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n832), .A2(KEYINPUT59), .A3(new_n213), .ZN(new_n833));
  XOR2_X1   g632(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n834));
  NAND2_X1  g633(.A1(new_n805), .A2(KEYINPUT57), .ZN(new_n835));
  INV_X1    g634(.A(new_n777), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n814), .A2(new_n637), .ZN(new_n837));
  INV_X1    g636(.A(new_n764), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n774), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n616), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n819), .B(new_n256), .C1(new_n836), .C2(new_n840), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n835), .A2(new_n711), .A3(new_n812), .A4(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n834), .B1(new_n842), .B2(G148gat), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n830), .B1(new_n833), .B2(new_n843), .ZN(G1345gat));
  INV_X1    g643(.A(G155gat), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n831), .A2(new_n845), .A3(new_n712), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n808), .A2(new_n642), .A3(new_n810), .A4(new_n616), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n847), .B2(new_n845), .ZN(G1346gat));
  NOR2_X1   g647(.A1(new_n637), .A2(G162gat), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n808), .A2(new_n642), .A3(new_n810), .A4(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(G162gat), .B1(new_n831), .B2(new_n637), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(G1347gat));
  NOR2_X1   g651(.A1(new_n642), .A2(new_n674), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n649), .A2(new_n256), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n779), .A2(new_n781), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(G169gat), .B1(new_n855), .B2(new_n789), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT124), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n779), .A2(new_n781), .A3(new_n853), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n363), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n859), .A2(G169gat), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n857), .B1(new_n860), .B2(new_n550), .ZN(new_n861));
  NOR4_X1   g660(.A1(new_n859), .A2(KEYINPUT124), .A3(G169gat), .A4(new_n789), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n856), .B1(new_n861), .B2(new_n862), .ZN(G1348gat));
  NOR3_X1   g662(.A1(new_n855), .A2(new_n286), .A3(new_n601), .ZN(new_n864));
  INV_X1    g663(.A(new_n859), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n711), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n864), .B1(new_n866), .B2(new_n286), .ZN(G1349gat));
  NAND4_X1  g666(.A1(new_n858), .A2(new_n315), .A3(new_n363), .A4(new_n616), .ZN(new_n868));
  OAI21_X1  g667(.A(G183gat), .B1(new_n855), .B2(new_n712), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g670(.A1(new_n865), .A2(new_n280), .A3(new_n636), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n858), .A2(new_n636), .A3(new_n854), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT61), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n873), .A2(new_n874), .A3(G190gat), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n874), .B1(new_n873), .B2(G190gat), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n872), .B1(new_n876), .B2(new_n877), .ZN(G1351gat));
  AND2_X1   g677(.A1(new_n835), .A2(new_n841), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n853), .A2(new_n503), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n550), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(G197gat), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n779), .A2(new_n256), .A3(new_n781), .A4(new_n880), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(new_n542), .A3(new_n550), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT125), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n882), .A2(new_n886), .ZN(G1352gat));
  NOR3_X1   g686(.A1(new_n883), .A2(G204gat), .A3(new_n601), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT62), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n835), .A2(new_n711), .A3(new_n841), .A4(new_n880), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G204gat), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n889), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT126), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT62), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n894), .B1(new_n888), .B2(new_n895), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n890), .B(new_n892), .C1(new_n893), .C2(new_n896), .ZN(G1353gat));
  NAND3_X1  g696(.A1(new_n884), .A2(new_n204), .A3(new_n616), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n835), .A2(new_n616), .A3(new_n841), .A4(new_n880), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n899), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT63), .B1(new_n899), .B2(G211gat), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(G1354gat));
  NAND3_X1  g701(.A1(new_n884), .A2(new_n205), .A3(new_n636), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n879), .A2(new_n636), .A3(new_n880), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(new_n205), .ZN(G1355gat));
endmodule


