

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U553 ( .A(n539), .B(KEYINPUT65), .ZN(G160) );
  XOR2_X1 U554 ( .A(KEYINPUT17), .B(n520), .Z(n891) );
  NOR2_X1 U555 ( .A1(n738), .A2(n737), .ZN(n727) );
  INV_X1 U556 ( .A(KEYINPUT102), .ZN(n754) );
  NOR2_X1 U557 ( .A1(G651), .A2(n623), .ZN(n652) );
  AND2_X1 U558 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U559 ( .A(G2105), .ZN(n523) );
  INV_X1 U560 ( .A(G2104), .ZN(n527) );
  NOR2_X1 U561 ( .A1(n523), .A2(n527), .ZN(n895) );
  NAND2_X1 U562 ( .A1(G111), .A2(n895), .ZN(n522) );
  NOR2_X1 U563 ( .A1(G2105), .A2(G2104), .ZN(n520) );
  NAND2_X1 U564 ( .A1(G135), .A2(n891), .ZN(n521) );
  NAND2_X1 U565 ( .A1(n522), .A2(n521), .ZN(n526) );
  NOR2_X1 U566 ( .A1(G2104), .A2(n523), .ZN(n896) );
  NAND2_X1 U567 ( .A1(n896), .A2(G123), .ZN(n524) );
  XOR2_X1 U568 ( .A(KEYINPUT18), .B(n524), .Z(n525) );
  NOR2_X1 U569 ( .A1(n526), .A2(n525), .ZN(n530) );
  NOR2_X1 U570 ( .A1(n527), .A2(G2105), .ZN(n528) );
  XNOR2_X1 U571 ( .A(n528), .B(KEYINPUT66), .ZN(n709) );
  BUF_X1 U572 ( .A(n709), .Z(n892) );
  NAND2_X1 U573 ( .A1(G99), .A2(n892), .ZN(n529) );
  NAND2_X1 U574 ( .A1(n530), .A2(n529), .ZN(n923) );
  XNOR2_X1 U575 ( .A(G2096), .B(n923), .ZN(n531) );
  OR2_X1 U576 ( .A1(G2100), .A2(n531), .ZN(G156) );
  INV_X1 U577 ( .A(G57), .ZN(G237) );
  NAND2_X1 U578 ( .A1(n891), .A2(G137), .ZN(n538) );
  NAND2_X1 U579 ( .A1(G113), .A2(n895), .ZN(n533) );
  NAND2_X1 U580 ( .A1(G125), .A2(n896), .ZN(n532) );
  NAND2_X1 U581 ( .A1(n533), .A2(n532), .ZN(n536) );
  NAND2_X1 U582 ( .A1(G101), .A2(n709), .ZN(n534) );
  XNOR2_X1 U583 ( .A(KEYINPUT23), .B(n534), .ZN(n535) );
  NOR2_X1 U584 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U585 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U586 ( .A1(G543), .A2(G651), .ZN(n540) );
  XNOR2_X1 U587 ( .A(n540), .B(KEYINPUT64), .ZN(n642) );
  NAND2_X1 U588 ( .A1(n642), .A2(G89), .ZN(n541) );
  XNOR2_X1 U589 ( .A(n541), .B(KEYINPUT4), .ZN(n542) );
  XNOR2_X1 U590 ( .A(KEYINPUT78), .B(n542), .ZN(n546) );
  INV_X1 U591 ( .A(G651), .ZN(n548) );
  XOR2_X1 U592 ( .A(KEYINPUT0), .B(G543), .Z(n623) );
  OR2_X1 U593 ( .A1(n548), .A2(n623), .ZN(n543) );
  XOR2_X1 U594 ( .A(KEYINPUT68), .B(n543), .Z(n645) );
  NAND2_X1 U595 ( .A1(G76), .A2(n645), .ZN(n544) );
  XOR2_X1 U596 ( .A(KEYINPUT79), .B(n544), .Z(n545) );
  NAND2_X1 U597 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U598 ( .A(KEYINPUT5), .B(n547), .ZN(n555) );
  NOR2_X1 U599 ( .A1(G543), .A2(n548), .ZN(n549) );
  XOR2_X1 U600 ( .A(KEYINPUT1), .B(n549), .Z(n641) );
  NAND2_X1 U601 ( .A1(n641), .A2(G63), .ZN(n550) );
  XNOR2_X1 U602 ( .A(n550), .B(KEYINPUT80), .ZN(n552) );
  NAND2_X1 U603 ( .A1(G51), .A2(n652), .ZN(n551) );
  NAND2_X1 U604 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U605 ( .A(KEYINPUT6), .B(n553), .Z(n554) );
  NAND2_X1 U606 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U607 ( .A(KEYINPUT7), .B(n556), .ZN(G168) );
  XOR2_X1 U608 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U609 ( .A1(G7), .A2(G661), .ZN(n557) );
  XOR2_X1 U610 ( .A(n557), .B(KEYINPUT10), .Z(n921) );
  NAND2_X1 U611 ( .A1(n921), .A2(G567), .ZN(n558) );
  XOR2_X1 U612 ( .A(KEYINPUT11), .B(n558), .Z(G234) );
  XNOR2_X1 U613 ( .A(KEYINPUT13), .B(KEYINPUT75), .ZN(n563) );
  NAND2_X1 U614 ( .A1(G81), .A2(n642), .ZN(n559) );
  XNOR2_X1 U615 ( .A(n559), .B(KEYINPUT12), .ZN(n561) );
  NAND2_X1 U616 ( .A1(G68), .A2(n645), .ZN(n560) );
  NAND2_X1 U617 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U618 ( .A(n563), .B(n562), .ZN(n566) );
  NAND2_X1 U619 ( .A1(n641), .A2(G56), .ZN(n564) );
  XOR2_X1 U620 ( .A(KEYINPUT14), .B(n564), .Z(n565) );
  NOR2_X1 U621 ( .A1(n566), .A2(n565), .ZN(n568) );
  NAND2_X1 U622 ( .A1(n652), .A2(G43), .ZN(n567) );
  NAND2_X1 U623 ( .A1(n568), .A2(n567), .ZN(n1011) );
  INV_X1 U624 ( .A(G860), .ZN(n601) );
  OR2_X1 U625 ( .A1(n1011), .A2(n601), .ZN(G153) );
  XNOR2_X1 U626 ( .A(KEYINPUT9), .B(KEYINPUT72), .ZN(n573) );
  NAND2_X1 U627 ( .A1(G77), .A2(n645), .ZN(n571) );
  NAND2_X1 U628 ( .A1(G90), .A2(n642), .ZN(n569) );
  XOR2_X1 U629 ( .A(KEYINPUT71), .B(n569), .Z(n570) );
  NAND2_X1 U630 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U631 ( .A(n573), .B(n572), .Z(n576) );
  NAND2_X1 U632 ( .A1(n652), .A2(G52), .ZN(n574) );
  XOR2_X1 U633 ( .A(KEYINPUT70), .B(n574), .Z(n575) );
  NOR2_X1 U634 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U635 ( .A1(n641), .A2(G64), .ZN(n577) );
  NAND2_X1 U636 ( .A1(n578), .A2(n577), .ZN(G301) );
  NAND2_X1 U637 ( .A1(n652), .A2(G54), .ZN(n585) );
  NAND2_X1 U638 ( .A1(n641), .A2(G66), .ZN(n580) );
  NAND2_X1 U639 ( .A1(G92), .A2(n642), .ZN(n579) );
  NAND2_X1 U640 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U641 ( .A1(n645), .A2(G79), .ZN(n581) );
  XOR2_X1 U642 ( .A(KEYINPUT76), .B(n581), .Z(n582) );
  NOR2_X1 U643 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U644 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U645 ( .A(KEYINPUT15), .B(n586), .ZN(n995) );
  NOR2_X1 U646 ( .A1(n995), .A2(G868), .ZN(n587) );
  XNOR2_X1 U647 ( .A(n587), .B(KEYINPUT77), .ZN(n589) );
  NAND2_X1 U648 ( .A1(G868), .A2(G301), .ZN(n588) );
  NAND2_X1 U649 ( .A1(n589), .A2(n588), .ZN(G284) );
  NAND2_X1 U650 ( .A1(G53), .A2(n652), .ZN(n596) );
  NAND2_X1 U651 ( .A1(G91), .A2(n642), .ZN(n591) );
  NAND2_X1 U652 ( .A1(G78), .A2(n645), .ZN(n590) );
  NAND2_X1 U653 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U654 ( .A1(G65), .A2(n641), .ZN(n592) );
  XNOR2_X1 U655 ( .A(KEYINPUT73), .B(n592), .ZN(n593) );
  NOR2_X1 U656 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U657 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U658 ( .A(n597), .B(KEYINPUT74), .Z(n922) );
  INV_X1 U659 ( .A(G868), .ZN(n663) );
  NAND2_X1 U660 ( .A1(n922), .A2(n663), .ZN(n598) );
  XNOR2_X1 U661 ( .A(n598), .B(KEYINPUT81), .ZN(n600) );
  NOR2_X1 U662 ( .A1(n663), .A2(G286), .ZN(n599) );
  NOR2_X1 U663 ( .A1(n600), .A2(n599), .ZN(G297) );
  NAND2_X1 U664 ( .A1(n601), .A2(G559), .ZN(n602) );
  NAND2_X1 U665 ( .A1(n602), .A2(n995), .ZN(n603) );
  XNOR2_X1 U666 ( .A(n603), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U667 ( .A1(n995), .A2(G868), .ZN(n604) );
  NOR2_X1 U668 ( .A1(G559), .A2(n604), .ZN(n605) );
  XNOR2_X1 U669 ( .A(n605), .B(KEYINPUT82), .ZN(n607) );
  NOR2_X1 U670 ( .A1(n1011), .A2(G868), .ZN(n606) );
  NOR2_X1 U671 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U672 ( .A(KEYINPUT83), .B(n608), .Z(G282) );
  XNOR2_X1 U673 ( .A(n1011), .B(KEYINPUT84), .ZN(n610) );
  NAND2_X1 U674 ( .A1(n995), .A2(G559), .ZN(n609) );
  XNOR2_X1 U675 ( .A(n610), .B(n609), .ZN(n661) );
  NOR2_X1 U676 ( .A1(G860), .A2(n661), .ZN(n619) );
  NAND2_X1 U677 ( .A1(n641), .A2(G67), .ZN(n611) );
  XOR2_X1 U678 ( .A(KEYINPUT85), .B(n611), .Z(n613) );
  NAND2_X1 U679 ( .A1(n652), .A2(G55), .ZN(n612) );
  NAND2_X1 U680 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U681 ( .A(KEYINPUT86), .B(n614), .ZN(n618) );
  NAND2_X1 U682 ( .A1(G93), .A2(n642), .ZN(n616) );
  NAND2_X1 U683 ( .A1(G80), .A2(n645), .ZN(n615) );
  NAND2_X1 U684 ( .A1(n616), .A2(n615), .ZN(n617) );
  OR2_X1 U685 ( .A1(n618), .A2(n617), .ZN(n664) );
  XOR2_X1 U686 ( .A(n619), .B(n664), .Z(G145) );
  NAND2_X1 U687 ( .A1(G49), .A2(n652), .ZN(n621) );
  NAND2_X1 U688 ( .A1(G74), .A2(G651), .ZN(n620) );
  NAND2_X1 U689 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U690 ( .A1(n641), .A2(n622), .ZN(n625) );
  NAND2_X1 U691 ( .A1(n623), .A2(G87), .ZN(n624) );
  NAND2_X1 U692 ( .A1(n625), .A2(n624), .ZN(G288) );
  NAND2_X1 U693 ( .A1(n641), .A2(G62), .ZN(n627) );
  NAND2_X1 U694 ( .A1(G75), .A2(n645), .ZN(n626) );
  NAND2_X1 U695 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U696 ( .A1(G88), .A2(n642), .ZN(n628) );
  XNOR2_X1 U697 ( .A(KEYINPUT91), .B(n628), .ZN(n629) );
  NOR2_X1 U698 ( .A1(n630), .A2(n629), .ZN(n632) );
  NAND2_X1 U699 ( .A1(n652), .A2(G50), .ZN(n631) );
  NAND2_X1 U700 ( .A1(n632), .A2(n631), .ZN(G303) );
  INV_X1 U701 ( .A(G303), .ZN(G166) );
  NAND2_X1 U702 ( .A1(G85), .A2(n642), .ZN(n633) );
  XOR2_X1 U703 ( .A(KEYINPUT67), .B(n633), .Z(n635) );
  NAND2_X1 U704 ( .A1(G72), .A2(n645), .ZN(n634) );
  NAND2_X1 U705 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U706 ( .A(KEYINPUT69), .B(n636), .ZN(n640) );
  NAND2_X1 U707 ( .A1(G60), .A2(n641), .ZN(n638) );
  NAND2_X1 U708 ( .A1(G47), .A2(n652), .ZN(n637) );
  AND2_X1 U709 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U710 ( .A1(n640), .A2(n639), .ZN(G290) );
  NAND2_X1 U711 ( .A1(n641), .A2(G61), .ZN(n644) );
  NAND2_X1 U712 ( .A1(G86), .A2(n642), .ZN(n643) );
  NAND2_X1 U713 ( .A1(n644), .A2(n643), .ZN(n650) );
  XOR2_X1 U714 ( .A(KEYINPUT88), .B(KEYINPUT2), .Z(n647) );
  NAND2_X1 U715 ( .A1(G73), .A2(n645), .ZN(n646) );
  XNOR2_X1 U716 ( .A(n647), .B(n646), .ZN(n648) );
  XOR2_X1 U717 ( .A(KEYINPUT87), .B(n648), .Z(n649) );
  NOR2_X1 U718 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U719 ( .A(KEYINPUT89), .B(n651), .Z(n654) );
  NAND2_X1 U720 ( .A1(n652), .A2(G48), .ZN(n653) );
  NAND2_X1 U721 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U722 ( .A(KEYINPUT90), .B(n655), .ZN(G305) );
  XNOR2_X1 U723 ( .A(G288), .B(KEYINPUT19), .ZN(n657) );
  XOR2_X1 U724 ( .A(n922), .B(G166), .Z(n656) );
  XNOR2_X1 U725 ( .A(n657), .B(n656), .ZN(n658) );
  XOR2_X1 U726 ( .A(n664), .B(n658), .Z(n660) );
  XNOR2_X1 U727 ( .A(G290), .B(G305), .ZN(n659) );
  XNOR2_X1 U728 ( .A(n660), .B(n659), .ZN(n910) );
  XOR2_X1 U729 ( .A(n910), .B(n661), .Z(n662) );
  NOR2_X1 U730 ( .A1(n663), .A2(n662), .ZN(n666) );
  NOR2_X1 U731 ( .A1(G868), .A2(n664), .ZN(n665) );
  NOR2_X1 U732 ( .A1(n666), .A2(n665), .ZN(G295) );
  NAND2_X1 U733 ( .A1(G2084), .A2(G2078), .ZN(n668) );
  XOR2_X1 U734 ( .A(KEYINPUT20), .B(KEYINPUT92), .Z(n667) );
  XNOR2_X1 U735 ( .A(n668), .B(n667), .ZN(n669) );
  NAND2_X1 U736 ( .A1(G2090), .A2(n669), .ZN(n670) );
  XNOR2_X1 U737 ( .A(KEYINPUT21), .B(n670), .ZN(n671) );
  NAND2_X1 U738 ( .A1(n671), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U739 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U740 ( .A(KEYINPUT22), .B(KEYINPUT93), .Z(n673) );
  NAND2_X1 U741 ( .A1(G132), .A2(G82), .ZN(n672) );
  XNOR2_X1 U742 ( .A(n673), .B(n672), .ZN(n674) );
  NOR2_X1 U743 ( .A1(n674), .A2(G218), .ZN(n675) );
  NAND2_X1 U744 ( .A1(G96), .A2(n675), .ZN(n832) );
  NAND2_X1 U745 ( .A1(n832), .A2(G2106), .ZN(n679) );
  NAND2_X1 U746 ( .A1(G69), .A2(G120), .ZN(n676) );
  NOR2_X1 U747 ( .A1(G237), .A2(n676), .ZN(n677) );
  NAND2_X1 U748 ( .A1(G108), .A2(n677), .ZN(n833) );
  NAND2_X1 U749 ( .A1(n833), .A2(G567), .ZN(n678) );
  NAND2_X1 U750 ( .A1(n679), .A2(n678), .ZN(n920) );
  NAND2_X1 U751 ( .A1(G661), .A2(G483), .ZN(n680) );
  NOR2_X1 U752 ( .A1(n920), .A2(n680), .ZN(n831) );
  NAND2_X1 U753 ( .A1(n831), .A2(G36), .ZN(G176) );
  NAND2_X1 U754 ( .A1(G114), .A2(n895), .ZN(n682) );
  NAND2_X1 U755 ( .A1(G126), .A2(n896), .ZN(n681) );
  NAND2_X1 U756 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U757 ( .A(KEYINPUT94), .B(n683), .Z(n685) );
  NAND2_X1 U758 ( .A1(n891), .A2(G138), .ZN(n684) );
  NAND2_X1 U759 ( .A1(n685), .A2(n684), .ZN(n688) );
  NAND2_X1 U760 ( .A1(G102), .A2(n709), .ZN(n686) );
  XNOR2_X1 U761 ( .A(KEYINPUT95), .B(n686), .ZN(n687) );
  NOR2_X1 U762 ( .A1(n688), .A2(n687), .ZN(G164) );
  NAND2_X1 U763 ( .A1(G160), .A2(G40), .ZN(n689) );
  XNOR2_X1 U764 ( .A(n689), .B(KEYINPUT96), .ZN(n718) );
  NOR2_X1 U765 ( .A1(G164), .A2(G1384), .ZN(n721) );
  NOR2_X1 U766 ( .A1(n718), .A2(n721), .ZN(n824) );
  NAND2_X1 U767 ( .A1(n891), .A2(G140), .ZN(n691) );
  NAND2_X1 U768 ( .A1(G104), .A2(n892), .ZN(n690) );
  NAND2_X1 U769 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U770 ( .A(KEYINPUT34), .B(n692), .ZN(n698) );
  NAND2_X1 U771 ( .A1(n895), .A2(G116), .ZN(n693) );
  XNOR2_X1 U772 ( .A(n693), .B(KEYINPUT98), .ZN(n695) );
  NAND2_X1 U773 ( .A1(G128), .A2(n896), .ZN(n694) );
  NAND2_X1 U774 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U775 ( .A(KEYINPUT35), .B(n696), .Z(n697) );
  NOR2_X1 U776 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U777 ( .A(KEYINPUT36), .B(n699), .ZN(n906) );
  XOR2_X1 U778 ( .A(G2067), .B(KEYINPUT37), .Z(n700) );
  XNOR2_X1 U779 ( .A(KEYINPUT97), .B(n700), .ZN(n822) );
  NOR2_X1 U780 ( .A1(n906), .A2(n822), .ZN(n940) );
  NAND2_X1 U781 ( .A1(n824), .A2(n940), .ZN(n820) );
  NAND2_X1 U782 ( .A1(G107), .A2(n895), .ZN(n702) );
  NAND2_X1 U783 ( .A1(G131), .A2(n891), .ZN(n701) );
  NAND2_X1 U784 ( .A1(n702), .A2(n701), .ZN(n706) );
  NAND2_X1 U785 ( .A1(n896), .A2(G119), .ZN(n704) );
  NAND2_X1 U786 ( .A1(G95), .A2(n892), .ZN(n703) );
  NAND2_X1 U787 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U788 ( .A1(n706), .A2(n705), .ZN(n884) );
  INV_X1 U789 ( .A(G1991), .ZN(n857) );
  NOR2_X1 U790 ( .A1(n884), .A2(n857), .ZN(n716) );
  NAND2_X1 U791 ( .A1(G117), .A2(n895), .ZN(n708) );
  NAND2_X1 U792 ( .A1(G129), .A2(n896), .ZN(n707) );
  NAND2_X1 U793 ( .A1(n708), .A2(n707), .ZN(n712) );
  NAND2_X1 U794 ( .A1(n709), .A2(G105), .ZN(n710) );
  XOR2_X1 U795 ( .A(KEYINPUT38), .B(n710), .Z(n711) );
  NOR2_X1 U796 ( .A1(n712), .A2(n711), .ZN(n714) );
  NAND2_X1 U797 ( .A1(n891), .A2(G141), .ZN(n713) );
  NAND2_X1 U798 ( .A1(n714), .A2(n713), .ZN(n903) );
  AND2_X1 U799 ( .A1(G1996), .A2(n903), .ZN(n715) );
  NOR2_X1 U800 ( .A1(n716), .A2(n715), .ZN(n928) );
  INV_X1 U801 ( .A(n928), .ZN(n717) );
  NAND2_X1 U802 ( .A1(n717), .A2(n824), .ZN(n813) );
  NAND2_X1 U803 ( .A1(n820), .A2(n813), .ZN(n810) );
  XNOR2_X1 U804 ( .A(n718), .B(KEYINPUT99), .ZN(n722) );
  NAND2_X1 U805 ( .A1(n722), .A2(n721), .ZN(n764) );
  NAND2_X1 U806 ( .A1(G8), .A2(n764), .ZN(n796) );
  NOR2_X1 U807 ( .A1(G1981), .A2(G305), .ZN(n719) );
  XOR2_X1 U808 ( .A(n719), .B(KEYINPUT24), .Z(n720) );
  NOR2_X1 U809 ( .A1(n796), .A2(n720), .ZN(n808) );
  AND2_X2 U810 ( .A1(n722), .A2(n721), .ZN(n749) );
  NAND2_X1 U811 ( .A1(G1996), .A2(n749), .ZN(n723) );
  XNOR2_X1 U812 ( .A(KEYINPUT26), .B(n723), .ZN(n725) );
  NAND2_X1 U813 ( .A1(G1341), .A2(n764), .ZN(n724) );
  NAND2_X1 U814 ( .A1(n725), .A2(n724), .ZN(n726) );
  OR2_X1 U815 ( .A1(n1011), .A2(n726), .ZN(n738) );
  INV_X1 U816 ( .A(n995), .ZN(n737) );
  XNOR2_X1 U817 ( .A(n727), .B(KEYINPUT101), .ZN(n735) );
  NOR2_X1 U818 ( .A1(n749), .A2(G1348), .ZN(n729) );
  NOR2_X1 U819 ( .A1(G2067), .A2(n764), .ZN(n728) );
  NOR2_X1 U820 ( .A1(n729), .A2(n728), .ZN(n733) );
  NAND2_X1 U821 ( .A1(n749), .A2(G2072), .ZN(n730) );
  XNOR2_X1 U822 ( .A(n730), .B(KEYINPUT27), .ZN(n732) );
  AND2_X1 U823 ( .A1(G1956), .A2(n764), .ZN(n731) );
  NOR2_X1 U824 ( .A1(n732), .A2(n731), .ZN(n741) );
  NAND2_X1 U825 ( .A1(n741), .A2(n922), .ZN(n736) );
  AND2_X1 U826 ( .A1(n733), .A2(n736), .ZN(n734) );
  NAND2_X1 U827 ( .A1(n735), .A2(n734), .ZN(n747) );
  INV_X1 U828 ( .A(n736), .ZN(n740) );
  NAND2_X1 U829 ( .A1(n738), .A2(n737), .ZN(n739) );
  OR2_X1 U830 ( .A1(n740), .A2(n739), .ZN(n745) );
  NOR2_X1 U831 ( .A1(n741), .A2(n922), .ZN(n743) );
  XOR2_X1 U832 ( .A(KEYINPUT28), .B(KEYINPUT100), .Z(n742) );
  XNOR2_X1 U833 ( .A(n743), .B(n742), .ZN(n744) );
  AND2_X1 U834 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U835 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U836 ( .A(n748), .B(KEYINPUT29), .ZN(n753) );
  NAND2_X1 U837 ( .A1(G1961), .A2(n764), .ZN(n751) );
  XOR2_X1 U838 ( .A(KEYINPUT25), .B(G2078), .Z(n975) );
  NAND2_X1 U839 ( .A1(n749), .A2(n975), .ZN(n750) );
  NAND2_X1 U840 ( .A1(n751), .A2(n750), .ZN(n759) );
  NOR2_X1 U841 ( .A1(G301), .A2(n759), .ZN(n752) );
  NOR2_X1 U842 ( .A1(n753), .A2(n752), .ZN(n755) );
  XNOR2_X1 U843 ( .A(n755), .B(n754), .ZN(n778) );
  NOR2_X1 U844 ( .A1(G1966), .A2(n796), .ZN(n779) );
  NOR2_X1 U845 ( .A1(G2084), .A2(n764), .ZN(n781) );
  NOR2_X1 U846 ( .A1(n779), .A2(n781), .ZN(n756) );
  NAND2_X1 U847 ( .A1(G8), .A2(n756), .ZN(n757) );
  XNOR2_X1 U848 ( .A(KEYINPUT30), .B(n757), .ZN(n758) );
  NOR2_X1 U849 ( .A1(G168), .A2(n758), .ZN(n761) );
  AND2_X1 U850 ( .A1(G301), .A2(n759), .ZN(n760) );
  NOR2_X1 U851 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U852 ( .A(KEYINPUT31), .B(n762), .Z(n777) );
  INV_X1 U853 ( .A(G8), .ZN(n770) );
  NOR2_X1 U854 ( .A1(G1971), .A2(n796), .ZN(n763) );
  XNOR2_X1 U855 ( .A(KEYINPUT103), .B(n763), .ZN(n768) );
  NOR2_X1 U856 ( .A1(G2090), .A2(n764), .ZN(n765) );
  XNOR2_X1 U857 ( .A(KEYINPUT104), .B(n765), .ZN(n766) );
  NOR2_X1 U858 ( .A1(G166), .A2(n766), .ZN(n767) );
  NAND2_X1 U859 ( .A1(n768), .A2(n767), .ZN(n769) );
  OR2_X1 U860 ( .A1(n770), .A2(n769), .ZN(n772) );
  AND2_X1 U861 ( .A1(n777), .A2(n772), .ZN(n771) );
  NAND2_X1 U862 ( .A1(n778), .A2(n771), .ZN(n775) );
  INV_X1 U863 ( .A(n772), .ZN(n773) );
  OR2_X1 U864 ( .A1(n773), .A2(G286), .ZN(n774) );
  NAND2_X1 U865 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U866 ( .A(n776), .B(KEYINPUT32), .ZN(n785) );
  AND2_X1 U867 ( .A1(n778), .A2(n777), .ZN(n780) );
  NOR2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n783) );
  NAND2_X1 U869 ( .A1(G8), .A2(n781), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U871 ( .A1(n785), .A2(n784), .ZN(n793) );
  NOR2_X1 U872 ( .A1(G2090), .A2(G303), .ZN(n786) );
  NAND2_X1 U873 ( .A1(G8), .A2(n786), .ZN(n787) );
  NAND2_X1 U874 ( .A1(n793), .A2(n787), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n788), .A2(n796), .ZN(n806) );
  NOR2_X1 U876 ( .A1(G1976), .A2(G288), .ZN(n998) );
  NOR2_X1 U877 ( .A1(G1971), .A2(G303), .ZN(n789) );
  NOR2_X1 U878 ( .A1(n998), .A2(n789), .ZN(n791) );
  INV_X1 U879 ( .A(KEYINPUT33), .ZN(n790) );
  AND2_X1 U880 ( .A1(n791), .A2(n790), .ZN(n792) );
  NAND2_X1 U881 ( .A1(n793), .A2(n792), .ZN(n804) );
  NAND2_X1 U882 ( .A1(G1976), .A2(G288), .ZN(n1000) );
  INV_X1 U883 ( .A(n1000), .ZN(n794) );
  NOR2_X1 U884 ( .A1(n794), .A2(n796), .ZN(n795) );
  OR2_X1 U885 ( .A1(KEYINPUT33), .A2(n795), .ZN(n802) );
  NAND2_X1 U886 ( .A1(n998), .A2(KEYINPUT33), .ZN(n797) );
  NOR2_X1 U887 ( .A1(n797), .A2(n796), .ZN(n800) );
  XNOR2_X1 U888 ( .A(G1981), .B(G305), .ZN(n798) );
  XNOR2_X1 U889 ( .A(n798), .B(KEYINPUT105), .ZN(n1008) );
  INV_X1 U890 ( .A(n1008), .ZN(n799) );
  NOR2_X1 U891 ( .A1(n800), .A2(n799), .ZN(n801) );
  AND2_X1 U892 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U893 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U894 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U895 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U896 ( .A1(n810), .A2(n809), .ZN(n812) );
  XNOR2_X1 U897 ( .A(G1986), .B(G290), .ZN(n997) );
  NAND2_X1 U898 ( .A1(n997), .A2(n824), .ZN(n811) );
  NAND2_X1 U899 ( .A1(n812), .A2(n811), .ZN(n827) );
  NOR2_X1 U900 ( .A1(G1996), .A2(n903), .ZN(n936) );
  INV_X1 U901 ( .A(n813), .ZN(n817) );
  AND2_X1 U902 ( .A1(n857), .A2(n884), .ZN(n926) );
  NOR2_X1 U903 ( .A1(G1986), .A2(G290), .ZN(n814) );
  XNOR2_X1 U904 ( .A(KEYINPUT106), .B(n814), .ZN(n815) );
  NOR2_X1 U905 ( .A1(n926), .A2(n815), .ZN(n816) );
  NOR2_X1 U906 ( .A1(n817), .A2(n816), .ZN(n818) );
  NOR2_X1 U907 ( .A1(n936), .A2(n818), .ZN(n819) );
  XNOR2_X1 U908 ( .A(n819), .B(KEYINPUT39), .ZN(n821) );
  NAND2_X1 U909 ( .A1(n821), .A2(n820), .ZN(n823) );
  NAND2_X1 U910 ( .A1(n906), .A2(n822), .ZN(n938) );
  NAND2_X1 U911 ( .A1(n823), .A2(n938), .ZN(n825) );
  NAND2_X1 U912 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U913 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U914 ( .A(n828), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n921), .ZN(G217) );
  AND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U917 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U919 ( .A1(n831), .A2(n830), .ZN(G188) );
  NOR2_X1 U920 ( .A1(n833), .A2(n832), .ZN(G325) );
  XNOR2_X1 U921 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  INV_X1 U923 ( .A(G132), .ZN(G219) );
  INV_X1 U924 ( .A(G120), .ZN(G236) );
  INV_X1 U925 ( .A(G96), .ZN(G221) );
  INV_X1 U926 ( .A(G82), .ZN(G220) );
  INV_X1 U927 ( .A(G69), .ZN(G235) );
  XOR2_X1 U928 ( .A(G2454), .B(G2435), .Z(n835) );
  XNOR2_X1 U929 ( .A(G2438), .B(G2427), .ZN(n834) );
  XNOR2_X1 U930 ( .A(n835), .B(n834), .ZN(n842) );
  XOR2_X1 U931 ( .A(KEYINPUT107), .B(G2446), .Z(n837) );
  XNOR2_X1 U932 ( .A(G2443), .B(G2430), .ZN(n836) );
  XNOR2_X1 U933 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U934 ( .A(n838), .B(G2451), .Z(n840) );
  XNOR2_X1 U935 ( .A(G1341), .B(G1348), .ZN(n839) );
  XNOR2_X1 U936 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U937 ( .A(n842), .B(n841), .ZN(n843) );
  NAND2_X1 U938 ( .A1(n843), .A2(G14), .ZN(n844) );
  XOR2_X1 U939 ( .A(KEYINPUT108), .B(n844), .Z(G401) );
  XOR2_X1 U940 ( .A(G2100), .B(G2096), .Z(n846) );
  XNOR2_X1 U941 ( .A(KEYINPUT42), .B(G2678), .ZN(n845) );
  XNOR2_X1 U942 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U943 ( .A(KEYINPUT43), .B(G2090), .Z(n848) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2072), .ZN(n847) );
  XNOR2_X1 U945 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U946 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U947 ( .A(G2084), .B(G2078), .ZN(n851) );
  XNOR2_X1 U948 ( .A(n852), .B(n851), .ZN(G227) );
  XOR2_X1 U949 ( .A(G1981), .B(G1971), .Z(n854) );
  XNOR2_X1 U950 ( .A(G1966), .B(G1961), .ZN(n853) );
  XNOR2_X1 U951 ( .A(n854), .B(n853), .ZN(n865) );
  XOR2_X1 U952 ( .A(KEYINPUT110), .B(KEYINPUT41), .Z(n856) );
  XNOR2_X1 U953 ( .A(G1996), .B(KEYINPUT112), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(n861) );
  XOR2_X1 U955 ( .A(G1976), .B(G1956), .Z(n859) );
  XOR2_X1 U956 ( .A(n857), .B(G1986), .Z(n858) );
  XNOR2_X1 U957 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U958 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U959 ( .A(KEYINPUT111), .B(G2474), .ZN(n862) );
  XNOR2_X1 U960 ( .A(n863), .B(n862), .ZN(n864) );
  XNOR2_X1 U961 ( .A(n865), .B(n864), .ZN(G229) );
  NAND2_X1 U962 ( .A1(G124), .A2(n896), .ZN(n866) );
  XNOR2_X1 U963 ( .A(n866), .B(KEYINPUT44), .ZN(n868) );
  NAND2_X1 U964 ( .A1(n895), .A2(G112), .ZN(n867) );
  NAND2_X1 U965 ( .A1(n868), .A2(n867), .ZN(n872) );
  NAND2_X1 U966 ( .A1(n891), .A2(G136), .ZN(n870) );
  NAND2_X1 U967 ( .A1(G100), .A2(n892), .ZN(n869) );
  NAND2_X1 U968 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U969 ( .A1(n872), .A2(n871), .ZN(G162) );
  NAND2_X1 U970 ( .A1(G118), .A2(n895), .ZN(n874) );
  NAND2_X1 U971 ( .A1(G130), .A2(n896), .ZN(n873) );
  NAND2_X1 U972 ( .A1(n874), .A2(n873), .ZN(n879) );
  NAND2_X1 U973 ( .A1(n891), .A2(G142), .ZN(n876) );
  NAND2_X1 U974 ( .A1(G106), .A2(n892), .ZN(n875) );
  NAND2_X1 U975 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U976 ( .A(n877), .B(KEYINPUT45), .Z(n878) );
  NOR2_X1 U977 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U978 ( .A(n880), .B(n923), .ZN(n888) );
  XOR2_X1 U979 ( .A(KEYINPUT48), .B(KEYINPUT114), .Z(n882) );
  XNOR2_X1 U980 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n881) );
  XNOR2_X1 U981 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U982 ( .A(n883), .B(KEYINPUT46), .Z(n886) );
  XNOR2_X1 U983 ( .A(n884), .B(KEYINPUT113), .ZN(n885) );
  XNOR2_X1 U984 ( .A(n886), .B(n885), .ZN(n887) );
  XOR2_X1 U985 ( .A(n888), .B(n887), .Z(n890) );
  XNOR2_X1 U986 ( .A(G164), .B(G162), .ZN(n889) );
  XNOR2_X1 U987 ( .A(n890), .B(n889), .ZN(n902) );
  NAND2_X1 U988 ( .A1(n891), .A2(G139), .ZN(n894) );
  NAND2_X1 U989 ( .A1(G103), .A2(n892), .ZN(n893) );
  NAND2_X1 U990 ( .A1(n894), .A2(n893), .ZN(n901) );
  NAND2_X1 U991 ( .A1(G115), .A2(n895), .ZN(n898) );
  NAND2_X1 U992 ( .A1(G127), .A2(n896), .ZN(n897) );
  NAND2_X1 U993 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U994 ( .A(KEYINPUT47), .B(n899), .Z(n900) );
  NOR2_X1 U995 ( .A1(n901), .A2(n900), .ZN(n929) );
  XOR2_X1 U996 ( .A(n902), .B(n929), .Z(n905) );
  XOR2_X1 U997 ( .A(G160), .B(n903), .Z(n904) );
  XNOR2_X1 U998 ( .A(n905), .B(n904), .ZN(n907) );
  XOR2_X1 U999 ( .A(n907), .B(n906), .Z(n908) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n908), .ZN(G395) );
  INV_X1 U1001 ( .A(G301), .ZN(G171) );
  XOR2_X1 U1002 ( .A(G286), .B(G171), .Z(n909) );
  XNOR2_X1 U1003 ( .A(n909), .B(n1011), .ZN(n912) );
  XOR2_X1 U1004 ( .A(n995), .B(n910), .Z(n911) );
  XNOR2_X1 U1005 ( .A(n912), .B(n911), .ZN(n913) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n913), .ZN(G397) );
  OR2_X1 U1007 ( .A1(n920), .A2(G401), .ZN(n917) );
  NOR2_X1 U1008 ( .A1(G227), .A2(G229), .ZN(n914) );
  XOR2_X1 U1009 ( .A(KEYINPUT49), .B(n914), .Z(n915) );
  XNOR2_X1 U1010 ( .A(n915), .B(KEYINPUT117), .ZN(n916) );
  NOR2_X1 U1011 ( .A1(n917), .A2(n916), .ZN(n919) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1013 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(n920), .ZN(G319) );
  INV_X1 U1016 ( .A(G108), .ZN(G238) );
  INV_X1 U1017 ( .A(n921), .ZN(G223) );
  INV_X1 U1018 ( .A(n922), .ZN(G299) );
  XNOR2_X1 U1019 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n1029) );
  XNOR2_X1 U1020 ( .A(G160), .B(G2084), .ZN(n924) );
  NAND2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(n934) );
  XOR2_X1 U1024 ( .A(G2072), .B(n929), .Z(n931) );
  XOR2_X1 U1025 ( .A(G164), .B(G2078), .Z(n930) );
  NOR2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1027 ( .A(KEYINPUT50), .B(n932), .Z(n933) );
  NOR2_X1 U1028 ( .A1(n934), .A2(n933), .ZN(n943) );
  XOR2_X1 U1029 ( .A(G2090), .B(G162), .Z(n935) );
  NOR2_X1 U1030 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1031 ( .A(KEYINPUT51), .B(n937), .Z(n939) );
  NAND2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n941) );
  NOR2_X1 U1033 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1034 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1035 ( .A(KEYINPUT52), .B(n944), .ZN(n945) );
  XOR2_X1 U1036 ( .A(KEYINPUT118), .B(n945), .Z(n946) );
  INV_X1 U1037 ( .A(KEYINPUT55), .ZN(n990) );
  NAND2_X1 U1038 ( .A1(n946), .A2(n990), .ZN(n947) );
  NAND2_X1 U1039 ( .A1(n947), .A2(G29), .ZN(n1027) );
  XOR2_X1 U1040 ( .A(G4), .B(KEYINPUT125), .Z(n949) );
  XNOR2_X1 U1041 ( .A(G1348), .B(KEYINPUT59), .ZN(n948) );
  XNOR2_X1 U1042 ( .A(n949), .B(n948), .ZN(n953) );
  XNOR2_X1 U1043 ( .A(G1956), .B(G20), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(G1981), .B(G6), .ZN(n950) );
  NOR2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n956) );
  XNOR2_X1 U1047 ( .A(KEYINPUT124), .B(G1341), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(G19), .B(n954), .ZN(n955) );
  NOR2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(KEYINPUT60), .B(n957), .ZN(n961) );
  XNOR2_X1 U1051 ( .A(G1966), .B(G21), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(G5), .B(G1961), .ZN(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n968) );
  XNOR2_X1 U1055 ( .A(G1971), .B(G22), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(G23), .B(G1976), .ZN(n962) );
  NOR2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n965) );
  XOR2_X1 U1058 ( .A(G1986), .B(G24), .Z(n964) );
  NAND2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(KEYINPUT58), .B(n966), .ZN(n967) );
  NOR2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1062 ( .A(KEYINPUT61), .B(n969), .Z(n970) );
  NOR2_X1 U1063 ( .A1(G16), .A2(n970), .ZN(n1024) );
  XOR2_X1 U1064 ( .A(G2067), .B(G26), .Z(n972) );
  XOR2_X1 U1065 ( .A(G1996), .B(G32), .Z(n971) );
  NAND2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n982) );
  XNOR2_X1 U1067 ( .A(KEYINPUT119), .B(G2072), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(n973), .B(G33), .ZN(n980) );
  XOR2_X1 U1069 ( .A(G25), .B(G1991), .Z(n974) );
  NAND2_X1 U1070 ( .A1(n974), .A2(G28), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(G27), .B(n975), .ZN(n976) );
  XNOR2_X1 U1072 ( .A(KEYINPUT120), .B(n976), .ZN(n977) );
  NOR2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1076 ( .A(KEYINPUT53), .B(n983), .Z(n986) );
  XOR2_X1 U1077 ( .A(KEYINPUT54), .B(G34), .Z(n984) );
  XNOR2_X1 U1078 ( .A(G2084), .B(n984), .ZN(n985) );
  NAND2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n988) );
  XNOR2_X1 U1080 ( .A(G35), .B(G2090), .ZN(n987) );
  NOR2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1082 ( .A(n990), .B(n989), .Z(n992) );
  INV_X1 U1083 ( .A(G29), .ZN(n991) );
  NAND2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1085 ( .A1(n993), .A2(G11), .ZN(n994) );
  XNOR2_X1 U1086 ( .A(n994), .B(KEYINPUT121), .ZN(n1022) );
  XNOR2_X1 U1087 ( .A(G16), .B(KEYINPUT56), .ZN(n1020) );
  XOR2_X1 U1088 ( .A(G1348), .B(n995), .Z(n996) );
  NOR2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n1007) );
  INV_X1 U1090 ( .A(n998), .ZN(n999) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(n1001), .B(KEYINPUT122), .ZN(n1005) );
  XOR2_X1 U1093 ( .A(G303), .B(G1971), .Z(n1003) );
  XOR2_X1 U1094 ( .A(G299), .B(G1956), .Z(n1002) );
  NAND2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1017) );
  XNOR2_X1 U1098 ( .A(G1966), .B(G168), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(n1010), .B(KEYINPUT57), .ZN(n1015) );
  XOR2_X1 U1101 ( .A(G171), .B(G1961), .Z(n1013) );
  XNOR2_X1 U1102 ( .A(n1011), .B(G1341), .ZN(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(KEYINPUT123), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1110 ( .A(KEYINPUT126), .B(n1025), .ZN(n1026) );
  NAND2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1112 ( .A(n1029), .B(n1028), .Z(G150) );
  INV_X1 U1113 ( .A(G150), .ZN(G311) );
endmodule

