//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 0 0 0 1 1 1 1 1 1 1 1 0 1 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n565,
    new_n566, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n582,
    new_n583, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n622, new_n624, new_n625, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  OR2_X1    g031(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n457), .A2(KEYINPUT67), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(KEYINPUT67), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  XNOR2_X1  g038(.A(KEYINPUT68), .B(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(G137), .A3(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n464), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n471), .A2(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n465), .A2(new_n467), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(new_n472), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n479), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT69), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n482), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  NAND2_X1  g065(.A1(G114), .A2(G2104), .ZN(new_n491));
  INV_X1    g066(.A(G126), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n491), .B1(new_n478), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n473), .A2(G138), .A3(new_n472), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n493), .A2(G2105), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(G102), .A2(G2104), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT4), .A2(G138), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n478), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(new_n472), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n496), .A2(new_n500), .ZN(G164));
  NAND2_X1  g076(.A1(G75), .A2(G543), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(new_n507), .A2(G62), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n502), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n507), .A2(new_n509), .A3(G62), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  OAI21_X1  g087(.A(G651), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT73), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n516), .B2(G651), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n516), .A2(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n507), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AND3_X1   g099(.A1(new_n518), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n525));
  AOI21_X1  g100(.A(KEYINPUT70), .B1(new_n518), .B2(KEYINPUT6), .ZN(new_n526));
  OAI211_X1 g101(.A(G543), .B(new_n521), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n524), .A2(G88), .B1(new_n528), .B2(G50), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n529), .B(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n514), .A2(new_n531), .ZN(G303));
  INV_X1    g107(.A(G303), .ZN(G166));
  NAND2_X1  g108(.A1(new_n527), .A2(KEYINPUT74), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT74), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n520), .A2(new_n535), .A3(G543), .A4(new_n521), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n534), .A2(G51), .A3(new_n536), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n520), .A2(G89), .A3(new_n507), .A4(new_n521), .ZN(new_n538));
  AND2_X1   g113(.A1(G63), .A2(G651), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(KEYINPUT7), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT7), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n542), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n507), .A2(new_n539), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n537), .A2(new_n545), .ZN(G168));
  NAND3_X1  g121(.A1(new_n534), .A2(G52), .A3(new_n536), .ZN(new_n547));
  INV_X1    g122(.A(G64), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n548), .B1(new_n505), .B2(new_n506), .ZN(new_n549));
  AND2_X1   g124(.A1(G77), .A2(G543), .ZN(new_n550));
  OAI21_X1  g125(.A(G651), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n520), .A2(G90), .A3(new_n507), .A4(new_n521), .ZN(new_n552));
  AND2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n547), .A2(new_n553), .ZN(G171));
  NAND3_X1  g129(.A1(new_n534), .A2(G43), .A3(new_n536), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n556), .B1(new_n505), .B2(new_n506), .ZN(new_n557));
  AND2_X1   g132(.A1(G68), .A2(G543), .ZN(new_n558));
  OAI21_X1  g133(.A(G651), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n520), .A2(G81), .A3(new_n507), .A4(new_n521), .ZN(new_n560));
  AND2_X1   g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AND2_X1   g136(.A1(new_n555), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  AOI22_X1  g142(.A1(new_n507), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n568), .A2(new_n518), .ZN(new_n569));
  INV_X1    g144(.A(new_n522), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n570), .A2(G53), .A3(G543), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n571), .A2(KEYINPUT75), .A3(KEYINPUT9), .ZN(new_n572));
  NAND2_X1  g147(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n570), .A2(G53), .A3(G543), .A4(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n569), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n570), .A2(new_n507), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT76), .ZN(new_n577));
  OR3_X1    g152(.A1(new_n522), .A2(KEYINPUT76), .A3(new_n523), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n577), .A2(G91), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n575), .A2(new_n579), .ZN(G299));
  NAND2_X1  g155(.A1(new_n547), .A2(new_n553), .ZN(G301));
  AND3_X1   g156(.A1(new_n537), .A2(KEYINPUT77), .A3(new_n545), .ZN(new_n582));
  AOI21_X1  g157(.A(KEYINPUT77), .B1(new_n537), .B2(new_n545), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n582), .A2(new_n583), .ZN(G286));
  AND2_X1   g159(.A1(new_n577), .A2(new_n578), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G87), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n507), .A2(G74), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n528), .A2(G49), .B1(new_n587), .B2(G651), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n586), .A2(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(new_n585), .A2(G86), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n507), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n518), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n570), .A2(G48), .A3(G543), .ZN(new_n594));
  AND2_X1   g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n590), .A2(new_n595), .ZN(G305));
  AND2_X1   g171(.A1(new_n534), .A2(new_n536), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(G47), .ZN(new_n598));
  NAND2_X1  g173(.A1(G72), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G60), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n523), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n524), .A2(G85), .B1(new_n601), .B2(G651), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n598), .A2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n577), .A2(G92), .A3(new_n578), .ZN(new_n605));
  XOR2_X1   g180(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n523), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n597), .A2(G54), .B1(G651), .B2(new_n612), .ZN(new_n613));
  NAND4_X1  g188(.A1(new_n577), .A2(G92), .A3(new_n578), .A4(new_n606), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n609), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n604), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n604), .B1(new_n616), .B2(G868), .ZN(G321));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  MUX2_X1   g194(.A(G286), .B(G299), .S(new_n619), .Z(G297));
  MUX2_X1   g195(.A(G286), .B(G299), .S(new_n619), .Z(G280));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n616), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND2_X1  g198(.A1(new_n616), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n562), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT79), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g203(.A(KEYINPUT80), .ZN(new_n629));
  OR3_X1    g204(.A1(new_n629), .A2(new_n472), .A3(G111), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n472), .B2(G111), .ZN(new_n631));
  OR2_X1    g206(.A1(G99), .A2(G2105), .ZN(new_n632));
  NAND4_X1  g207(.A1(new_n630), .A2(G2104), .A3(new_n631), .A4(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(G135), .ZN(new_n634));
  INV_X1    g209(.A(G123), .ZN(new_n635));
  OAI221_X1 g210(.A(new_n633), .B1(new_n480), .B2(new_n634), .C1(new_n635), .C2(new_n483), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT81), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(G2096), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(G2096), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n469), .A2(new_n472), .A3(new_n473), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2100), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n639), .A2(new_n640), .A3(new_n644), .ZN(G156));
  XNOR2_X1  g220(.A(G2427), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2430), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(KEYINPUT14), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT83), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2451), .B(G2454), .Z(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(G14), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n656), .A2(new_n659), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(G401));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2072), .B(G2078), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT18), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n667), .B(KEYINPUT17), .Z(new_n671));
  INV_X1    g246(.A(new_n664), .ZN(new_n672));
  INV_X1    g247(.A(new_n665), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n672), .A2(new_n668), .A3(new_n673), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(new_n666), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n670), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT84), .ZN(new_n678));
  XOR2_X1   g253(.A(G2096), .B(G2100), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G227));
  XOR2_X1   g255(.A(G1971), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1956), .B(G2474), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1961), .B(G1966), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  NOR3_X1   g261(.A1(new_n682), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n682), .A2(new_n685), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT20), .Z(new_n689));
  AOI211_X1 g264(.A(new_n687), .B(new_n689), .C1(new_n682), .C2(new_n686), .ZN(new_n690));
  INV_X1    g265(.A(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  INV_X1    g270(.A(G1981), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n694), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(G229));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G23), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n586), .A2(new_n588), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(new_n700), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT33), .B(G1976), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n700), .A2(G6), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n590), .A2(new_n595), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(new_n700), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT32), .B(G1981), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n700), .A2(G22), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G166), .B2(new_n700), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT87), .B(G1971), .Z(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n712), .A2(new_n714), .ZN(new_n716));
  NAND4_X1  g291(.A1(new_n705), .A2(new_n710), .A3(new_n715), .A4(new_n716), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(KEYINPUT34), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(KEYINPUT34), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n720), .A2(G25), .ZN(new_n721));
  OAI21_X1  g296(.A(KEYINPUT85), .B1(G95), .B2(G2105), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  NOR3_X1   g298(.A1(KEYINPUT85), .A2(G95), .A3(G2105), .ZN(new_n724));
  OAI221_X1 g299(.A(G2104), .B1(G107), .B2(new_n472), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G131), .ZN(new_n726));
  INV_X1    g301(.A(G119), .ZN(new_n727));
  OAI221_X1 g302(.A(new_n725), .B1(new_n480), .B2(new_n726), .C1(new_n727), .C2(new_n483), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT86), .Z(new_n729));
  AOI21_X1  g304(.A(new_n721), .B1(new_n729), .B2(G29), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT35), .B(G1991), .Z(new_n731));
  AND2_X1   g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n700), .A2(G24), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(G290), .B2(G16), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n735), .A2(new_n691), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n735), .A2(new_n691), .ZN(new_n737));
  NOR4_X1   g312(.A1(new_n732), .A2(new_n733), .A3(new_n736), .A4(new_n737), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n718), .A2(new_n719), .A3(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT88), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(KEYINPUT36), .B1(new_n739), .B2(new_n740), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n720), .A2(G35), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G162), .B2(new_n720), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT29), .Z(new_n746));
  INV_X1    g321(.A(G2090), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n700), .A2(G5), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G171), .B2(new_n700), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G1961), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT96), .B(KEYINPUT23), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n700), .A2(G20), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G299), .B2(G16), .ZN(new_n755));
  INV_X1    g330(.A(G1956), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NOR3_X1   g332(.A1(new_n748), .A2(new_n751), .A3(new_n757), .ZN(new_n758));
  OR2_X1    g333(.A1(G104), .A2(G2105), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n759), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n760));
  INV_X1    g335(.A(G140), .ZN(new_n761));
  INV_X1    g336(.A(G128), .ZN(new_n762));
  OAI221_X1 g337(.A(new_n760), .B1(new_n480), .B2(new_n761), .C1(new_n762), .C2(new_n483), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(G29), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n720), .A2(G26), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G2067), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n720), .A2(G33), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT25), .Z(new_n773));
  AOI22_X1  g348(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n774));
  INV_X1    g349(.A(G139), .ZN(new_n775));
  OAI221_X1 g350(.A(new_n773), .B1(new_n472), .B2(new_n774), .C1(new_n480), .C2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n771), .B1(new_n776), .B2(G29), .ZN(new_n777));
  INV_X1    g352(.A(G2072), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT91), .ZN(new_n780));
  NOR2_X1   g355(.A1(G168), .A2(new_n700), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n700), .B2(G21), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT92), .B(G1966), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n770), .B(new_n780), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n700), .A2(G4), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n616), .B2(new_n700), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT89), .B(G1348), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n787), .A2(new_n788), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n784), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT93), .B(KEYINPUT31), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G11), .ZN(new_n794));
  INV_X1    g369(.A(G28), .ZN(new_n795));
  AOI21_X1  g370(.A(G29), .B1(new_n795), .B2(KEYINPUT30), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT94), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI22_X1  g373(.A1(new_n796), .A2(new_n797), .B1(KEYINPUT30), .B2(new_n795), .ZN(new_n799));
  OAI221_X1 g374(.A(new_n794), .B1(new_n798), .B2(new_n799), .C1(new_n777), .C2(new_n778), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT24), .ZN(new_n801));
  INV_X1    g376(.A(G34), .ZN(new_n802));
  AOI21_X1  g377(.A(G29), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n801), .B2(new_n802), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G160), .B2(new_n720), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n800), .B1(G2084), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n720), .A2(G27), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT95), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G164), .B2(new_n720), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n806), .B1(G2078), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n562), .A2(new_n700), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(new_n700), .B2(G19), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n813), .A2(G1341), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(G1341), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n809), .A2(G2078), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n782), .A2(new_n783), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n814), .A2(new_n815), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  OAI22_X1  g393(.A1(new_n638), .A2(new_n720), .B1(G2084), .B2(new_n805), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n720), .A2(G32), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n481), .A2(G141), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n484), .A2(G129), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n472), .A2(G105), .ZN(new_n823));
  NAND3_X1  g398(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT26), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n469), .A2(new_n823), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n821), .A2(new_n822), .A3(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n820), .B1(new_n830), .B2(new_n720), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT27), .B(G1996), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NOR4_X1   g408(.A1(new_n810), .A2(new_n818), .A3(new_n819), .A4(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n758), .A2(new_n792), .A3(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT97), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n741), .A2(new_n742), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n743), .A2(new_n836), .A3(new_n837), .ZN(G150));
  INV_X1    g413(.A(G150), .ZN(G311));
  NAND2_X1  g414(.A1(new_n616), .A2(G559), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n555), .A2(new_n561), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(KEYINPUT99), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT99), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n555), .A2(new_n561), .A3(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT98), .ZN(new_n845));
  AND2_X1   g420(.A1(G80), .A2(G543), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(new_n507), .B2(G67), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n845), .B1(new_n847), .B2(new_n518), .ZN(new_n848));
  INV_X1    g423(.A(G67), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(new_n505), .B2(new_n506), .ZN(new_n850));
  OAI211_X1 g425(.A(KEYINPUT98), .B(G651), .C1(new_n850), .C2(new_n846), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n534), .A2(G55), .A3(new_n536), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n524), .A2(G93), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n842), .A2(new_n844), .A3(new_n855), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n848), .A2(new_n851), .B1(new_n524), .B2(G93), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n562), .A2(new_n843), .A3(new_n853), .A4(new_n857), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n840), .B(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT39), .ZN(new_n863));
  AOI21_X1  g438(.A(G860), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n863), .B2(new_n862), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT101), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n855), .A2(G860), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT37), .Z(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(G145));
  XNOR2_X1  g444(.A(G164), .B(new_n763), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(new_n776), .Z(new_n871));
  XNOR2_X1  g446(.A(new_n728), .B(KEYINPUT103), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(new_n642), .Z(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n870), .B(new_n776), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n872), .B(new_n642), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n481), .A2(G142), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n484), .A2(G130), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n881));
  NOR3_X1   g456(.A1(new_n881), .A2(new_n472), .A3(G118), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n881), .B1(new_n472), .B2(G118), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n883), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n879), .B(new_n880), .C1(new_n882), .C2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n829), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n878), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n874), .A2(new_n886), .A3(new_n877), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n638), .B(G160), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(G162), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(KEYINPUT104), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n888), .A2(new_n895), .A3(new_n892), .A4(new_n889), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(KEYINPUT105), .B(G37), .Z(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n892), .B(KEYINPUT106), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n899), .B1(new_n900), .B2(new_n890), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g478(.A1(new_n855), .A2(new_n619), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n859), .B(KEYINPUT107), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(new_n624), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n579), .B(new_n575), .C1(new_n609), .C2(new_n615), .ZN(new_n907));
  NAND4_X1  g482(.A1(G299), .A2(new_n608), .A3(new_n614), .A4(new_n613), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n907), .A2(KEYINPUT41), .A3(new_n908), .ZN(new_n911));
  AOI21_X1  g486(.A(KEYINPUT41), .B1(new_n907), .B2(new_n908), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n910), .B1(new_n906), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n707), .A2(G303), .ZN(new_n915));
  NAND3_X1  g490(.A1(G305), .A2(new_n531), .A3(new_n514), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n702), .A2(G290), .ZN(new_n918));
  NAND3_X1  g493(.A1(G288), .A2(new_n598), .A3(new_n602), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n915), .A2(new_n918), .A3(new_n919), .A4(new_n916), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT42), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n914), .B(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n904), .B1(new_n925), .B2(new_n619), .ZN(G295));
  OAI21_X1  g501(.A(new_n904), .B1(new_n925), .B2(new_n619), .ZN(G331));
  INV_X1    g502(.A(KEYINPUT112), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n537), .A2(new_n545), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT77), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n537), .A2(KEYINPUT77), .A3(new_n545), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(G171), .A3(new_n932), .ZN(new_n933));
  NOR3_X1   g508(.A1(G171), .A2(KEYINPUT108), .A3(new_n929), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n935), .B1(G168), .B2(G301), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n933), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n859), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n856), .A2(new_n858), .ZN(new_n939));
  OAI21_X1  g514(.A(KEYINPUT108), .B1(G171), .B2(new_n929), .ZN(new_n940));
  NAND3_X1  g515(.A1(G168), .A2(new_n935), .A3(G301), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n939), .A2(new_n942), .A3(new_n933), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n909), .A2(new_n938), .A3(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n938), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n859), .A2(new_n937), .A3(KEYINPUT110), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n943), .A2(KEYINPUT109), .ZN(new_n948));
  AOI22_X1  g523(.A1(new_n940), .A2(new_n941), .B1(G286), .B2(G171), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(new_n950), .A3(new_n939), .ZN(new_n951));
  AOI22_X1  g526(.A1(new_n946), .A2(new_n947), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n923), .B(new_n944), .C1(new_n952), .C2(new_n913), .ZN(new_n953));
  INV_X1    g528(.A(G37), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT110), .B1(new_n859), .B2(new_n937), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n949), .A2(new_n945), .A3(new_n939), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n950), .B1(new_n949), .B2(new_n939), .ZN(new_n958));
  AND4_X1   g533(.A1(new_n950), .A2(new_n939), .A3(new_n933), .A4(new_n942), .ZN(new_n959));
  OAI22_X1  g534(.A1(new_n956), .A2(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT41), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n909), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n907), .A2(new_n908), .A3(KEYINPUT41), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n960), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n923), .B1(new_n965), .B2(new_n944), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT43), .B1(new_n955), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT111), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT111), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n969), .B(KEYINPUT43), .C1(new_n955), .C2(new_n966), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n907), .A2(new_n908), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n938), .A2(new_n943), .ZN(new_n972));
  OAI22_X1  g547(.A1(new_n960), .A2(new_n971), .B1(new_n913), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n923), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT43), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n975), .A2(new_n976), .A3(new_n898), .A4(new_n953), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n968), .A2(new_n970), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n976), .B1(new_n955), .B2(new_n966), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n975), .A2(KEYINPUT43), .A3(new_n898), .A4(new_n953), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n928), .B1(new_n980), .B2(new_n984), .ZN(new_n985));
  AOI211_X1 g560(.A(KEYINPUT112), .B(new_n983), .C1(new_n978), .C2(new_n979), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(G397));
  NAND2_X1  g562(.A1(new_n496), .A2(new_n500), .ZN(new_n988));
  INV_X1    g563(.A(G1384), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(KEYINPUT113), .B(G40), .ZN(new_n993));
  NOR4_X1   g568(.A1(new_n471), .A2(KEYINPUT114), .A3(new_n476), .A4(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n471), .A2(new_n476), .A3(new_n993), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n997));
  OR2_X1    g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n992), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G1996), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n999), .A2(new_n1000), .A3(new_n830), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT115), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n763), .B(G2067), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n830), .A2(new_n1000), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n999), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n999), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n728), .B(new_n731), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1003), .B(new_n1006), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(G290), .B(G1986), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1009), .B1(new_n999), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n998), .A2(new_n995), .ZN(new_n1013));
  AOI21_X1  g588(.A(G1384), .B1(new_n496), .B2(new_n500), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT45), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1013), .A2(new_n992), .A3(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1012), .B1(new_n1016), .B2(G2078), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n992), .A2(new_n1015), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1012), .A2(G2078), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(new_n1013), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1961), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n996), .A2(new_n997), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n1023));
  OAI22_X1  g598(.A1(new_n994), .A2(new_n1022), .B1(new_n1014), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n990), .A2(KEYINPUT50), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1021), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1017), .A2(new_n1020), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(G171), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1029));
  INV_X1    g604(.A(G2084), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1966), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1016), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(G168), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(G8), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n1029), .A2(new_n1030), .B1(new_n1016), .B2(new_n1032), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1036), .A2(G168), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT51), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1034), .A2(new_n1039), .A3(G8), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1028), .B1(new_n1041), .B2(KEYINPUT62), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n1043));
  NOR2_X1   g618(.A1(G305), .A2(G1981), .ZN(new_n1044));
  XOR2_X1   g619(.A(KEYINPUT118), .B(G86), .Z(new_n1045));
  OAI21_X1  g620(.A(new_n594), .B1(new_n576), .B2(new_n1045), .ZN(new_n1046));
  OR2_X1    g621(.A1(new_n1046), .A2(KEYINPUT119), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n592), .B1(new_n1046), .B2(KEYINPUT119), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n696), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1043), .B1(new_n1044), .B2(new_n1049), .ZN(new_n1050));
  OR2_X1    g625(.A1(new_n1050), .A2(KEYINPUT49), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1014), .B1(new_n1022), .B2(new_n994), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G8), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1050), .A2(KEYINPUT49), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1051), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1029), .A2(new_n747), .ZN(new_n1058));
  XOR2_X1   g633(.A(KEYINPUT116), .B(G1971), .Z(new_n1059));
  NAND2_X1  g634(.A1(new_n1016), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1054), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(G303), .A2(G8), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1062), .A2(KEYINPUT55), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1062), .A2(KEYINPUT55), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1061), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G1976), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1052), .B(G8), .C1(new_n1067), .C2(G288), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n1070));
  OR3_X1    g645(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(G288), .A2(new_n1070), .A3(new_n1067), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1068), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1057), .A2(new_n1066), .A3(new_n1074), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1013), .B(KEYINPUT121), .C1(new_n1023), .C2(new_n1014), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT121), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1024), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1025), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n747), .B1(new_n1079), .B2(KEYINPUT122), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n1081));
  AOI211_X1 g656(.A(new_n1081), .B(new_n1025), .C1(new_n1076), .C2(new_n1078), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1060), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(G8), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1065), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1075), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT62), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1038), .A2(new_n1087), .A3(new_n1040), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1042), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1057), .A2(new_n1067), .A3(new_n702), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(G1981), .B2(G305), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1066), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1057), .A2(new_n1074), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1091), .A2(new_n1055), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1036), .A2(new_n1054), .A3(G286), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT63), .B1(new_n1086), .B2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1095), .B(KEYINPUT63), .C1(new_n1065), .C2(new_n1061), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1097), .A2(new_n1075), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1089), .B(new_n1094), .C1(new_n1096), .C2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1018), .A2(G40), .A3(G160), .A4(new_n1019), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1100), .A2(new_n1017), .A3(G301), .A4(new_n1026), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT54), .B1(new_n1028), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1102), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1100), .A2(new_n1017), .A3(new_n1026), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1017), .A2(new_n1020), .A3(G301), .A4(new_n1026), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT125), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1108));
  OAI221_X1 g683(.A(KEYINPUT54), .B1(G301), .B2(new_n1104), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1086), .A2(new_n1103), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT61), .ZN(new_n1111));
  XOR2_X1   g686(.A(G299), .B(KEYINPUT57), .Z(new_n1112));
  INV_X1    g687(.A(new_n1025), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1024), .A2(new_n1077), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1024), .A2(new_n1077), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(new_n1117), .A3(new_n756), .ZN(new_n1118));
  OAI21_X1  g693(.A(KEYINPUT123), .B1(new_n1079), .B2(G1956), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1016), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT56), .B(G2072), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1112), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1123), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1112), .ZN(new_n1126));
  AOI211_X1 g701(.A(new_n1125), .B(new_n1126), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1111), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g703(.A(KEYINPUT58), .B(G1341), .ZN(new_n1129));
  OAI22_X1  g704(.A1(new_n1016), .A2(G1996), .B1(new_n1053), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n562), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1131), .A2(KEYINPUT59), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1131), .A2(KEYINPUT59), .ZN(new_n1133));
  INV_X1    g708(.A(new_n788), .ZN(new_n1134));
  OAI22_X1  g709(.A1(new_n1029), .A2(new_n1134), .B1(G2067), .B2(new_n1052), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT60), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n616), .A2(new_n1136), .ZN(new_n1137));
  OAI22_X1  g712(.A1(new_n1132), .A2(new_n1133), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  OR2_X1    g713(.A1(new_n1135), .A2(new_n616), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1135), .A2(new_n616), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1136), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1120), .A2(new_n1123), .A3(new_n1112), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1125), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1144));
  XOR2_X1   g719(.A(new_n1112), .B(KEYINPUT124), .Z(new_n1145));
  OAI211_X1 g720(.A(new_n1143), .B(KEYINPUT61), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1128), .A2(new_n1142), .A3(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1140), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(new_n1143), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1110), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1011), .B1(new_n1099), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n999), .B1(new_n829), .B2(new_n1004), .ZN(new_n1152));
  XOR2_X1   g727(.A(new_n1152), .B(KEYINPUT126), .Z(new_n1153));
  NAND2_X1  g728(.A1(new_n999), .A2(new_n1000), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT46), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  XOR2_X1   g731(.A(new_n1156), .B(KEYINPUT47), .Z(new_n1157));
  INV_X1    g732(.A(new_n731), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n729), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1003), .A2(new_n1006), .A3(new_n1159), .ZN(new_n1160));
  OR2_X1    g735(.A1(new_n763), .A2(G2067), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1007), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1007), .A2(G1986), .A3(G290), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1163), .B(KEYINPUT48), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1009), .A2(new_n1164), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1157), .A2(new_n1162), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1151), .A2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g742(.A1(new_n462), .A2(G227), .ZN(new_n1169));
  OAI21_X1  g743(.A(new_n1169), .B1(new_n661), .B2(new_n662), .ZN(new_n1170));
  OR2_X1    g744(.A1(new_n1170), .A2(KEYINPUT127), .ZN(new_n1171));
  NAND2_X1  g745(.A1(new_n1170), .A2(KEYINPUT127), .ZN(new_n1172));
  AND3_X1   g746(.A1(new_n1171), .A2(new_n698), .A3(new_n1172), .ZN(new_n1173));
  NAND3_X1  g747(.A1(new_n1173), .A2(new_n902), .A3(new_n978), .ZN(G225));
  INV_X1    g748(.A(G225), .ZN(G308));
endmodule


