//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0 0 1 1 1 0 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1257, new_n1258, new_n1259, new_n1260, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n203), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(new_n212), .A2(KEYINPUT0), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n218), .B1(KEYINPUT0), .B2(new_n212), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT64), .Z(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n205), .C2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT65), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n225), .A2(new_n226), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n209), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n232), .A2(KEYINPUT1), .ZN(new_n233));
  AND2_X1   g0033(.A1(new_n232), .A2(KEYINPUT1), .ZN(new_n234));
  NOR3_X1   g0034(.A1(new_n220), .A2(new_n233), .A3(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT66), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(KEYINPUT70), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(KEYINPUT67), .A3(new_n213), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(KEYINPUT67), .B1(new_n254), .B2(new_n213), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT8), .B(G58), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n214), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G150), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI22_X1  g0063(.A1(new_n259), .A2(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n203), .A2(G50), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n214), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n258), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n254), .A2(new_n213), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT67), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n255), .ZN(new_n271));
  INV_X1    g0071(.A(G1), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G13), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G20), .ZN(new_n275));
  INV_X1    g0075(.A(G50), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n276), .B1(new_n272), .B2(G20), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n271), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT68), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n273), .A2(new_n214), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n276), .ZN(new_n281));
  AND3_X1   g0081(.A1(new_n278), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n279), .B1(new_n278), .B2(new_n281), .ZN(new_n283));
  OAI211_X1 g0083(.A(KEYINPUT9), .B(new_n267), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  INV_X1    g0085(.A(G45), .ZN(new_n286));
  AOI21_X1  g0086(.A(G1), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G41), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(G1), .A3(G13), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n287), .A2(new_n289), .A3(G274), .ZN(new_n290));
  INV_X1    g0090(.A(G226), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n272), .B1(G41), .B2(G45), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n290), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT3), .B(G33), .ZN(new_n295));
  INV_X1    g0095(.A(G1698), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n295), .A2(G222), .A3(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n295), .A2(G223), .A3(G1698), .ZN(new_n298));
  INV_X1    g0098(.A(G77), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n297), .B(new_n298), .C1(new_n299), .C2(new_n295), .ZN(new_n300));
  INV_X1    g0100(.A(new_n289), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n294), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G190), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT69), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n300), .A2(new_n301), .ZN(new_n305));
  INV_X1    g0105(.A(new_n294), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n304), .B1(new_n307), .B2(G200), .ZN(new_n308));
  INV_X1    g0108(.A(G200), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n302), .A2(KEYINPUT69), .A3(new_n309), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n284), .B(new_n303), .C1(new_n308), .C2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n267), .B1(new_n282), .B2(new_n283), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT9), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT10), .B1(new_n311), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n307), .A2(new_n304), .A3(G200), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT69), .B1(new_n302), .B2(new_n309), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n317), .A2(new_n318), .B1(G190), .B2(new_n302), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT10), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n319), .A2(new_n320), .A3(new_n314), .A4(new_n284), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G169), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n307), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G179), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n302), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n312), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n301), .B1(new_n295), .B2(G107), .ZN(new_n328));
  INV_X1    g0128(.A(G238), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G1698), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(G232), .B2(G1698), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n328), .B1(new_n295), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G244), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n290), .B1(new_n333), .B2(new_n293), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G200), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n258), .A2(new_n280), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n338), .B(G77), .C1(G1), .C2(new_n214), .ZN(new_n339));
  NAND2_X1  g0139(.A1(G20), .A2(G77), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT15), .B(G87), .ZN(new_n341));
  OAI221_X1 g0141(.A(new_n340), .B1(new_n259), .B2(new_n263), .C1(new_n260), .C2(new_n341), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n342), .A2(new_n258), .B1(new_n299), .B2(new_n280), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n335), .A2(G190), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n337), .A2(new_n339), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n336), .A2(new_n323), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n339), .A2(new_n343), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n335), .A2(new_n325), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  AND4_X1   g0150(.A1(new_n253), .A2(new_n322), .A3(new_n327), .A4(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n327), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(new_n316), .B2(new_n321), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n253), .B1(new_n353), .B2(new_n350), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT3), .ZN(new_n356));
  INV_X1    g0156(.A(G33), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(KEYINPUT3), .A2(G33), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(new_n214), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT7), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT7), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n358), .A2(new_n362), .A3(new_n214), .A4(new_n359), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n361), .A2(G68), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G159), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT75), .B1(new_n263), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT75), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n262), .A2(new_n367), .A3(G159), .ZN(new_n368));
  XNOR2_X1  g0168(.A(G58), .B(G68), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n366), .A2(new_n368), .B1(new_n369), .B2(G20), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n364), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT16), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT74), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n374), .B1(new_n361), .B2(new_n363), .ZN(new_n375));
  AND2_X1   g0175(.A1(KEYINPUT3), .A2(G33), .ZN(new_n376));
  NOR2_X1   g0176(.A1(KEYINPUT3), .A2(G33), .ZN(new_n377));
  NOR3_X1   g0177(.A1(new_n376), .A2(new_n377), .A3(G20), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n374), .A2(new_n362), .ZN(new_n379));
  OAI21_X1  g0179(.A(G68), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI211_X1 g0180(.A(KEYINPUT16), .B(new_n370), .C1(new_n375), .C2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n373), .A2(new_n381), .A3(new_n258), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n259), .B1(new_n272), .B2(G20), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n338), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n280), .A2(new_n259), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI211_X1 g0186(.A(G223), .B(new_n296), .C1(new_n376), .C2(new_n377), .ZN(new_n387));
  OAI211_X1 g0187(.A(G226), .B(G1698), .C1(new_n376), .C2(new_n377), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G33), .A2(G87), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n301), .ZN(new_n391));
  INV_X1    g0191(.A(G190), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n289), .A2(G232), .A3(new_n292), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n290), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n391), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n394), .B1(new_n301), .B2(new_n390), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n396), .B1(G200), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n382), .A2(new_n386), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT17), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n384), .A2(new_n385), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n271), .B1(new_n371), .B2(new_n372), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n402), .B1(new_n403), .B2(new_n381), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n404), .A2(KEYINPUT17), .A3(new_n398), .ZN(new_n405));
  AND2_X1   g0205(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n391), .A2(G179), .A3(new_n395), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n323), .B2(new_n397), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n382), .A2(new_n386), .B1(new_n408), .B2(KEYINPUT76), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT76), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n407), .B(new_n410), .C1(new_n323), .C2(new_n397), .ZN(new_n411));
  NAND2_X1  g0211(.A1(KEYINPUT77), .A2(KEYINPUT18), .ZN(new_n412));
  OR2_X1    g0212(.A1(KEYINPUT77), .A2(KEYINPUT18), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n409), .A2(new_n411), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n382), .A2(new_n386), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n408), .A2(KEYINPUT76), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n415), .A2(new_n411), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(KEYINPUT77), .A3(KEYINPUT18), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n406), .A2(new_n414), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT73), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n214), .A2(G33), .A3(G77), .ZN(new_n421));
  OAI221_X1 g0221(.A(new_n421), .B1(new_n214), .B2(G68), .C1(new_n263), .C2(new_n276), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n258), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT11), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n280), .A2(new_n202), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n426), .B(KEYINPUT12), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n258), .A2(KEYINPUT11), .A3(new_n422), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n202), .B1(new_n272), .B2(G20), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n271), .A2(new_n275), .A3(new_n429), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n425), .A2(new_n427), .A3(new_n428), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT72), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n428), .A2(new_n430), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT72), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n433), .A2(new_n434), .A3(new_n425), .A4(new_n427), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT14), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT13), .ZN(new_n438));
  OAI211_X1 g0238(.A(G232), .B(G1698), .C1(new_n376), .C2(new_n377), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT71), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT71), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n295), .A2(new_n441), .A3(G232), .A4(G1698), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G97), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n295), .A2(G226), .A3(new_n296), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n440), .A2(new_n442), .A3(new_n443), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n301), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n290), .B1(new_n329), .B2(new_n293), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n438), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  AOI211_X1 g0249(.A(KEYINPUT13), .B(new_n447), .C1(new_n445), .C2(new_n301), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n437), .B(G169), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n446), .A2(new_n448), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT13), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n446), .A2(new_n438), .A3(new_n448), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n453), .A2(G179), .A3(new_n454), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n449), .A2(new_n450), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT14), .B1(new_n457), .B2(new_n323), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n436), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n431), .B1(new_n457), .B2(G190), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n453), .A2(new_n454), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G200), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n420), .B1(new_n459), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n437), .B1(new_n461), .B2(G169), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n451), .A2(new_n455), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n432), .B(new_n435), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(KEYINPUT73), .A3(new_n463), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n419), .B1(new_n465), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n355), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT19), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n214), .B1(new_n443), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(G87), .B2(new_n207), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n214), .B(G68), .C1(new_n376), .C2(new_n377), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n473), .B1(new_n260), .B2(new_n205), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n258), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n272), .A2(G33), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n271), .A2(G87), .A3(new_n275), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n280), .A2(new_n341), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n479), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n272), .A2(G45), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n289), .A2(G250), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n289), .A2(G274), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n485), .B1(new_n486), .B2(new_n484), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n295), .A2(G244), .A3(G1698), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G33), .A2(G116), .ZN(new_n489));
  OAI211_X1 g0289(.A(G238), .B(new_n296), .C1(new_n376), .C2(new_n377), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n487), .B1(new_n491), .B2(new_n301), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G190), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n483), .B(new_n493), .C1(new_n309), .C2(new_n492), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n275), .B(new_n480), .C1(new_n256), .C2(new_n257), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n479), .B(new_n482), .C1(new_n341), .C2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n492), .A2(new_n325), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n496), .B(new_n497), .C1(G169), .C2(new_n492), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n214), .B(G87), .C1(new_n376), .C2(new_n377), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT22), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT22), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n295), .A2(new_n502), .A3(new_n214), .A4(G87), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT24), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n489), .A2(G20), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT23), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(new_n214), .B2(G107), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n504), .A2(new_n505), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n505), .B1(new_n504), .B2(new_n510), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n258), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n280), .A2(new_n206), .ZN(new_n514));
  XNOR2_X1  g0314(.A(new_n514), .B(KEYINPUT25), .ZN(new_n515));
  INV_X1    g0315(.A(new_n495), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n515), .B1(G107), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g0318(.A(KEYINPUT5), .B(G41), .ZN(new_n519));
  INV_X1    g0319(.A(new_n484), .ZN(new_n520));
  INV_X1    g0320(.A(new_n213), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n288), .ZN(new_n522));
  INV_X1    g0322(.A(G274), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n523), .B1(new_n521), .B2(new_n288), .ZN(new_n524));
  OR2_X1    g0324(.A1(KEYINPUT5), .A2(G41), .ZN(new_n525));
  NAND2_X1  g0325(.A1(KEYINPUT5), .A2(G41), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n484), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n522), .A2(G264), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(G250), .A2(G1698), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n529), .B1(new_n224), .B2(G1698), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n530), .A2(new_n295), .B1(G33), .B2(G294), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n301), .B1(new_n531), .B2(KEYINPUT82), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n223), .A2(new_n296), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n224), .A2(G1698), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n533), .B(new_n534), .C1(new_n376), .C2(new_n377), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G33), .A2(G294), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT82), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(G179), .B(new_n528), .C1(new_n532), .C2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT83), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n519), .A2(new_n520), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n542), .A2(G264), .A3(new_n289), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n527), .A2(new_n524), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n531), .A2(KEYINPUT82), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n289), .B1(new_n537), .B2(new_n538), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n540), .B(new_n541), .C1(new_n548), .C2(new_n323), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n548), .A2(KEYINPUT83), .A3(G179), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n518), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n548), .A2(new_n392), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n548), .A2(G200), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n513), .B(new_n517), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n499), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(G116), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n274), .A2(G20), .A3(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n254), .A2(new_n213), .B1(G20), .B2(new_n556), .ZN(new_n558));
  NAND2_X1  g0358(.A1(G33), .A2(G283), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n559), .B(new_n214), .C1(G33), .C2(new_n205), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n558), .A2(KEYINPUT20), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT20), .B1(new_n558), .B2(new_n560), .ZN(new_n562));
  OAI221_X1 g0362(.A(new_n557), .B1(new_n561), .B2(new_n562), .C1(new_n495), .C2(new_n556), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n522), .A2(G270), .B1(new_n524), .B2(new_n527), .ZN(new_n564));
  OAI211_X1 g0364(.A(G264), .B(G1698), .C1(new_n376), .C2(new_n377), .ZN(new_n565));
  OAI211_X1 g0365(.A(G257), .B(new_n296), .C1(new_n376), .C2(new_n377), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n358), .A2(G303), .A3(new_n359), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n301), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n323), .B1(new_n564), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n563), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT21), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n564), .A2(G179), .A3(new_n569), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n563), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n563), .A2(KEYINPUT21), .A3(new_n570), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n564), .A2(new_n569), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G200), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n495), .A2(new_n556), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n557), .B1(new_n561), .B2(new_n562), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n564), .A2(new_n569), .A3(G190), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n579), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT81), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OR2_X1    g0386(.A1(new_n584), .A2(new_n585), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n577), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n527), .A2(new_n301), .A3(new_n224), .ZN(new_n589));
  OAI211_X1 g0389(.A(G244), .B(new_n296), .C1(new_n376), .C2(new_n377), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT4), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n295), .A2(KEYINPUT4), .A3(G244), .A4(new_n296), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n295), .A2(G250), .A3(G1698), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n559), .A4(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n589), .B1(new_n595), .B2(new_n301), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n544), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G169), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n596), .A2(G179), .A3(new_n544), .ZN(new_n599));
  XNOR2_X1  g0399(.A(G97), .B(G107), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT6), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT78), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT78), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(KEYINPUT6), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT79), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n603), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(G97), .B1(new_n603), .B2(new_n605), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n601), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n603), .A2(new_n605), .A3(new_n606), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n600), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n609), .A2(G20), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n361), .A2(G107), .A3(new_n363), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n263), .A2(new_n299), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n258), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n280), .A2(new_n205), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(new_n495), .B2(new_n205), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n598), .A2(new_n599), .B1(new_n617), .B2(new_n620), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n613), .A2(new_n615), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n609), .A2(G20), .A3(new_n611), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n271), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n624), .A2(KEYINPUT80), .A3(new_n619), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT80), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n626), .B1(new_n617), .B2(new_n620), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n597), .A2(G200), .ZN(new_n629));
  INV_X1    g0429(.A(new_n544), .ZN(new_n630));
  AOI211_X1 g0430(.A(new_n589), .B(new_n630), .C1(new_n595), .C2(new_n301), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(G190), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n621), .B1(new_n628), .B2(new_n633), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n472), .A2(new_n555), .A3(new_n588), .A4(new_n634), .ZN(G372));
  NAND2_X1  g0435(.A1(new_n401), .A2(new_n405), .ZN(new_n636));
  INV_X1    g0436(.A(new_n349), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n463), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n636), .B1(new_n468), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n415), .A2(new_n408), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT18), .ZN(new_n641));
  XNOR2_X1  g0441(.A(new_n640), .B(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n322), .B1(new_n639), .B2(new_n643), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n551), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n491), .A2(new_n301), .ZN(new_n648));
  INV_X1    g0448(.A(new_n487), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n650), .A2(KEYINPUT84), .A3(G200), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT84), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n492), .B2(new_n309), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n651), .A2(new_n653), .A3(new_n493), .A4(new_n483), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n654), .A2(new_n498), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT80), .B1(new_n624), .B2(new_n619), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n617), .A2(new_n626), .A3(new_n620), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n656), .A2(new_n657), .A3(new_n629), .A4(new_n632), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n599), .B1(new_n631), .B2(new_n323), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n617), .A2(new_n620), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n655), .A2(new_n658), .A3(new_n554), .A4(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n647), .A2(new_n662), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n656), .A2(new_n657), .B1(new_n598), .B2(new_n599), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n655), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n659), .A2(new_n494), .A3(new_n498), .A4(new_n660), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT26), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n666), .A2(new_n498), .A3(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n663), .A2(new_n669), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n327), .B(new_n644), .C1(new_n471), .C2(new_n670), .ZN(G369));
  INV_X1    g0471(.A(new_n518), .ZN(new_n672));
  OR3_X1    g0472(.A1(new_n273), .A2(KEYINPUT27), .A3(G20), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT27), .B1(new_n273), .B2(G20), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n551), .B(new_n554), .C1(new_n672), .C2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n551), .B2(new_n678), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n582), .A2(new_n678), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT85), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n588), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT86), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n682), .A2(new_n645), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n684), .B1(new_n683), .B2(new_n685), .ZN(new_n687));
  OAI211_X1 g0487(.A(G330), .B(new_n680), .C1(new_n686), .C2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n551), .A2(new_n677), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n645), .A2(new_n677), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n551), .A2(new_n554), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n688), .A2(new_n692), .ZN(G399));
  INV_X1    g0493(.A(new_n210), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G41), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(G1), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n216), .B2(new_n696), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT87), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n665), .B1(new_n655), .B2(new_n664), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n498), .B1(new_n667), .B2(KEYINPUT26), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n654), .A2(new_n498), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n552), .A2(new_n553), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n705), .B1(new_n672), .B2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n634), .A2(new_n707), .A3(new_n646), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n677), .B1(new_n704), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(KEYINPUT29), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n670), .A2(new_n677), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n710), .B1(new_n711), .B2(KEYINPUT29), .ZN(new_n712));
  INV_X1    g0512(.A(G330), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n574), .A2(new_n548), .A3(new_n492), .A4(new_n596), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT30), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n547), .A2(new_n546), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n717), .A2(new_n528), .A3(new_n492), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(KEYINPUT30), .A3(new_n574), .A4(new_n596), .ZN(new_n719));
  AOI21_X1  g0519(.A(G179), .B1(new_n717), .B2(new_n528), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n720), .A2(new_n597), .A3(new_n650), .A4(new_n578), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n716), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n722), .A2(KEYINPUT31), .A3(new_n677), .ZN(new_n723));
  AOI21_X1  g0523(.A(KEYINPUT31), .B1(new_n722), .B2(new_n677), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n555), .A2(new_n634), .A3(new_n588), .A4(new_n678), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n713), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n712), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n701), .B1(new_n730), .B2(G1), .ZN(G364));
  OR3_X1    g0531(.A1(new_n686), .A2(new_n687), .A3(G330), .ZN(new_n732));
  OAI21_X1  g0532(.A(G330), .B1(new_n686), .B2(new_n687), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n214), .A2(G13), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n272), .B1(new_n734), .B2(G45), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n695), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n732), .A2(new_n733), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n295), .A2(new_n210), .ZN(new_n740));
  INV_X1    g0540(.A(G355), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n740), .A2(new_n741), .B1(G116), .B2(new_n210), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n694), .A2(new_n295), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n744), .B1(new_n286), .B2(new_n217), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n251), .A2(G45), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n742), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OR3_X1    g0547(.A1(KEYINPUT88), .A2(G13), .A3(G33), .ZN(new_n748));
  OAI21_X1  g0548(.A(KEYINPUT88), .B1(G13), .B2(G33), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n214), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n213), .B1(G20), .B2(new_n323), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n737), .B1(new_n747), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n295), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n214), .A2(new_n392), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(new_n325), .A3(G200), .ZN(new_n758));
  INV_X1    g0558(.A(G303), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n756), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  XOR2_X1   g0560(.A(new_n760), .B(KEYINPUT93), .Z(new_n761));
  NOR2_X1   g0561(.A1(new_n325), .A2(G200), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G322), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n214), .A2(G190), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(new_n762), .ZN(new_n766));
  INV_X1    g0566(.A(G311), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n763), .A2(new_n764), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G190), .ZN(new_n770));
  NOR2_X1   g0570(.A1(KEYINPUT33), .A2(G317), .ZN(new_n771));
  AND2_X1   g0571(.A1(KEYINPUT33), .A2(G317), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(G294), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G179), .A2(G200), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n214), .B1(new_n775), .B2(G190), .ZN(new_n776));
  INV_X1    g0576(.A(G326), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n769), .A2(new_n392), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n773), .B1(new_n774), .B2(new_n776), .C1(new_n777), .C2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n765), .A2(new_n775), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n768), .B(new_n780), .C1(G329), .C2(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n765), .A2(new_n325), .A3(G200), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT91), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT92), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G283), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n761), .B(new_n783), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n790), .A2(new_n206), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n781), .A2(new_n365), .ZN(new_n794));
  INV_X1    g0594(.A(KEYINPUT32), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n295), .B1(new_n222), .B2(new_n758), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n776), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n794), .A2(new_n795), .B1(new_n797), .B2(G97), .ZN(new_n798));
  INV_X1    g0598(.A(new_n770), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n202), .B2(new_n799), .ZN(new_n800));
  OR3_X1    g0600(.A1(new_n793), .A2(new_n796), .A3(new_n800), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n763), .A2(new_n201), .B1(new_n766), .B2(new_n299), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT89), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n802), .A2(new_n803), .B1(new_n276), .B2(new_n779), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(new_n803), .B2(new_n802), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT90), .Z(new_n806));
  OAI21_X1  g0606(.A(new_n792), .B1(new_n801), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n755), .B1(new_n807), .B2(new_n752), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n683), .A2(new_n685), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n808), .B1(new_n809), .B2(new_n751), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n739), .A2(new_n810), .ZN(G396));
  NAND2_X1  g0611(.A1(new_n347), .A2(new_n677), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n637), .B1(new_n345), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n637), .A2(new_n678), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n711), .B(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n737), .B1(new_n817), .B2(new_n728), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n728), .B2(new_n817), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n750), .A2(new_n752), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n738), .B1(new_n299), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n750), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n789), .A2(G68), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n276), .B2(new_n758), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT95), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n756), .B1(new_n782), .B2(G132), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n825), .B(new_n826), .C1(new_n201), .C2(new_n776), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(KEYINPUT96), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n763), .ZN(new_n831));
  XOR2_X1   g0631(.A(KEYINPUT94), .B(G143), .Z(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n766), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n831), .A2(new_n833), .B1(new_n834), .B2(G159), .ZN(new_n835));
  INV_X1    g0635(.A(G137), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n835), .B1(new_n799), .B2(new_n261), .C1(new_n836), .C2(new_n779), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT34), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(new_n828), .B2(KEYINPUT96), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n789), .A2(G87), .ZN(new_n841));
  INV_X1    g0641(.A(new_n758), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n842), .A2(G107), .B1(new_n782), .B2(G311), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n556), .B2(new_n766), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n799), .A2(new_n791), .B1(new_n779), .B2(new_n759), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n756), .B1(new_n776), .B2(new_n205), .C1(new_n774), .C2(new_n763), .ZN(new_n846));
  NOR3_X1   g0646(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n830), .A2(new_n840), .B1(new_n841), .B2(new_n847), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n821), .B1(new_n822), .B2(new_n816), .C1(new_n848), .C2(new_n753), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n819), .A2(new_n849), .ZN(G384));
  NAND2_X1  g0650(.A1(new_n725), .A2(new_n726), .ZN(new_n851));
  INV_X1    g0651(.A(new_n813), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n814), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n432), .A2(new_n435), .A3(new_n677), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT97), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n459), .B2(new_n464), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT97), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n854), .B(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n468), .A2(new_n463), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n853), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n417), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n399), .B1(new_n404), .B2(new_n675), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT98), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT37), .B1(new_n409), .B2(new_n411), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n382), .A2(new_n386), .A3(new_n398), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n675), .B1(new_n382), .B2(new_n386), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT98), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n865), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n370), .B1(new_n375), .B2(new_n380), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n372), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(new_n381), .A3(new_n258), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n386), .ZN(new_n874));
  INV_X1    g0674(.A(new_n675), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n408), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(new_n877), .A3(new_n399), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n864), .A2(new_n870), .B1(KEYINPUT37), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n412), .B1(new_n409), .B2(new_n411), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n636), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n876), .B1(new_n881), .B2(new_n414), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  NOR3_X1   g0683(.A1(new_n879), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n878), .A2(KEYINPUT37), .ZN(new_n885));
  NOR3_X1   g0685(.A1(new_n862), .A2(KEYINPUT98), .A3(new_n863), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n869), .B1(new_n865), .B2(new_n868), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n876), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n419), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT38), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n851), .B(new_n860), .C1(new_n884), .C2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT40), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n856), .A2(new_n859), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n894), .A2(new_n851), .A3(new_n816), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n861), .B1(new_n868), .B2(new_n640), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(new_n864), .B2(new_n870), .ZN(new_n897));
  INV_X1    g0697(.A(new_n867), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n642), .B2(new_n406), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n883), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n888), .A2(KEYINPUT38), .A3(new_n890), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n893), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n892), .A2(new_n893), .B1(new_n895), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n472), .A2(new_n851), .ZN(new_n905));
  OAI21_X1  g0705(.A(G330), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n904), .B2(new_n905), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n900), .A2(new_n901), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT39), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n459), .A2(new_n678), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n883), .B1(new_n879), .B2(new_n882), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(new_n901), .A3(KEYINPUT39), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n910), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n856), .A2(new_n859), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n816), .B(new_n678), .C1(new_n663), .C2(new_n669), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n916), .B1(new_n814), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n913), .A2(new_n901), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n918), .A2(new_n919), .B1(new_n643), .B2(new_n675), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n915), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n644), .A2(new_n327), .ZN(new_n922));
  OR2_X1    g0722(.A1(new_n663), .A2(new_n669), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT29), .B1(new_n923), .B2(new_n678), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n709), .A2(KEYINPUT29), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n922), .B1(new_n926), .B2(new_n472), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n921), .B(new_n927), .Z(new_n928));
  OAI22_X1  g0728(.A1(new_n907), .A2(new_n928), .B1(new_n272), .B2(new_n734), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n928), .B2(new_n907), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n609), .A2(new_n611), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT35), .ZN(new_n932));
  OAI211_X1 g0732(.A(G116), .B(new_n215), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(new_n932), .B2(new_n931), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT36), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n217), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n276), .A2(G68), .ZN(new_n937));
  AOI211_X1 g0737(.A(new_n272), .B(G13), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  OR3_X1    g0738(.A1(new_n930), .A2(new_n935), .A3(new_n938), .ZN(G367));
  AND2_X1   g0739(.A1(new_n690), .A2(new_n691), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT42), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n658), .B(new_n661), .C1(new_n628), .C2(new_n678), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n664), .A2(new_n677), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n940), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n551), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n677), .B1(new_n947), .B2(new_n661), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n941), .B1(new_n940), .B2(new_n944), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n948), .A2(KEYINPUT99), .A3(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT99), .ZN(new_n951));
  INV_X1    g0751(.A(new_n944), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n690), .A2(new_n691), .ZN(new_n953));
  OAI21_X1  g0753(.A(KEYINPUT42), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n551), .B1(new_n942), .B2(new_n943), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n678), .B1(new_n955), .B2(new_n621), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n951), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n945), .B1(new_n950), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(KEYINPUT100), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n483), .A2(new_n678), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n655), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n498), .B2(new_n960), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n963));
  OAI21_X1  g0763(.A(KEYINPUT99), .B1(new_n948), .B2(new_n949), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n954), .A2(new_n956), .A3(new_n951), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT100), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n966), .A2(new_n967), .A3(new_n945), .ZN(new_n968));
  AND3_X1   g0768(.A1(new_n959), .A2(new_n963), .A3(new_n968), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n962), .B(KEYINPUT43), .Z(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(new_n959), .B2(new_n968), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n969), .A2(new_n972), .B1(new_n688), .B2(new_n952), .ZN(new_n973));
  INV_X1    g0773(.A(new_n688), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n692), .A2(new_n944), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT45), .ZN(new_n976));
  XNOR2_X1  g0776(.A(KEYINPUT101), .B(KEYINPUT44), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n952), .B(new_n977), .C1(new_n940), .C2(new_n689), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT101), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n979), .B(KEYINPUT44), .C1(new_n692), .C2(new_n944), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n974), .B1(new_n976), .B2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT45), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n975), .B(new_n983), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n984), .A2(new_n688), .A3(new_n980), .A4(new_n978), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n953), .B1(new_n680), .B2(new_n690), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n733), .A2(new_n988), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n987), .B(G330), .C1(new_n686), .C2(new_n687), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n991), .A2(new_n728), .A3(new_n712), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n730), .B1(new_n986), .B2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n695), .B(KEYINPUT41), .Z(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n735), .ZN(new_n997));
  INV_X1    g0797(.A(new_n968), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n967), .B1(new_n966), .B2(new_n945), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n970), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n688), .A2(new_n952), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n959), .A2(new_n968), .A3(new_n963), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n973), .A2(new_n997), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n341), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n754), .B1(new_n694), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n243), .A2(new_n743), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n738), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n758), .A2(new_n556), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n1009), .A2(KEYINPUT46), .B1(new_n767), .B2(new_n779), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(KEYINPUT46), .B2(new_n1009), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n766), .A2(new_n791), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n756), .B1(new_n763), .B2(new_n759), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1012), .B(new_n1013), .C1(G317), .C2(new_n782), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n788), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(G97), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n797), .A2(G107), .B1(G294), .B2(new_n770), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1011), .A2(new_n1014), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n295), .B1(new_n788), .B2(new_n299), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1019), .A2(KEYINPUT103), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(KEYINPUT103), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n766), .A2(new_n276), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n758), .A2(new_n201), .B1(new_n781), .B2(new_n836), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1022), .B(new_n1023), .C1(G159), .C2(new_n770), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1020), .A2(new_n1021), .A3(new_n1024), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n779), .A2(new_n832), .B1(new_n763), .B2(new_n261), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n776), .A2(new_n202), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT102), .Z(new_n1029));
  OAI21_X1  g0829(.A(new_n1018), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT47), .Z(new_n1031));
  OAI221_X1 g0831(.A(new_n1008), .B1(new_n962), .B2(new_n751), .C1(new_n1031), .C2(new_n753), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1004), .A2(new_n1032), .ZN(G387));
  NAND2_X1  g0833(.A1(new_n991), .A2(new_n736), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT104), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n680), .A2(new_n751), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n740), .A2(new_n697), .B1(G107), .B2(new_n210), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n240), .A2(new_n286), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n697), .ZN(new_n1039));
  AOI211_X1 g0839(.A(G45), .B(new_n1039), .C1(G68), .C2(G77), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n259), .A2(G50), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT50), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n744), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1037), .B1(new_n1038), .B2(new_n1043), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n758), .A2(new_n774), .B1(new_n776), .B2(new_n791), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G317), .A2(new_n831), .B1(new_n834), .B2(G303), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n799), .B2(new_n767), .C1(new_n764), .C2(new_n779), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT48), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1045), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n1048), .B2(new_n1047), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT49), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n756), .B1(new_n781), .B2(new_n777), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n1015), .B2(G116), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n789), .A2(G97), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n842), .A2(G77), .B1(new_n782), .B2(G150), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n276), .B2(new_n763), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n295), .B1(new_n766), .B2(new_n202), .C1(new_n799), .C2(new_n259), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n779), .A2(new_n365), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n776), .A2(new_n341), .ZN(new_n1059));
  NOR4_X1   g0859(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1051), .A2(new_n1053), .B1(new_n1054), .B2(new_n1060), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n737), .B1(new_n754), .B2(new_n1044), .C1(new_n1061), .C2(new_n753), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT105), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1035), .B1(new_n1036), .B2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n729), .A2(new_n990), .A3(new_n989), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1065), .A2(new_n695), .A3(new_n992), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1064), .A2(new_n1066), .ZN(G393));
  OR2_X1    g0867(.A1(new_n986), .A2(new_n992), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n986), .A2(new_n992), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1068), .A2(new_n695), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n735), .B1(new_n986), .B2(KEYINPUT106), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(KEYINPUT106), .B2(new_n986), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n793), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n831), .A2(G311), .B1(G317), .B2(new_n778), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT52), .Z(new_n1075));
  NOR2_X1   g0875(.A1(new_n776), .A2(new_n556), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n756), .B1(new_n766), .B2(new_n774), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1076), .B(new_n1077), .C1(G303), .C2(new_n770), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n758), .A2(new_n791), .B1(new_n781), .B2(new_n764), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT108), .Z(new_n1080));
  NAND4_X1  g0880(.A1(new_n1073), .A2(new_n1075), .A3(new_n1078), .A4(new_n1080), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n779), .A2(new_n261), .B1(new_n763), .B2(new_n365), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT51), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n758), .A2(new_n202), .B1(new_n832), .B2(new_n781), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n799), .A2(new_n276), .B1(new_n776), .B2(new_n299), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n295), .B1(new_n766), .B2(new_n259), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n841), .A2(new_n1083), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n753), .B1(new_n1081), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n248), .A2(new_n743), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n754), .B1(G97), .B2(new_n694), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n738), .B(new_n1089), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT109), .ZN(new_n1093));
  OAI21_X1  g0893(.A(KEYINPUT107), .B1(new_n944), .B2(new_n751), .ZN(new_n1094));
  OR3_X1    g0894(.A1(new_n944), .A2(KEYINPUT107), .A3(new_n751), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1070), .A2(new_n1072), .A3(new_n1096), .ZN(G390));
  INV_X1    g0897(.A(new_n914), .ZN(new_n1098));
  AOI21_X1  g0898(.A(KEYINPUT39), .B1(new_n900), .B2(new_n901), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n1098), .A2(new_n1099), .B1(new_n918), .B2(new_n912), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n677), .B(new_n813), .C1(new_n704), .C2(new_n708), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n894), .B1(new_n1101), .B2(new_n815), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n912), .B1(new_n900), .B2(new_n901), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n1102), .A2(KEYINPUT110), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(KEYINPUT110), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1100), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n860), .A2(new_n727), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n851), .A2(G330), .A3(new_n816), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n916), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n815), .B1(new_n709), .B2(new_n852), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1111), .A2(new_n1112), .A3(new_n1107), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n917), .A2(new_n814), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1110), .A2(new_n916), .B1(new_n860), .B2(new_n727), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT111), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n471), .B2(new_n728), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n355), .A2(KEYINPUT111), .A3(new_n470), .A4(new_n727), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1116), .A2(new_n927), .A3(new_n1120), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1100), .B(new_n1107), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1109), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1116), .A2(new_n927), .A3(new_n1120), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT112), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1124), .B(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1109), .A2(new_n1122), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n695), .B(new_n1123), .C1(new_n1126), .C2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n750), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n295), .B1(new_n788), .B2(new_n276), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1131), .A2(KEYINPUT113), .B1(G125), .B2(new_n782), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(KEYINPUT113), .B2(new_n1131), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT114), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(KEYINPUT54), .B(G143), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n831), .A2(G132), .B1(new_n834), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n842), .A2(G150), .ZN(new_n1138));
  XOR2_X1   g0938(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1137), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1138), .A2(new_n1140), .B1(new_n778), .B2(G128), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1142), .B1(new_n836), .B2(new_n799), .C1(new_n365), .C2(new_n776), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n1134), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(G116), .A2(new_n831), .B1(new_n782), .B2(G294), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n205), .B2(new_n766), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n799), .A2(new_n206), .B1(new_n779), .B2(new_n791), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n756), .B1(new_n776), .B2(new_n299), .C1(new_n758), .C2(new_n222), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n823), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n752), .B1(new_n1144), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n738), .B1(new_n259), .B2(new_n820), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n1130), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n1128), .B2(new_n736), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1129), .A2(new_n1154), .ZN(G378));
  AND2_X1   g0955(.A1(new_n927), .A2(new_n1120), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1123), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n895), .A2(new_n908), .A3(KEYINPUT40), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n894), .A2(new_n851), .A3(new_n816), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n901), .B2(new_n913), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1158), .B(G330), .C1(new_n1160), .C2(KEYINPUT40), .ZN(new_n1161));
  XOR2_X1   g0961(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT117), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n312), .A2(new_n875), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n353), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1165), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n352), .B(new_n1167), .C1(new_n316), .C2(new_n321), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1164), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n353), .A2(new_n1165), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1171), .A2(new_n1168), .A3(KEYINPUT117), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1163), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1166), .A2(new_n1169), .A3(new_n1164), .ZN(new_n1174));
  OAI21_X1  g0974(.A(KEYINPUT117), .B1(new_n1171), .B2(new_n1168), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1174), .A2(new_n1175), .A3(new_n1162), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1161), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n892), .A2(new_n893), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1177), .A2(new_n1180), .A3(G330), .A4(new_n1158), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n1179), .A2(new_n921), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n921), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1183));
  OAI21_X1  g0983(.A(KEYINPUT57), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n695), .B1(new_n1157), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1123), .A2(new_n1156), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n921), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1161), .A2(new_n1178), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1177), .B1(new_n903), .B2(G330), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1187), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1179), .A2(new_n921), .A3(new_n1181), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(KEYINPUT57), .B1(new_n1186), .B2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n735), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1178), .A2(new_n750), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1015), .A2(G58), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n756), .A2(new_n285), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1027), .B(new_n1197), .C1(G77), .C2(new_n842), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n770), .A2(G97), .B1(new_n778), .B2(G116), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n763), .A2(new_n206), .B1(new_n781), .B2(new_n791), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n1005), .B2(new_n834), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1196), .A2(new_n1198), .A3(new_n1199), .A4(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT58), .ZN(new_n1203));
  AOI21_X1  g1003(.A(G50), .B1(new_n357), .B2(new_n285), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1202), .A2(new_n1203), .B1(new_n1197), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(G128), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n763), .A2(new_n1206), .B1(new_n766), .B2(new_n836), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n758), .A2(new_n1135), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1208), .A2(KEYINPUT116), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G125), .B2(new_n778), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n797), .A2(G150), .B1(G132), .B2(new_n770), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1207), .B(new_n1212), .C1(KEYINPUT116), .C2(new_n1208), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1015), .A2(G159), .ZN(new_n1216));
  AOI211_X1 g1016(.A(G33), .B(G41), .C1(new_n782), .C2(G124), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1205), .B1(new_n1203), .B2(new_n1202), .C1(new_n1218), .C2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n752), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n820), .A2(new_n276), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1195), .A2(new_n737), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(new_n1194), .A2(KEYINPUT118), .A3(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT118), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n736), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1226), .B1(new_n1227), .B2(new_n1223), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n1185), .A2(new_n1193), .B1(new_n1225), .B2(new_n1228), .ZN(G375));
  OAI22_X1  g1029(.A1(new_n763), .A2(new_n836), .B1(new_n766), .B2(new_n261), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(G159), .B2(new_n842), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n295), .B1(new_n781), .B2(new_n1206), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(G50), .B2(new_n797), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1136), .A2(new_n770), .B1(G132), .B2(new_n778), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1196), .A2(new_n1231), .A3(new_n1233), .A4(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n790), .A2(new_n299), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n295), .B(new_n1059), .C1(G97), .C2(new_n842), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n763), .A2(new_n791), .B1(new_n781), .B2(new_n759), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(G107), .B2(new_n834), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n770), .A2(G116), .B1(new_n778), .B2(G294), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1237), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1235), .B1(new_n1236), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n752), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n738), .B1(new_n202), .B2(new_n820), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1243), .B(new_n1244), .C1(new_n894), .C2(new_n822), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1116), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1246), .A2(new_n735), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1245), .B1(new_n1247), .B2(KEYINPUT119), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(KEYINPUT119), .B2(new_n1247), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n995), .B1(new_n1156), .B2(new_n1116), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1249), .B1(new_n1126), .B2(new_n1250), .ZN(G381));
  XOR2_X1   g1051(.A(G375), .B(KEYINPUT120), .Z(new_n1252));
  NAND4_X1  g1052(.A1(new_n1064), .A2(new_n810), .A3(new_n739), .A4(new_n1066), .ZN(new_n1253));
  OR2_X1    g1053(.A1(G390), .A2(G384), .ZN(new_n1254));
  OR4_X1    g1054(.A1(G387), .A2(G381), .A3(new_n1253), .A4(new_n1254), .ZN(new_n1255));
  OR3_X1    g1055(.A1(new_n1252), .A2(G378), .A3(new_n1255), .ZN(G407));
  INV_X1    g1056(.A(G378), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n676), .A2(G213), .ZN(new_n1258));
  XOR2_X1   g1058(.A(new_n1258), .B(KEYINPUT121), .Z(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(G407), .B(G213), .C1(new_n1252), .C2(new_n1260), .ZN(G409));
  NAND2_X1  g1061(.A1(new_n1227), .A2(new_n1223), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1123), .A2(new_n1156), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1263), .A2(new_n995), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1257), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT57), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1186), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1268), .B(new_n695), .C1(KEYINPUT57), .C2(new_n1263), .ZN(new_n1269));
  OAI21_X1  g1069(.A(KEYINPUT118), .B1(new_n1194), .B2(new_n1224), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1227), .A2(new_n1226), .A3(new_n1223), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1269), .A2(new_n1272), .A3(G378), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1265), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1259), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  AND2_X1   g1077(.A1(new_n1124), .A2(KEYINPUT60), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1156), .A2(new_n1116), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n696), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n1279), .B2(new_n1278), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1281), .A2(G384), .A3(new_n1249), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(G384), .B1(new_n1281), .B2(new_n1249), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1277), .A2(KEYINPUT63), .A3(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1274), .A2(new_n1258), .A3(new_n1285), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT63), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1281), .A2(new_n1249), .ZN(new_n1290));
  INV_X1    g1090(.A(G384), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n1282), .ZN(new_n1293));
  INV_X1    g1093(.A(G2897), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1293), .B1(new_n1294), .B2(new_n1275), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1258), .A2(new_n1294), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1295), .B1(new_n1293), .B2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1274), .A2(new_n1258), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT122), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1004), .A2(new_n1032), .A3(G390), .ZN(new_n1302));
  AOI21_X1  g1102(.A(G390), .B1(new_n1004), .B2(new_n1032), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1301), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(G393), .A2(G396), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1253), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1304), .A2(new_n1307), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1306), .B(new_n1301), .C1(new_n1302), .C2(new_n1303), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1310), .A2(KEYINPUT61), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1286), .A2(new_n1289), .A3(new_n1300), .A4(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1277), .A2(KEYINPUT62), .A3(new_n1285), .ZN(new_n1313));
  XOR2_X1   g1113(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n1314));
  NAND2_X1  g1114(.A1(new_n1287), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1313), .A2(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(KEYINPUT61), .B1(new_n1298), .B2(new_n1276), .ZN(new_n1317));
  AND2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1310), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1312), .B1(new_n1318), .B2(new_n1319), .ZN(G405));
  INV_X1    g1120(.A(KEYINPUT126), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1269), .A2(new_n1272), .A3(G378), .ZN(new_n1322));
  AOI21_X1  g1122(.A(G378), .B1(new_n1269), .B2(new_n1272), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1285), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(G375), .A2(new_n1257), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1325), .A2(new_n1293), .A3(new_n1273), .ZN(new_n1326));
  AOI211_X1 g1126(.A(KEYINPUT125), .B(new_n1310), .C1(new_n1324), .C2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT125), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1324), .A2(new_n1326), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1328), .B1(new_n1329), .B2(new_n1319), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1327), .A2(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1324), .A2(new_n1326), .A3(new_n1310), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT124), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1324), .A2(new_n1326), .A3(new_n1310), .A4(KEYINPUT124), .ZN(new_n1335));
  AND2_X1   g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1321), .B1(new_n1331), .B2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1338));
  OAI211_X1 g1138(.A(new_n1338), .B(KEYINPUT126), .C1(new_n1330), .C2(new_n1327), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1337), .A2(new_n1339), .ZN(G402));
endmodule


