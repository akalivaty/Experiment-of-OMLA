//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n441, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n559,
    new_n561, new_n562, new_n563, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1149, new_n1150, new_n1151;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XNOR2_X1  g015(.A(KEYINPUT66), .B(G57), .ZN(new_n441));
  INV_X1    g016(.A(new_n441), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(new_n441), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT67), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(new_n455), .B2(G567), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n460), .A2(new_n462), .A3(G137), .ZN(new_n463));
  NAND2_X1  g038(.A1(G101), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n460), .A2(new_n462), .A3(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT68), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n460), .A2(new_n462), .A3(new_n469), .A4(G125), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n467), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n465), .B1(new_n471), .B2(G2105), .ZN(G160));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n460), .A2(new_n462), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n477), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT70), .Z(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n474), .A2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n459), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  NOR2_X1   g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n490), .A2(KEYINPUT71), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(new_n475), .B2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(new_n491), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n477), .A2(G126), .A3(G2105), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n460), .A2(new_n462), .A3(G138), .A4(new_n475), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n477), .A2(KEYINPUT4), .A3(G138), .A4(new_n475), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n497), .A2(new_n498), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT73), .B1(new_n505), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(new_n508), .A3(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n505), .A2(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G88), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G50), .ZN(new_n518));
  XOR2_X1   g093(.A(new_n518), .B(KEYINPUT72), .Z(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n512), .A2(G62), .ZN(new_n521));
  NAND2_X1  g096(.A1(G75), .A2(G543), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n523), .A2(KEYINPUT74), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n523), .A2(KEYINPUT74), .ZN(new_n525));
  OAI211_X1 g100(.A(new_n515), .B(new_n519), .C1(new_n524), .C2(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND2_X1  g102(.A1(new_n514), .A2(G89), .ZN(new_n528));
  XOR2_X1   g103(.A(KEYINPUT75), .B(KEYINPUT7), .Z(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n529), .B(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(G63), .A2(G651), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n512), .A2(new_n532), .B1(new_n517), .B2(G51), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n528), .A2(new_n531), .A3(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  AOI22_X1  g110(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n520), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT76), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n537), .B(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n514), .A2(G90), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n517), .A2(G52), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(new_n517), .A2(G43), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n512), .A2(new_n513), .ZN(new_n546));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n510), .A2(new_n511), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G651), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(KEYINPUT77), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(KEYINPUT77), .ZN(new_n555));
  AOI211_X1 g130(.A(new_n545), .B(new_n548), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(new_n557));
  XOR2_X1   g132(.A(new_n557), .B(KEYINPUT78), .Z(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(G176));
  XOR2_X1   g135(.A(KEYINPUT79), .B(KEYINPUT8), .Z(new_n561));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n559), .A2(new_n563), .ZN(G188));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n565), .A2(KEYINPUT80), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n517), .A2(G53), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(KEYINPUT80), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT81), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n550), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n514), .A2(G91), .B1(G651), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n569), .A2(new_n574), .ZN(G299));
  OAI21_X1  g150(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n517), .A2(G49), .ZN(new_n577));
  INV_X1    g152(.A(G87), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n576), .B(new_n577), .C1(new_n578), .C2(new_n546), .ZN(G288));
  NAND2_X1  g154(.A1(new_n514), .A2(G86), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n550), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n583), .A2(G651), .B1(new_n517), .B2(G48), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n580), .A2(new_n584), .ZN(G305));
  AOI22_X1  g160(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(new_n520), .ZN(new_n587));
  INV_X1    g162(.A(G85), .ZN(new_n588));
  INV_X1    g163(.A(G47), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n546), .A2(new_n588), .B1(new_n589), .B2(new_n516), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(new_n514), .A2(G92), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n517), .A2(G54), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n512), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(new_n520), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(G171), .B2(new_n600), .ZN(G284));
  OAI21_X1  g177(.A(new_n601), .B1(G171), .B2(new_n600), .ZN(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  INV_X1    g179(.A(G299), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G280));
  XNOR2_X1  g181(.A(G280), .B(KEYINPUT82), .ZN(G297));
  AND3_X1   g182(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(new_n608));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G860), .ZN(G148));
  NOR2_X1   g185(.A1(new_n599), .A2(G559), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n611), .A2(new_n600), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n556), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(KEYINPUT83), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(KEYINPUT83), .B2(new_n612), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g191(.A1(new_n485), .A2(G135), .ZN(new_n617));
  OAI21_X1  g192(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT86), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n620), .B(new_n621), .C1(G111), .C2(new_n475), .ZN(new_n622));
  INV_X1    g197(.A(G123), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n617), .B(new_n622), .C1(new_n479), .C2(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(G2096), .Z(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n626));
  NOR3_X1   g201(.A1(new_n461), .A2(new_n459), .A3(G2105), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  AND2_X1   g204(.A1(KEYINPUT85), .A2(G2100), .ZN(new_n630));
  NOR2_X1   g205(.A1(KEYINPUT85), .A2(G2100), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n625), .B(new_n632), .C1(new_n629), .C2(new_n630), .ZN(G156));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XOR2_X1   g210(.A(G2443), .B(G2446), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XOR2_X1   g216(.A(KEYINPUT15), .B(G2435), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(KEYINPUT14), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n639), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(G14), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(G401));
  XOR2_X1   g222(.A(G2067), .B(G2678), .Z(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT87), .Z(new_n649));
  XOR2_X1   g224(.A(G2072), .B(G2078), .Z(new_n650));
  NOR2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT88), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT18), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n652), .B1(new_n649), .B2(new_n650), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n650), .B(KEYINPUT17), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n656), .B1(new_n649), .B2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT89), .Z(new_n660));
  NAND3_X1  g235(.A1(new_n658), .A2(new_n652), .A3(new_n649), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n655), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2096), .B(G2100), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(G227));
  INV_X1    g240(.A(KEYINPUT20), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1961), .B(G1966), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT90), .ZN(new_n668));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n666), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n668), .A2(new_n669), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n675), .A2(new_n672), .A3(new_n670), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n670), .A2(new_n666), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n677), .A2(new_n674), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n673), .B(new_n676), .C1(new_n678), .C2(new_n672), .ZN(new_n679));
  XOR2_X1   g254(.A(G1991), .B(G1996), .Z(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT91), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n683), .B(new_n685), .ZN(G229));
  INV_X1    g261(.A(G29), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G32), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n485), .A2(G141), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT99), .Z(new_n690));
  NAND2_X1  g265(.A1(new_n480), .A2(G129), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n475), .A2(G105), .A3(G2104), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT100), .ZN(new_n693));
  NAND3_X1  g268(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT26), .Z(new_n695));
  NAND4_X1  g270(.A1(new_n690), .A2(new_n691), .A3(new_n693), .A4(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n688), .B1(new_n697), .B2(new_n687), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT101), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT27), .B(G1996), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G19), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(new_n556), .B2(new_n702), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(G1341), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n702), .A2(G4), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(new_n608), .B2(new_n702), .ZN(new_n707));
  INV_X1    g282(.A(G1348), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n687), .A2(G26), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n480), .A2(G128), .B1(G140), .B2(new_n485), .ZN(new_n711));
  OR2_X1    g286(.A1(G104), .A2(G2105), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n712), .B(G2104), .C1(G116), .C2(new_n475), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT96), .Z(new_n714));
  NAND2_X1  g289(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n710), .B1(new_n715), .B2(G29), .ZN(new_n716));
  MUX2_X1   g291(.A(new_n710), .B(new_n716), .S(KEYINPUT28), .Z(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT97), .B(G2067), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n709), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(G2090), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n687), .A2(G35), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n487), .B2(G29), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT29), .ZN(new_n724));
  AOI211_X1 g299(.A(new_n705), .B(new_n720), .C1(new_n721), .C2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n702), .A2(G20), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT102), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT23), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n605), .B2(new_n702), .ZN(new_n729));
  INV_X1    g304(.A(G1956), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n724), .B2(new_n721), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT103), .ZN(new_n733));
  INV_X1    g308(.A(G28), .ZN(new_n734));
  AOI21_X1  g309(.A(G29), .B1(new_n734), .B2(KEYINPUT30), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(KEYINPUT30), .B2(new_n734), .ZN(new_n736));
  NAND2_X1  g311(.A1(G168), .A2(G16), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G16), .B2(G21), .ZN(new_n738));
  INV_X1    g313(.A(G1966), .ZN(new_n739));
  OAI221_X1 g314(.A(new_n736), .B1(new_n687), .B2(new_n624), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(G29), .A2(G33), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT25), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n485), .A2(G139), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n743), .B(new_n744), .C1(new_n475), .C2(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT98), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n741), .B1(new_n748), .B2(G29), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n740), .B1(G2072), .B2(new_n749), .ZN(new_n750));
  OR2_X1    g325(.A1(KEYINPUT24), .A2(G34), .ZN(new_n751));
  NAND2_X1  g326(.A1(KEYINPUT24), .A2(G34), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n751), .A2(new_n687), .A3(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G160), .B2(new_n687), .ZN(new_n754));
  OAI22_X1  g329(.A1(new_n749), .A2(G2072), .B1(G2084), .B2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G2084), .B2(new_n754), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n687), .A2(G27), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G164), .B2(new_n687), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2078), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n738), .B2(new_n739), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n750), .A2(new_n756), .A3(new_n760), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT31), .B(G11), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n702), .A2(G5), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G171), .B2(new_n702), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G1961), .ZN(new_n765));
  NOR3_X1   g340(.A1(new_n761), .A2(new_n762), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n725), .A2(new_n733), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n485), .A2(G131), .ZN(new_n768));
  NOR2_X1   g343(.A1(G95), .A2(G2105), .ZN(new_n769));
  OAI21_X1  g344(.A(G2104), .B1(new_n475), .B2(G107), .ZN(new_n770));
  INV_X1    g345(.A(G119), .ZN(new_n771));
  OAI221_X1 g346(.A(new_n768), .B1(new_n769), .B2(new_n770), .C1(new_n479), .C2(new_n771), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT92), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G29), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G25), .B2(G29), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT35), .B(G1991), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT93), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n775), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n702), .A2(G6), .ZN(new_n779));
  INV_X1    g354(.A(G305), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n780), .B2(new_n702), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT94), .Z(new_n782));
  XOR2_X1   g357(.A(KEYINPUT32), .B(G1981), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT34), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n702), .A2(G22), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G166), .B2(new_n702), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(G1971), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(G1971), .ZN(new_n789));
  NOR2_X1   g364(.A1(G16), .A2(G23), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT95), .ZN(new_n791));
  NAND2_X1  g366(.A1(G288), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n514), .A2(G87), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n793), .A2(KEYINPUT95), .A3(new_n576), .A4(new_n577), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n790), .B1(new_n795), .B2(G16), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT33), .B(G1976), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n788), .A2(new_n789), .A3(new_n798), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n784), .A2(new_n785), .A3(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n785), .B1(new_n784), .B2(new_n799), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n778), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT36), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n702), .A2(G24), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n591), .B2(new_n702), .ZN(new_n806));
  INV_X1    g381(.A(G1986), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n803), .A2(new_n804), .A3(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n778), .ZN(new_n810));
  INV_X1    g385(.A(new_n802), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n808), .B(new_n810), .C1(new_n811), .C2(new_n800), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(KEYINPUT36), .ZN(new_n813));
  AOI211_X1 g388(.A(new_n701), .B(new_n767), .C1(new_n809), .C2(new_n813), .ZN(G311));
  AOI21_X1  g389(.A(new_n767), .B1(new_n809), .B2(new_n813), .ZN(new_n815));
  INV_X1    g390(.A(new_n701), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(G150));
  AOI22_X1  g392(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n818), .A2(new_n520), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n512), .A2(G93), .A3(new_n513), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n517), .A2(G55), .ZN(new_n821));
  AND3_X1   g396(.A1(new_n820), .A2(KEYINPUT104), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(KEYINPUT104), .B1(new_n820), .B2(new_n821), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n819), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(G860), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT37), .Z(new_n826));
  NOR2_X1   g401(.A1(new_n599), .A2(new_n609), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n824), .A2(KEYINPUT105), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT105), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n819), .B(new_n831), .C1(new_n822), .C2(new_n823), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n556), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n556), .B1(new_n830), .B2(new_n832), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n829), .B(new_n836), .Z(new_n837));
  OAI21_X1  g412(.A(new_n826), .B1(new_n837), .B2(G860), .ZN(G145));
  XOR2_X1   g413(.A(new_n487), .B(G160), .Z(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n748), .A2(new_n503), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n747), .A2(G164), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n485), .A2(G142), .ZN(new_n843));
  NOR2_X1   g418(.A1(G106), .A2(G2105), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(new_n475), .B2(G118), .ZN(new_n845));
  INV_X1    g420(.A(G130), .ZN(new_n846));
  OAI221_X1 g421(.A(new_n843), .B1(new_n844), .B2(new_n845), .C1(new_n479), .C2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT106), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n841), .A2(new_n842), .A3(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n715), .B(new_n772), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n848), .B1(new_n841), .B2(new_n842), .ZN(new_n853));
  NOR3_X1   g428(.A1(new_n850), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n841), .A2(new_n842), .ZN(new_n855));
  INV_X1    g430(.A(new_n848), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n851), .B1(new_n857), .B2(new_n849), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n697), .B1(new_n854), .B2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n624), .B(new_n628), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n852), .B1(new_n850), .B2(new_n853), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n857), .A2(new_n851), .A3(new_n849), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n861), .A2(new_n696), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n859), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n860), .B1(new_n859), .B2(new_n863), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n840), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(G37), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n859), .A2(new_n863), .ZN(new_n869));
  INV_X1    g444(.A(new_n860), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n871), .A2(new_n839), .A3(new_n864), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n867), .A2(new_n868), .A3(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g449(.A1(new_n824), .A2(new_n600), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n608), .A2(new_n605), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n599), .A2(G299), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n876), .A2(KEYINPUT41), .A3(new_n877), .ZN(new_n880));
  AOI21_X1  g455(.A(KEYINPUT41), .B1(new_n876), .B2(new_n877), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n836), .B(new_n611), .ZN(new_n883));
  MUX2_X1   g458(.A(new_n879), .B(new_n882), .S(new_n883), .Z(new_n884));
  NAND2_X1  g459(.A1(new_n795), .A2(new_n591), .ZN(new_n885));
  NAND3_X1  g460(.A1(G290), .A2(new_n792), .A3(new_n794), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n887), .A2(new_n780), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n780), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n889), .A2(G166), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(G166), .B1(new_n889), .B2(new_n890), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OR2_X1    g468(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n894));
  NAND2_X1  g469(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(new_n895), .B2(new_n893), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n884), .B(new_n897), .Z(new_n898));
  OAI21_X1  g473(.A(new_n875), .B1(new_n898), .B2(new_n600), .ZN(G295));
  OAI21_X1  g474(.A(new_n875), .B1(new_n898), .B2(new_n600), .ZN(G331));
  NOR2_X1   g475(.A1(G168), .A2(KEYINPUT108), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n545), .B1(new_n554), .B2(new_n555), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(new_n547), .B2(new_n546), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n824), .A2(KEYINPUT105), .ZN(new_n905));
  INV_X1    g480(.A(new_n832), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(G168), .A2(KEYINPUT108), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n908), .A2(new_n539), .A3(new_n540), .A4(new_n541), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n907), .A2(new_n833), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n909), .B1(new_n907), .B2(new_n833), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n902), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI211_X1 g487(.A(G171), .B(new_n908), .C1(new_n834), .C2(new_n835), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n907), .A2(new_n833), .A3(new_n909), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(new_n914), .A3(new_n901), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n912), .A2(new_n915), .A3(new_n882), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n878), .B1(new_n912), .B2(new_n915), .ZN(new_n917));
  OAI22_X1  g492(.A1(new_n916), .A2(new_n917), .B1(new_n891), .B2(new_n892), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n912), .A2(new_n915), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n879), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n912), .A2(new_n915), .A3(new_n882), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(new_n893), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n918), .A2(new_n922), .A3(new_n868), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT43), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n918), .A2(new_n922), .A3(new_n925), .A4(new_n868), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n924), .A2(KEYINPUT44), .A3(new_n926), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(G397));
  INV_X1    g506(.A(G1384), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT71), .B1(new_n490), .B2(new_n492), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n495), .A2(new_n494), .A3(new_n491), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n498), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n501), .A2(new_n502), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT109), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT45), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n471), .A2(G2105), .ZN(new_n941));
  INV_X1    g516(.A(new_n465), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n941), .A2(G40), .A3(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n945), .A2(G1996), .ZN(new_n946));
  OR2_X1    g521(.A1(new_n946), .A2(KEYINPUT46), .ZN(new_n947));
  INV_X1    g522(.A(G2067), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n711), .A2(new_n948), .A3(new_n714), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n715), .A2(G2067), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n697), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n944), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n946), .A2(KEYINPUT46), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n947), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n954), .B(KEYINPUT47), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n944), .A2(new_n807), .A3(new_n591), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n956), .B(KEYINPUT48), .ZN(new_n957));
  INV_X1    g532(.A(G1996), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n696), .B(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(new_n949), .A3(new_n950), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n772), .B(new_n776), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n957), .B1(new_n945), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n776), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n773), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n949), .B1(new_n960), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n944), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n955), .A2(new_n963), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT126), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n968), .B(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n937), .A2(new_n939), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT110), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n937), .A2(new_n973), .A3(new_n939), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G40), .ZN(new_n976));
  AOI211_X1 g551(.A(new_n976), .B(new_n465), .C1(new_n471), .C2(G2105), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(new_n939), .B2(new_n937), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n975), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT111), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n978), .B1(new_n972), .B2(new_n974), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(G1971), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n937), .A2(KEYINPUT50), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n503), .B2(new_n932), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n989), .A2(new_n943), .A3(KEYINPUT116), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT116), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n937), .A2(KEYINPUT50), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n991), .B1(new_n992), .B2(new_n977), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n987), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n994), .A2(G2090), .ZN(new_n995));
  OAI21_X1  g570(.A(G8), .B1(new_n985), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n997));
  AND3_X1   g572(.A1(G303), .A2(new_n997), .A3(G8), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n997), .B1(G303), .B2(G8), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n996), .A2(new_n1001), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n986), .A2(new_n943), .A3(new_n989), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n1003), .A2(new_n721), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1000), .B(G8), .C1(new_n985), .C2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1981), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT113), .B(G86), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n514), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1006), .B1(new_n1009), .B2(new_n584), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT49), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(G305), .A2(G1981), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1013), .B1(new_n1015), .B2(new_n1010), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1012), .A2(KEYINPUT114), .A3(new_n1013), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1014), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n943), .A2(new_n937), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1022), .A2(G8), .ZN(new_n1023));
  INV_X1    g598(.A(G288), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1024), .A2(G1976), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT52), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT112), .B1(new_n795), .B2(G1976), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n1023), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1027), .B(new_n1023), .C1(KEYINPUT52), .C2(new_n1025), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n1020), .A2(new_n1023), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1002), .A2(new_n1005), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT62), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n979), .A2(new_n971), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n739), .ZN(new_n1035));
  INV_X1    g610(.A(G2084), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1003), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1035), .A2(G168), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(G8), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT51), .ZN(new_n1040));
  AOI21_X1  g615(.A(G168), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT51), .ZN(new_n1042));
  OAI211_X1 g617(.A(G8), .B(new_n1038), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1033), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1032), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1040), .A2(new_n1043), .A3(new_n1033), .ZN(new_n1046));
  INV_X1    g621(.A(G2078), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n981), .A2(new_n1047), .A3(new_n984), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OR2_X1    g625(.A1(new_n1003), .A2(KEYINPUT119), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1003), .A2(KEYINPUT119), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT123), .B(G1961), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1047), .A2(KEYINPUT53), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1050), .B(new_n1054), .C1(new_n1034), .C2(new_n1055), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1046), .A2(new_n1056), .A3(G171), .ZN(new_n1057));
  AOI21_X1  g632(.A(G1976), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n1024), .ZN(new_n1059));
  XNOR2_X1  g634(.A(new_n1007), .B(KEYINPUT115), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  AOI22_X1  g636(.A1(new_n1045), .A2(new_n1057), .B1(new_n1023), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1005), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n1031), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT63), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1039), .A2(G286), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1065), .B1(new_n1032), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(G8), .B1(new_n985), .B2(new_n1004), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1065), .B1(new_n1069), .B2(new_n1001), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1070), .A2(new_n1005), .A3(new_n1031), .A4(new_n1066), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1062), .A2(new_n1064), .A3(new_n1072), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT58), .B(G1341), .Z(new_n1074));
  AOI22_X1  g649(.A1(new_n982), .A2(new_n958), .B1(new_n1022), .B2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1075), .A2(new_n904), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT59), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1076), .B(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT56), .B(G2072), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n982), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1083), .B1(new_n994), .B2(new_n730), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n992), .A2(new_n991), .A3(new_n977), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT116), .B1(new_n989), .B2(new_n943), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n986), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1087), .A2(KEYINPUT117), .A3(G1956), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1082), .B1(new_n1084), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n605), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1093));
  NAND2_X1  g668(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n1094));
  NAND3_X1  g669(.A1(G299), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1089), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n994), .A2(new_n1083), .A3(new_n730), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT117), .B1(new_n1087), .B2(G1956), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1081), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1096), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1097), .A2(KEYINPUT61), .A3(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1051), .A2(new_n708), .A3(new_n1052), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1021), .A2(new_n948), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n599), .A2(KEYINPUT60), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1104), .A2(new_n599), .A3(new_n1105), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n599), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT60), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AND4_X1   g685(.A1(new_n1079), .A2(new_n1103), .A3(new_n1107), .A4(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(new_n1089), .B2(new_n1096), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n1100), .A2(KEYINPUT121), .A3(new_n1101), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1102), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT61), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT122), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AOI211_X1 g692(.A(new_n1096), .B(new_n1081), .C1(new_n1099), .C2(new_n1098), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1089), .A2(new_n1112), .A3(new_n1096), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT121), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1121), .A2(new_n1122), .A3(KEYINPUT61), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1111), .B1(new_n1117), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1097), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1125), .B1(new_n1109), .B2(new_n1102), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(G301), .B(KEYINPUT54), .ZN(new_n1128));
  AOI211_X1 g703(.A(new_n1055), .B(new_n978), .C1(new_n938), .C2(new_n939), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1054), .A2(KEYINPUT124), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1054), .A2(KEYINPUT124), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1130), .B(new_n1050), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1133), .A2(new_n1005), .A3(new_n1031), .A4(new_n1002), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1056), .A2(new_n1128), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT125), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1032), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1056), .A2(new_n1128), .B1(new_n1043), .B2(new_n1040), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT125), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .A4(new_n1133), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1138), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1073), .B1(new_n1127), .B2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n591), .B(G1986), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n945), .B1(new_n962), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n970), .B1(new_n1144), .B2(new_n1146), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g722(.A1(new_n873), .A2(new_n664), .ZN(new_n1149));
  NAND2_X1  g723(.A1(new_n646), .A2(G319), .ZN(new_n1150));
  NOR2_X1   g724(.A1(G229), .A2(new_n1150), .ZN(new_n1151));
  AND3_X1   g725(.A1(new_n1149), .A2(new_n927), .A3(new_n1151), .ZN(G308));
  NAND3_X1  g726(.A1(new_n1149), .A2(new_n927), .A3(new_n1151), .ZN(G225));
endmodule


