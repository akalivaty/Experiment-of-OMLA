

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734;

  NOR2_X1 U375 ( .A1(n612), .A2(n699), .ZN(n613) );
  NOR2_X2 U376 ( .A1(n734), .A2(n733), .ZN(n526) );
  XOR2_X2 U377 ( .A(KEYINPUT42), .B(n517), .Z(n734) );
  OR2_X2 U378 ( .A1(n516), .A2(n678), .ZN(n517) );
  XNOR2_X2 U379 ( .A(n590), .B(n497), .ZN(n583) );
  INV_X2 U380 ( .A(G953), .ZN(n603) );
  AND2_X1 U381 ( .A1(n691), .A2(n618), .ZN(n692) );
  XOR2_X1 U382 ( .A(n515), .B(n514), .Z(n678) );
  NOR2_X1 U383 ( .A1(n668), .A2(n665), .ZN(n515) );
  NOR2_X1 U384 ( .A1(n496), .A2(G902), .ZN(n390) );
  XNOR2_X1 U385 ( .A(n688), .B(KEYINPUT59), .ZN(n689) );
  XNOR2_X1 U386 ( .A(n411), .B(n429), .ZN(n365) );
  XNOR2_X1 U387 ( .A(n413), .B(n412), .ZN(n411) );
  XNOR2_X1 U388 ( .A(n406), .B(G140), .ZN(n481) );
  NOR2_X1 U389 ( .A1(n646), .A2(n575), .ZN(n582) );
  XNOR2_X1 U390 ( .A(G146), .B(G125), .ZN(n450) );
  XNOR2_X1 U391 ( .A(n434), .B(n705), .ZN(n444) );
  XNOR2_X1 U392 ( .A(n432), .B(n431), .ZN(n434) );
  XNOR2_X1 U393 ( .A(n371), .B(n370), .ZN(n408) );
  INV_X1 U394 ( .A(KEYINPUT48), .ZN(n370) );
  XNOR2_X1 U395 ( .A(n730), .B(n373), .ZN(n372) );
  OR2_X1 U396 ( .A1(n614), .A2(G902), .ZN(n392) );
  XNOR2_X1 U397 ( .A(n570), .B(n569), .ZN(n575) );
  XNOR2_X1 U398 ( .A(KEYINPUT64), .B(KEYINPUT22), .ZN(n569) );
  XNOR2_X1 U399 ( .A(n436), .B(n383), .ZN(n382) );
  INV_X1 U400 ( .A(KEYINPUT16), .ZN(n383) );
  XNOR2_X1 U401 ( .A(n499), .B(KEYINPUT101), .ZN(n544) );
  XNOR2_X1 U402 ( .A(n481), .B(n405), .ZN(n442) );
  INV_X1 U403 ( .A(G107), .ZN(n405) );
  NAND2_X1 U404 ( .A1(n404), .A2(n621), .ZN(n403) );
  NAND2_X1 U405 ( .A1(n354), .A2(n527), .ZN(n404) );
  NOR2_X1 U406 ( .A1(G953), .A2(G237), .ZN(n419) );
  INV_X1 U407 ( .A(n644), .ZN(n409) );
  NAND2_X1 U408 ( .A1(n531), .A2(n532), .ZN(n665) );
  NAND2_X1 U409 ( .A1(n663), .A2(n662), .ZN(n668) );
  NAND2_X1 U410 ( .A1(n646), .A2(n647), .ZN(n589) );
  XNOR2_X1 U411 ( .A(n657), .B(n506), .ZN(n518) );
  XNOR2_X1 U412 ( .A(n417), .B(n416), .ZN(n652) );
  XNOR2_X1 U413 ( .A(n485), .B(KEYINPUT25), .ZN(n416) );
  OR2_X1 U414 ( .A1(n697), .A2(G902), .ZN(n417) );
  XNOR2_X1 U415 ( .A(n426), .B(n427), .ZN(n496) );
  NAND2_X1 U416 ( .A1(n408), .A2(n368), .ZN(n719) );
  XNOR2_X1 U417 ( .A(G143), .B(G104), .ZN(n455) );
  XNOR2_X1 U418 ( .A(G122), .B(G140), .ZN(n451) );
  XOR2_X1 U419 ( .A(KEYINPUT94), .B(KEYINPUT12), .Z(n448) );
  XNOR2_X1 U420 ( .A(n365), .B(n410), .ZN(n435) );
  NOR2_X1 U421 ( .A1(n575), .A2(n574), .ZN(n576) );
  INV_X1 U422 ( .A(KEYINPUT6), .ZN(n497) );
  INV_X1 U423 ( .A(n617), .ZN(n380) );
  NAND2_X1 U424 ( .A1(n395), .A2(n362), .ZN(n393) );
  INV_X1 U425 ( .A(KEYINPUT81), .ZN(n373) );
  AND2_X1 U426 ( .A1(n540), .A2(n541), .ZN(n374) );
  XOR2_X1 U427 ( .A(G137), .B(G116), .Z(n422) );
  XNOR2_X1 U428 ( .A(n715), .B(G146), .ZN(n446) );
  XNOR2_X1 U429 ( .A(n467), .B(n425), .ZN(n715) );
  XNOR2_X1 U430 ( .A(KEYINPUT4), .B(G131), .ZN(n425) );
  XNOR2_X1 U431 ( .A(n384), .B(G119), .ZN(n436) );
  XNOR2_X1 U432 ( .A(G113), .B(KEYINPUT3), .ZN(n384) );
  INV_X1 U433 ( .A(KEYINPUT72), .ZN(n400) );
  INV_X1 U434 ( .A(G137), .ZN(n406) );
  XNOR2_X1 U435 ( .A(n430), .B(G134), .ZN(n467) );
  XNOR2_X1 U436 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n428) );
  INV_X1 U437 ( .A(KEYINPUT4), .ZN(n412) );
  INV_X1 U438 ( .A(KEYINPUT79), .ZN(n387) );
  NAND2_X1 U439 ( .A1(G234), .A2(G237), .ZN(n486) );
  NOR2_X1 U440 ( .A1(n652), .A2(n651), .ZN(n647) );
  XNOR2_X1 U441 ( .A(G104), .B(KEYINPUT74), .ZN(n433) );
  INV_X1 U442 ( .A(n467), .ZN(n376) );
  XOR2_X1 U443 ( .A(G116), .B(G107), .Z(n437) );
  AND2_X1 U444 ( .A1(n617), .A2(G469), .ZN(n396) );
  XNOR2_X1 U445 ( .A(n391), .B(KEYINPUT39), .ZN(n548) );
  XNOR2_X1 U446 ( .A(n364), .B(n551), .ZN(n679) );
  XNOR2_X1 U447 ( .A(n542), .B(n361), .ZN(n559) );
  XNOR2_X1 U448 ( .A(n415), .B(n414), .ZN(n531) );
  INV_X1 U449 ( .A(G478), .ZN(n414) );
  OR2_X1 U450 ( .A1(n694), .A2(G902), .ZN(n415) );
  INV_X1 U451 ( .A(G472), .ZN(n389) );
  AND2_X1 U452 ( .A1(n531), .A2(n513), .ZN(n367) );
  XNOR2_X1 U453 ( .A(n377), .B(n375), .ZN(n694) );
  XNOR2_X1 U454 ( .A(n465), .B(n378), .ZN(n377) );
  XNOR2_X1 U455 ( .A(n470), .B(n376), .ZN(n375) );
  XNOR2_X1 U456 ( .A(n466), .B(KEYINPUT96), .ZN(n378) );
  XNOR2_X1 U457 ( .A(n460), .B(n459), .ZN(n688) );
  XNOR2_X1 U458 ( .A(n458), .B(n457), .ZN(n459) );
  AND2_X1 U459 ( .A1(n369), .A2(n512), .ZN(n644) );
  XNOR2_X1 U460 ( .A(n547), .B(KEYINPUT106), .ZN(n730) );
  XNOR2_X1 U461 ( .A(n545), .B(KEYINPUT36), .ZN(n546) );
  XNOR2_X1 U462 ( .A(KEYINPUT76), .B(KEYINPUT32), .ZN(n578) );
  XNOR2_X1 U463 ( .A(n386), .B(n385), .ZN(n641) );
  XNOR2_X1 U464 ( .A(KEYINPUT31), .B(KEYINPUT90), .ZN(n385) );
  NOR2_X1 U465 ( .A1(n397), .A2(n393), .ZN(n620) );
  XNOR2_X1 U466 ( .A(n610), .B(n611), .ZN(n612) );
  AND2_X1 U467 ( .A1(n523), .A2(n663), .ZN(n352) );
  XOR2_X1 U468 ( .A(KEYINPUT69), .B(G469), .Z(n353) );
  XNOR2_X1 U469 ( .A(KEYINPUT91), .B(n592), .ZN(n354) );
  AND2_X1 U470 ( .A1(n548), .A2(n367), .ZN(n355) );
  XNOR2_X1 U471 ( .A(n512), .B(KEYINPUT38), .ZN(n663) );
  AND2_X1 U472 ( .A1(n700), .A2(n387), .ZN(n356) );
  AND2_X1 U473 ( .A1(n581), .A2(KEYINPUT44), .ZN(n357) );
  AND2_X1 U474 ( .A1(n366), .A2(G475), .ZN(n358) );
  AND2_X1 U475 ( .A1(n366), .A2(G472), .ZN(n359) );
  AND2_X1 U476 ( .A1(n366), .A2(G210), .ZN(n360) );
  XOR2_X1 U477 ( .A(KEYINPUT65), .B(KEYINPUT19), .Z(n361) );
  XNOR2_X1 U478 ( .A(n367), .B(n471), .ZN(n637) );
  AND2_X1 U479 ( .A1(n394), .A2(n618), .ZN(n362) );
  XNOR2_X1 U480 ( .A(KEYINPUT43), .B(KEYINPUT104), .ZN(n363) );
  NOR2_X1 U481 ( .A1(G952), .A2(n603), .ZN(n699) );
  NAND2_X1 U482 ( .A1(n550), .A2(n549), .ZN(n364) );
  NAND2_X1 U483 ( .A1(n402), .A2(n399), .ZN(n398) );
  NAND2_X1 U484 ( .A1(n559), .A2(n560), .ZN(n562) );
  NOR2_X1 U485 ( .A1(n403), .A2(n357), .ZN(n402) );
  XNOR2_X1 U486 ( .A(n401), .B(n400), .ZN(n399) );
  NOR2_X1 U487 ( .A1(n539), .A2(n538), .ZN(n540) );
  INV_X1 U488 ( .A(n719), .ZN(n388) );
  XNOR2_X1 U489 ( .A(n482), .B(n714), .ZN(n697) );
  NAND2_X1 U490 ( .A1(n600), .A2(n366), .ZN(n381) );
  NAND2_X1 U491 ( .A1(n682), .A2(n366), .ZN(n683) );
  NAND2_X2 U492 ( .A1(n593), .A2(n594), .ZN(n366) );
  NOR2_X1 U493 ( .A1(n640), .A2(n367), .ZN(n667) );
  NOR2_X1 U494 ( .A1(n644), .A2(n407), .ZN(n368) );
  XNOR2_X1 U495 ( .A(n504), .B(n363), .ZN(n369) );
  NAND2_X1 U496 ( .A1(n374), .A2(n372), .ZN(n371) );
  NAND2_X1 U497 ( .A1(n358), .A2(n600), .ZN(n690) );
  INV_X1 U498 ( .A(n381), .ZN(n379) );
  NAND2_X1 U499 ( .A1(n359), .A2(n600), .ZN(n601) );
  NAND2_X1 U500 ( .A1(n360), .A2(n600), .ZN(n610) );
  NAND2_X1 U501 ( .A1(n379), .A2(n396), .ZN(n395) );
  NAND2_X1 U502 ( .A1(n379), .A2(G478), .ZN(n693) );
  NAND2_X1 U503 ( .A1(n379), .A2(G217), .ZN(n696) );
  AND2_X1 U504 ( .A1(n381), .A2(n380), .ZN(n397) );
  XNOR2_X1 U505 ( .A(n465), .B(n382), .ZN(n707) );
  INV_X1 U506 ( .A(n559), .ZN(n558) );
  NAND2_X1 U507 ( .A1(n505), .A2(n662), .ZN(n542) );
  XNOR2_X1 U508 ( .A(n440), .B(n439), .ZN(n505) );
  NOR2_X1 U509 ( .A1(n624), .A2(n641), .ZN(n592) );
  NAND2_X1 U510 ( .A1(n591), .A2(n659), .ZN(n386) );
  XNOR2_X2 U511 ( .A(G143), .B(G128), .ZN(n430) );
  NAND2_X1 U512 ( .A1(n388), .A2(n356), .ZN(n593) );
  XNOR2_X2 U513 ( .A(n390), .B(n389), .ZN(n657) );
  NAND2_X1 U514 ( .A1(n524), .A2(n523), .ZN(n534) );
  NAND2_X1 U515 ( .A1(n524), .A2(n352), .ZN(n391) );
  XNOR2_X2 U516 ( .A(n521), .B(KEYINPUT1), .ZN(n646) );
  XNOR2_X2 U517 ( .A(n392), .B(n353), .ZN(n521) );
  OR2_X1 U518 ( .A1(n617), .A2(G469), .ZN(n394) );
  XNOR2_X2 U519 ( .A(n398), .B(KEYINPUT45), .ZN(n700) );
  NOR2_X2 U520 ( .A1(n581), .A2(KEYINPUT44), .ZN(n401) );
  INV_X1 U521 ( .A(n643), .ZN(n407) );
  AND2_X1 U522 ( .A1(n409), .A2(n408), .ZN(n597) );
  XNOR2_X1 U523 ( .A(n430), .B(n428), .ZN(n410) );
  NAND2_X1 U524 ( .A1(n603), .A2(G224), .ZN(n413) );
  NAND2_X1 U525 ( .A1(n546), .A2(n646), .ZN(n547) );
  INV_X1 U526 ( .A(n657), .ZN(n590) );
  XNOR2_X1 U527 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U528 ( .A(n477), .B(n476), .ZN(n479) );
  AND2_X1 U529 ( .A1(G221), .A2(n478), .ZN(n418) );
  INV_X1 U530 ( .A(n450), .ZN(n429) );
  XNOR2_X1 U531 ( .A(n436), .B(n422), .ZN(n423) );
  INV_X1 U532 ( .A(KEYINPUT23), .ZN(n474) );
  XNOR2_X1 U533 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U534 ( .A(n424), .B(n423), .ZN(n427) );
  INV_X1 U535 ( .A(KEYINPUT97), .ZN(n506) );
  XNOR2_X1 U536 ( .A(n479), .B(n418), .ZN(n482) );
  INV_X1 U537 ( .A(n699), .ZN(n618) );
  XNOR2_X1 U538 ( .A(n579), .B(n578), .ZN(n729) );
  XOR2_X2 U539 ( .A(KEYINPUT66), .B(G101), .Z(n432) );
  XOR2_X1 U540 ( .A(n432), .B(KEYINPUT5), .Z(n421) );
  XOR2_X1 U541 ( .A(KEYINPUT75), .B(n419), .Z(n454) );
  NAND2_X1 U542 ( .A1(n454), .A2(G210), .ZN(n420) );
  XNOR2_X1 U543 ( .A(n421), .B(n420), .ZN(n424) );
  INV_X1 U544 ( .A(n446), .ZN(n426) );
  XNOR2_X1 U545 ( .A(n496), .B(KEYINPUT62), .ZN(n602) );
  XOR2_X1 U546 ( .A(G902), .B(KEYINPUT15), .Z(n483) );
  XOR2_X1 U547 ( .A(KEYINPUT71), .B(KEYINPUT70), .Z(n431) );
  XNOR2_X1 U548 ( .A(n433), .B(G110), .ZN(n705) );
  XNOR2_X1 U549 ( .A(n435), .B(n444), .ZN(n438) );
  XOR2_X1 U550 ( .A(G122), .B(n437), .Z(n465) );
  XNOR2_X1 U551 ( .A(n438), .B(n707), .ZN(n607) );
  NOR2_X1 U552 ( .A1(n483), .A2(n607), .ZN(n440) );
  OR2_X1 U553 ( .A1(G237), .A2(G902), .ZN(n500) );
  NAND2_X1 U554 ( .A1(G210), .A2(n500), .ZN(n439) );
  INV_X1 U555 ( .A(n505), .ZN(n512) );
  INV_X1 U556 ( .A(n512), .ZN(n536) );
  NAND2_X1 U557 ( .A1(G227), .A2(n603), .ZN(n441) );
  XNOR2_X1 U558 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U559 ( .A(n446), .B(n445), .ZN(n614) );
  INV_X1 U560 ( .A(KEYINPUT99), .ZN(n471) );
  XNOR2_X1 U561 ( .A(G131), .B(KEYINPUT93), .ZN(n447) );
  XNOR2_X1 U562 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U563 ( .A(G113), .B(n449), .ZN(n453) );
  XNOR2_X1 U564 ( .A(n450), .B(KEYINPUT10), .ZN(n480) );
  XNOR2_X1 U565 ( .A(n451), .B(n480), .ZN(n452) );
  XNOR2_X1 U566 ( .A(n453), .B(n452), .ZN(n460) );
  NAND2_X1 U567 ( .A1(G214), .A2(n454), .ZN(n458) );
  XOR2_X1 U568 ( .A(KEYINPUT92), .B(KEYINPUT11), .Z(n456) );
  XNOR2_X1 U569 ( .A(n456), .B(n455), .ZN(n457) );
  NOR2_X1 U570 ( .A1(n688), .A2(G902), .ZN(n462) );
  XNOR2_X1 U571 ( .A(KEYINPUT95), .B(KEYINPUT13), .ZN(n461) );
  XNOR2_X1 U572 ( .A(n462), .B(n461), .ZN(n464) );
  INV_X1 U573 ( .A(G475), .ZN(n463) );
  XNOR2_X1 U574 ( .A(n464), .B(n463), .ZN(n513) );
  XOR2_X1 U575 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n466) );
  XOR2_X1 U576 ( .A(KEYINPUT80), .B(KEYINPUT8), .Z(n469) );
  NAND2_X1 U577 ( .A1(G234), .A2(n603), .ZN(n468) );
  XNOR2_X1 U578 ( .A(n469), .B(n468), .ZN(n478) );
  NAND2_X1 U579 ( .A1(G217), .A2(n478), .ZN(n470) );
  XOR2_X1 U580 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n473) );
  XNOR2_X1 U581 ( .A(G110), .B(KEYINPUT24), .ZN(n472) );
  XNOR2_X1 U582 ( .A(n473), .B(n472), .ZN(n477) );
  XNOR2_X1 U583 ( .A(G128), .B(G119), .ZN(n475) );
  XOR2_X1 U584 ( .A(n481), .B(n480), .Z(n714) );
  INV_X1 U585 ( .A(n483), .ZN(n599) );
  NAND2_X1 U586 ( .A1(G234), .A2(n599), .ZN(n484) );
  XNOR2_X1 U587 ( .A(KEYINPUT20), .B(n484), .ZN(n492) );
  NAND2_X1 U588 ( .A1(G217), .A2(n492), .ZN(n485) );
  XNOR2_X1 U589 ( .A(KEYINPUT14), .B(n486), .ZN(n489) );
  AND2_X1 U590 ( .A1(G953), .A2(G902), .ZN(n487) );
  NAND2_X1 U591 ( .A1(n489), .A2(n487), .ZN(n552) );
  XNOR2_X1 U592 ( .A(KEYINPUT100), .B(n552), .ZN(n488) );
  NOR2_X1 U593 ( .A1(G900), .A2(n488), .ZN(n491) );
  NAND2_X1 U594 ( .A1(G952), .A2(n489), .ZN(n677) );
  NOR2_X1 U595 ( .A1(n677), .A2(G953), .ZN(n490) );
  XNOR2_X1 U596 ( .A(n490), .B(KEYINPUT84), .ZN(n554) );
  NOR2_X1 U597 ( .A1(n491), .A2(n554), .ZN(n522) );
  NAND2_X1 U598 ( .A1(n492), .A2(G221), .ZN(n493) );
  XNOR2_X1 U599 ( .A(n493), .B(KEYINPUT21), .ZN(n651) );
  NOR2_X1 U600 ( .A1(n522), .A2(n651), .ZN(n494) );
  NAND2_X1 U601 ( .A1(n652), .A2(n494), .ZN(n495) );
  XNOR2_X1 U602 ( .A(KEYINPUT68), .B(n495), .ZN(n507) );
  NOR2_X1 U603 ( .A1(n507), .A2(n583), .ZN(n498) );
  NAND2_X1 U604 ( .A1(n637), .A2(n498), .ZN(n499) );
  NAND2_X1 U605 ( .A1(G214), .A2(n500), .ZN(n662) );
  NAND2_X1 U606 ( .A1(n544), .A2(n662), .ZN(n501) );
  XNOR2_X1 U607 ( .A(KEYINPUT102), .B(n501), .ZN(n502) );
  NOR2_X1 U608 ( .A1(n646), .A2(n502), .ZN(n503) );
  XNOR2_X1 U609 ( .A(n503), .B(KEYINPUT103), .ZN(n504) );
  NOR2_X1 U610 ( .A1(n531), .A2(n513), .ZN(n640) );
  INV_X1 U611 ( .A(n667), .ZN(n527) );
  INV_X1 U612 ( .A(n518), .ZN(n571) );
  NOR2_X1 U613 ( .A1(n507), .A2(n571), .ZN(n508) );
  XNOR2_X1 U614 ( .A(KEYINPUT28), .B(n508), .ZN(n509) );
  NAND2_X1 U615 ( .A1(n509), .A2(n521), .ZN(n516) );
  NOR2_X1 U616 ( .A1(n558), .A2(n516), .ZN(n510) );
  XNOR2_X1 U617 ( .A(n510), .B(KEYINPUT78), .ZN(n635) );
  NAND2_X1 U618 ( .A1(n527), .A2(n635), .ZN(n511) );
  NAND2_X1 U619 ( .A1(n511), .A2(KEYINPUT47), .ZN(n541) );
  INV_X1 U620 ( .A(n513), .ZN(n532) );
  XNOR2_X1 U621 ( .A(KEYINPUT105), .B(KEYINPUT41), .ZN(n514) );
  INV_X1 U622 ( .A(KEYINPUT30), .ZN(n520) );
  NAND2_X1 U623 ( .A1(n518), .A2(n662), .ZN(n519) );
  XNOR2_X1 U624 ( .A(n520), .B(n519), .ZN(n524) );
  NAND2_X1 U625 ( .A1(n521), .A2(n647), .ZN(n586) );
  NOR2_X1 U626 ( .A1(n522), .A2(n586), .ZN(n523) );
  XNOR2_X1 U627 ( .A(n355), .B(KEYINPUT40), .ZN(n733) );
  INV_X1 U628 ( .A(KEYINPUT46), .ZN(n525) );
  XNOR2_X1 U629 ( .A(n526), .B(n525), .ZN(n539) );
  XNOR2_X1 U630 ( .A(KEYINPUT67), .B(KEYINPUT47), .ZN(n528) );
  NAND2_X1 U631 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U632 ( .A(n529), .B(KEYINPUT73), .ZN(n530) );
  NAND2_X1 U633 ( .A1(n530), .A2(n635), .ZN(n537) );
  NOR2_X1 U634 ( .A1(n532), .A2(n531), .ZN(n565) );
  INV_X1 U635 ( .A(n565), .ZN(n533) );
  NOR2_X1 U636 ( .A1(n534), .A2(n533), .ZN(n535) );
  NAND2_X1 U637 ( .A1(n536), .A2(n535), .ZN(n633) );
  NAND2_X1 U638 ( .A1(n537), .A2(n633), .ZN(n538) );
  INV_X1 U639 ( .A(n542), .ZN(n543) );
  AND2_X1 U640 ( .A1(n544), .A2(n543), .ZN(n545) );
  INV_X1 U641 ( .A(n646), .ZN(n574) );
  NAND2_X1 U642 ( .A1(n548), .A2(n640), .ZN(n643) );
  XOR2_X1 U643 ( .A(KEYINPUT98), .B(KEYINPUT33), .Z(n551) );
  INV_X1 U644 ( .A(n589), .ZN(n550) );
  INV_X1 U645 ( .A(n583), .ZN(n549) );
  NOR2_X1 U646 ( .A1(G898), .A2(n552), .ZN(n553) );
  XNOR2_X1 U647 ( .A(KEYINPUT85), .B(n553), .ZN(n556) );
  INV_X1 U648 ( .A(n554), .ZN(n555) );
  NAND2_X1 U649 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U650 ( .A(KEYINPUT86), .B(n557), .ZN(n560) );
  XOR2_X1 U651 ( .A(KEYINPUT82), .B(KEYINPUT0), .Z(n561) );
  XNOR2_X2 U652 ( .A(n562), .B(n561), .ZN(n591) );
  INV_X1 U653 ( .A(n591), .ZN(n563) );
  NOR2_X1 U654 ( .A1(n679), .A2(n563), .ZN(n564) );
  XNOR2_X1 U655 ( .A(n564), .B(KEYINPUT34), .ZN(n566) );
  NAND2_X1 U656 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U657 ( .A(n567), .B(KEYINPUT35), .ZN(n728) );
  INV_X1 U658 ( .A(n652), .ZN(n584) );
  NOR2_X1 U659 ( .A1(n665), .A2(n651), .ZN(n568) );
  NAND2_X1 U660 ( .A1(n591), .A2(n568), .ZN(n570) );
  NAND2_X1 U661 ( .A1(n582), .A2(n571), .ZN(n572) );
  NOR2_X1 U662 ( .A1(n584), .A2(n572), .ZN(n628) );
  NOR2_X1 U663 ( .A1(n728), .A2(n628), .ZN(n580) );
  XNOR2_X1 U664 ( .A(KEYINPUT77), .B(n583), .ZN(n573) );
  NOR2_X1 U665 ( .A1(n584), .A2(n573), .ZN(n577) );
  NAND2_X1 U666 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U667 ( .A1(n580), .A2(n729), .ZN(n581) );
  AND2_X1 U668 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U669 ( .A1(n585), .A2(n584), .ZN(n621) );
  NOR2_X1 U670 ( .A1(n586), .A2(n657), .ZN(n587) );
  NAND2_X1 U671 ( .A1(n591), .A2(n587), .ZN(n588) );
  XNOR2_X1 U672 ( .A(KEYINPUT89), .B(n588), .ZN(n624) );
  NOR2_X1 U673 ( .A1(n590), .A2(n589), .ZN(n659) );
  INV_X1 U674 ( .A(KEYINPUT2), .ZN(n594) );
  XOR2_X1 U675 ( .A(n643), .B(KEYINPUT79), .Z(n595) );
  AND2_X1 U676 ( .A1(n595), .A2(KEYINPUT2), .ZN(n596) );
  AND2_X1 U677 ( .A1(n700), .A2(n596), .ZN(n598) );
  NAND2_X1 U678 ( .A1(n598), .A2(n597), .ZN(n682) );
  AND2_X2 U679 ( .A1(n682), .A2(n483), .ZN(n600) );
  XNOR2_X1 U680 ( .A(n602), .B(n601), .ZN(n604) );
  NOR2_X2 U681 ( .A1(n604), .A2(n699), .ZN(n606) );
  XNOR2_X1 U682 ( .A(KEYINPUT63), .B(KEYINPUT83), .ZN(n605) );
  XNOR2_X1 U683 ( .A(n606), .B(n605), .ZN(G57) );
  XNOR2_X1 U684 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n609) );
  XNOR2_X1 U685 ( .A(n607), .B(KEYINPUT55), .ZN(n608) );
  XNOR2_X1 U686 ( .A(n609), .B(n608), .ZN(n611) );
  XNOR2_X1 U687 ( .A(n613), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U688 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n616) );
  XNOR2_X1 U689 ( .A(n614), .B(KEYINPUT57), .ZN(n615) );
  XNOR2_X1 U690 ( .A(n616), .B(n615), .ZN(n617) );
  INV_X1 U691 ( .A(KEYINPUT121), .ZN(n619) );
  XNOR2_X1 U692 ( .A(n620), .B(n619), .ZN(G54) );
  XNOR2_X1 U693 ( .A(G101), .B(n621), .ZN(G3) );
  XOR2_X1 U694 ( .A(G104), .B(KEYINPUT107), .Z(n623) );
  NAND2_X1 U695 ( .A1(n624), .A2(n637), .ZN(n622) );
  XNOR2_X1 U696 ( .A(n623), .B(n622), .ZN(G6) );
  XOR2_X1 U697 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n626) );
  NAND2_X1 U698 ( .A1(n624), .A2(n640), .ZN(n625) );
  XNOR2_X1 U699 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X1 U700 ( .A(G107), .B(n627), .ZN(G9) );
  XOR2_X1 U701 ( .A(n628), .B(G110), .Z(G12) );
  XOR2_X1 U702 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n630) );
  NAND2_X1 U703 ( .A1(n640), .A2(n635), .ZN(n629) );
  XNOR2_X1 U704 ( .A(n630), .B(n629), .ZN(n632) );
  XOR2_X1 U705 ( .A(G128), .B(KEYINPUT29), .Z(n631) );
  XNOR2_X1 U706 ( .A(n632), .B(n631), .ZN(G30) );
  XNOR2_X1 U707 ( .A(G143), .B(KEYINPUT110), .ZN(n634) );
  XNOR2_X1 U708 ( .A(n634), .B(n633), .ZN(G45) );
  NAND2_X1 U709 ( .A1(n635), .A2(n637), .ZN(n636) );
  XNOR2_X1 U710 ( .A(n636), .B(G146), .ZN(G48) );
  XOR2_X1 U711 ( .A(G113), .B(KEYINPUT111), .Z(n639) );
  NAND2_X1 U712 ( .A1(n637), .A2(n641), .ZN(n638) );
  XNOR2_X1 U713 ( .A(n639), .B(n638), .ZN(G15) );
  NAND2_X1 U714 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U715 ( .A(n642), .B(G116), .ZN(G18) );
  XNOR2_X1 U716 ( .A(G134), .B(n643), .ZN(G36) );
  XNOR2_X1 U717 ( .A(G140), .B(n644), .ZN(n645) );
  XNOR2_X1 U718 ( .A(n645), .B(KEYINPUT113), .ZN(G42) );
  NOR2_X1 U719 ( .A1(n647), .A2(n646), .ZN(n649) );
  XNOR2_X1 U720 ( .A(KEYINPUT50), .B(KEYINPUT115), .ZN(n648) );
  XNOR2_X1 U721 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U722 ( .A(KEYINPUT114), .B(n650), .ZN(n655) );
  NAND2_X1 U723 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U724 ( .A(KEYINPUT49), .B(n653), .Z(n654) );
  NAND2_X1 U725 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U726 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U727 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U728 ( .A(KEYINPUT51), .B(n660), .Z(n661) );
  NOR2_X1 U729 ( .A1(n678), .A2(n661), .ZN(n673) );
  NOR2_X1 U730 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U731 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U732 ( .A(n666), .B(KEYINPUT116), .ZN(n670) );
  NOR2_X1 U733 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U734 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U735 ( .A1(n679), .A2(n671), .ZN(n672) );
  NOR2_X1 U736 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U737 ( .A(n674), .B(KEYINPUT117), .Z(n675) );
  XNOR2_X1 U738 ( .A(KEYINPUT52), .B(n675), .ZN(n676) );
  NOR2_X1 U739 ( .A1(n677), .A2(n676), .ZN(n681) );
  NOR2_X1 U740 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U741 ( .A1(n681), .A2(n680), .ZN(n684) );
  NAND2_X1 U742 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U743 ( .A1(G953), .A2(n685), .ZN(n687) );
  XNOR2_X1 U744 ( .A(KEYINPUT118), .B(KEYINPUT53), .ZN(n686) );
  XNOR2_X1 U745 ( .A(n687), .B(n686), .ZN(G75) );
  XNOR2_X1 U746 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U747 ( .A(n692), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U748 ( .A(n694), .B(n693), .ZN(n695) );
  NOR2_X1 U749 ( .A1(n699), .A2(n695), .ZN(G63) );
  XNOR2_X1 U750 ( .A(n697), .B(n696), .ZN(n698) );
  NOR2_X1 U751 ( .A1(n699), .A2(n698), .ZN(G66) );
  NAND2_X1 U752 ( .A1(n603), .A2(n700), .ZN(n704) );
  NAND2_X1 U753 ( .A1(G953), .A2(G224), .ZN(n701) );
  XNOR2_X1 U754 ( .A(KEYINPUT61), .B(n701), .ZN(n702) );
  NAND2_X1 U755 ( .A1(n702), .A2(G898), .ZN(n703) );
  NAND2_X1 U756 ( .A1(n704), .A2(n703), .ZN(n711) );
  XOR2_X1 U757 ( .A(G101), .B(n705), .Z(n706) );
  XNOR2_X1 U758 ( .A(n707), .B(n706), .ZN(n709) );
  NOR2_X1 U759 ( .A1(G898), .A2(n603), .ZN(n708) );
  NOR2_X1 U760 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U761 ( .A(n711), .B(n710), .ZN(n713) );
  XOR2_X1 U762 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n712) );
  XNOR2_X1 U763 ( .A(n713), .B(n712), .ZN(G69) );
  XOR2_X1 U764 ( .A(n715), .B(n714), .Z(n716) );
  XNOR2_X1 U765 ( .A(KEYINPUT124), .B(n716), .ZN(n722) );
  INV_X1 U766 ( .A(n722), .ZN(n717) );
  XNOR2_X1 U767 ( .A(n717), .B(KEYINPUT125), .ZN(n718) );
  XNOR2_X1 U768 ( .A(n719), .B(n718), .ZN(n720) );
  NAND2_X1 U769 ( .A1(n603), .A2(n720), .ZN(n721) );
  XNOR2_X1 U770 ( .A(KEYINPUT126), .B(n721), .ZN(n727) );
  XNOR2_X1 U771 ( .A(G227), .B(n722), .ZN(n723) );
  NAND2_X1 U772 ( .A1(n723), .A2(G900), .ZN(n724) );
  NAND2_X1 U773 ( .A1(G953), .A2(n724), .ZN(n725) );
  XOR2_X1 U774 ( .A(KEYINPUT127), .B(n725), .Z(n726) );
  NAND2_X1 U775 ( .A1(n727), .A2(n726), .ZN(G72) );
  XOR2_X1 U776 ( .A(n728), .B(G122), .Z(G24) );
  XNOR2_X1 U777 ( .A(n729), .B(G119), .ZN(G21) );
  XOR2_X1 U778 ( .A(KEYINPUT37), .B(KEYINPUT112), .Z(n732) );
  XNOR2_X1 U779 ( .A(n730), .B(G125), .ZN(n731) );
  XNOR2_X1 U780 ( .A(n732), .B(n731), .ZN(G27) );
  XOR2_X1 U781 ( .A(n733), .B(G131), .Z(G33) );
  XOR2_X1 U782 ( .A(G137), .B(n734), .Z(G39) );
endmodule

