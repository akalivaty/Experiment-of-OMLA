

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580;

  XOR2_X1 U322 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n291) );
  XNOR2_X1 U323 ( .A(G1GAT), .B(G57GAT), .ZN(n290) );
  XNOR2_X1 U324 ( .A(n291), .B(n290), .ZN(n309) );
  XOR2_X1 U325 ( .A(G85GAT), .B(G155GAT), .Z(n293) );
  XNOR2_X1 U326 ( .A(G127GAT), .B(G148GAT), .ZN(n292) );
  XNOR2_X1 U327 ( .A(n293), .B(n292), .ZN(n295) );
  XOR2_X1 U328 ( .A(G29GAT), .B(G162GAT), .Z(n294) );
  XNOR2_X1 U329 ( .A(n295), .B(n294), .ZN(n305) );
  XOR2_X1 U330 ( .A(G120GAT), .B(KEYINPUT0), .Z(n297) );
  XNOR2_X1 U331 ( .A(G113GAT), .B(G134GAT), .ZN(n296) );
  XNOR2_X1 U332 ( .A(n297), .B(n296), .ZN(n345) );
  XOR2_X1 U333 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n299) );
  XNOR2_X1 U334 ( .A(G141GAT), .B(KEYINPUT89), .ZN(n298) );
  XNOR2_X1 U335 ( .A(n299), .B(n298), .ZN(n377) );
  XNOR2_X1 U336 ( .A(n345), .B(n377), .ZN(n303) );
  XOR2_X1 U337 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n301) );
  XNOR2_X1 U338 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n300) );
  XNOR2_X1 U339 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U340 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U341 ( .A(n305), .B(n304), .ZN(n307) );
  NAND2_X1 U342 ( .A1(G225GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U343 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U344 ( .A(n309), .B(n308), .Z(n543) );
  XOR2_X1 U345 ( .A(KEYINPUT75), .B(KEYINPUT33), .Z(n311) );
  NAND2_X1 U346 ( .A1(G230GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U347 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U348 ( .A(n312), .B(KEYINPUT31), .Z(n317) );
  XNOR2_X1 U349 ( .A(G71GAT), .B(G57GAT), .ZN(n313) );
  XNOR2_X1 U350 ( .A(n313), .B(KEYINPUT13), .ZN(n428) );
  XOR2_X1 U351 ( .A(KEYINPUT74), .B(G64GAT), .Z(n315) );
  XNOR2_X1 U352 ( .A(G176GAT), .B(G204GAT), .ZN(n314) );
  XNOR2_X1 U353 ( .A(n315), .B(n314), .ZN(n384) );
  XNOR2_X1 U354 ( .A(n428), .B(n384), .ZN(n316) );
  XNOR2_X1 U355 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U356 ( .A(KEYINPUT71), .B(KEYINPUT32), .Z(n319) );
  XNOR2_X1 U357 ( .A(G120GAT), .B(KEYINPUT70), .ZN(n318) );
  XNOR2_X1 U358 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U359 ( .A(n321), .B(n320), .Z(n327) );
  XOR2_X1 U360 ( .A(G78GAT), .B(G148GAT), .Z(n323) );
  XNOR2_X1 U361 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n322) );
  XNOR2_X1 U362 ( .A(n323), .B(n322), .ZN(n366) );
  XOR2_X1 U363 ( .A(G92GAT), .B(KEYINPUT73), .Z(n325) );
  XNOR2_X1 U364 ( .A(G99GAT), .B(G85GAT), .ZN(n324) );
  XNOR2_X1 U365 ( .A(n325), .B(n324), .ZN(n408) );
  XNOR2_X1 U366 ( .A(n366), .B(n408), .ZN(n326) );
  XNOR2_X1 U367 ( .A(n327), .B(n326), .ZN(n569) );
  XOR2_X1 U368 ( .A(G15GAT), .B(G113GAT), .Z(n329) );
  XOR2_X1 U369 ( .A(KEYINPUT68), .B(G1GAT), .Z(n432) );
  XOR2_X1 U370 ( .A(G169GAT), .B(G8GAT), .Z(n381) );
  XNOR2_X1 U371 ( .A(n432), .B(n381), .ZN(n328) );
  XNOR2_X1 U372 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U373 ( .A(n330), .B(G50GAT), .Z(n335) );
  XOR2_X1 U374 ( .A(KEYINPUT29), .B(G197GAT), .Z(n332) );
  XNOR2_X1 U375 ( .A(G22GAT), .B(G141GAT), .ZN(n331) );
  XNOR2_X1 U376 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U377 ( .A(n333), .B(G36GAT), .ZN(n334) );
  XNOR2_X1 U378 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U379 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n337) );
  NAND2_X1 U380 ( .A1(G229GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U381 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U382 ( .A(n339), .B(n338), .Z(n344) );
  XOR2_X1 U383 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n341) );
  XNOR2_X1 U384 ( .A(G43GAT), .B(G29GAT), .ZN(n340) );
  XNOR2_X1 U385 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U386 ( .A(KEYINPUT67), .B(n342), .Z(n419) );
  XNOR2_X1 U387 ( .A(n419), .B(KEYINPUT69), .ZN(n343) );
  XNOR2_X1 U388 ( .A(n344), .B(n343), .ZN(n566) );
  INV_X1 U389 ( .A(n566), .ZN(n472) );
  NOR2_X1 U390 ( .A1(n569), .A2(n472), .ZN(n456) );
  XOR2_X1 U391 ( .A(G15GAT), .B(G127GAT), .Z(n434) );
  XOR2_X1 U392 ( .A(n434), .B(n345), .Z(n347) );
  XNOR2_X1 U393 ( .A(G43GAT), .B(G190GAT), .ZN(n346) );
  XNOR2_X1 U394 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U395 ( .A(KEYINPUT20), .B(KEYINPUT83), .Z(n349) );
  NAND2_X1 U396 ( .A1(G227GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U397 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U398 ( .A(n351), .B(n350), .Z(n356) );
  XOR2_X1 U399 ( .A(G176GAT), .B(KEYINPUT82), .Z(n353) );
  XNOR2_X1 U400 ( .A(G99GAT), .B(G71GAT), .ZN(n352) );
  XNOR2_X1 U401 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U402 ( .A(G169GAT), .B(n354), .ZN(n355) );
  XNOR2_X1 U403 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U404 ( .A(KEYINPUT84), .B(KEYINPUT17), .Z(n358) );
  XNOR2_X1 U405 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n357) );
  XNOR2_X1 U406 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U407 ( .A(KEYINPUT19), .B(n359), .ZN(n380) );
  XOR2_X1 U408 ( .A(n360), .B(n380), .Z(n508) );
  INV_X1 U409 ( .A(n508), .ZN(n549) );
  XOR2_X1 U410 ( .A(KEYINPUT22), .B(KEYINPUT87), .Z(n362) );
  NAND2_X1 U411 ( .A1(G228GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U412 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U413 ( .A(n363), .B(KEYINPUT90), .Z(n368) );
  XOR2_X1 U414 ( .A(G211GAT), .B(KEYINPUT21), .Z(n365) );
  XNOR2_X1 U415 ( .A(G197GAT), .B(G218GAT), .ZN(n364) );
  XNOR2_X1 U416 ( .A(n365), .B(n364), .ZN(n386) );
  XNOR2_X1 U417 ( .A(n386), .B(n366), .ZN(n367) );
  XNOR2_X1 U418 ( .A(n368), .B(n367), .ZN(n375) );
  XOR2_X1 U419 ( .A(G204GAT), .B(KEYINPUT88), .Z(n370) );
  XNOR2_X1 U420 ( .A(KEYINPUT85), .B(KEYINPUT86), .ZN(n369) );
  XNOR2_X1 U421 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U422 ( .A(n371), .B(KEYINPUT23), .Z(n373) );
  XOR2_X1 U423 ( .A(G22GAT), .B(G155GAT), .Z(n433) );
  XNOR2_X1 U424 ( .A(n433), .B(KEYINPUT24), .ZN(n372) );
  XNOR2_X1 U425 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U426 ( .A(n375), .B(n374), .Z(n379) );
  XNOR2_X1 U427 ( .A(G50GAT), .B(KEYINPUT76), .ZN(n376) );
  XNOR2_X1 U428 ( .A(n376), .B(G162GAT), .ZN(n411) );
  XNOR2_X1 U429 ( .A(n411), .B(n377), .ZN(n378) );
  XNOR2_X1 U430 ( .A(n379), .B(n378), .ZN(n545) );
  XOR2_X1 U431 ( .A(n545), .B(KEYINPUT28), .Z(n491) );
  INV_X1 U432 ( .A(n491), .ZN(n469) );
  INV_X1 U433 ( .A(n380), .ZN(n392) );
  XOR2_X1 U434 ( .A(G36GAT), .B(G190GAT), .Z(n407) );
  XNOR2_X1 U435 ( .A(n381), .B(n407), .ZN(n390) );
  XOR2_X1 U436 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n383) );
  NAND2_X1 U437 ( .A1(G226GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U438 ( .A(n383), .B(n382), .ZN(n385) );
  XOR2_X1 U439 ( .A(n385), .B(n384), .Z(n388) );
  XNOR2_X1 U440 ( .A(n386), .B(G92GAT), .ZN(n387) );
  XNOR2_X1 U441 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U442 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U443 ( .A(n392), .B(n391), .Z(n462) );
  INV_X1 U444 ( .A(n462), .ZN(n540) );
  XNOR2_X1 U445 ( .A(KEYINPUT27), .B(n540), .ZN(n401) );
  OR2_X1 U446 ( .A1(n469), .A2(n401), .ZN(n393) );
  NOR2_X1 U447 ( .A1(n543), .A2(n393), .ZN(n509) );
  NAND2_X1 U448 ( .A1(n549), .A2(n509), .ZN(n394) );
  XNOR2_X1 U449 ( .A(n394), .B(KEYINPUT95), .ZN(n406) );
  INV_X1 U450 ( .A(n543), .ZN(n523) );
  NOR2_X1 U451 ( .A1(n549), .A2(n540), .ZN(n395) );
  XNOR2_X1 U452 ( .A(n395), .B(KEYINPUT98), .ZN(n396) );
  NOR2_X1 U453 ( .A1(n545), .A2(n396), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n397), .B(KEYINPUT25), .ZN(n398) );
  XNOR2_X1 U455 ( .A(n398), .B(KEYINPUT99), .ZN(n403) );
  NAND2_X1 U456 ( .A1(n545), .A2(n549), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n399), .B(KEYINPUT96), .ZN(n400) );
  XNOR2_X1 U458 ( .A(KEYINPUT26), .B(n400), .ZN(n564) );
  NOR2_X1 U459 ( .A1(n401), .A2(n564), .ZN(n524) );
  XOR2_X1 U460 ( .A(n524), .B(KEYINPUT97), .Z(n402) );
  NOR2_X1 U461 ( .A1(n403), .A2(n402), .ZN(n404) );
  NOR2_X1 U462 ( .A1(n523), .A2(n404), .ZN(n405) );
  NOR2_X1 U463 ( .A1(n406), .A2(n405), .ZN(n453) );
  XOR2_X1 U464 ( .A(KEYINPUT81), .B(KEYINPUT16), .Z(n442) );
  XOR2_X1 U465 ( .A(KEYINPUT10), .B(n407), .Z(n410) );
  XNOR2_X1 U466 ( .A(G218GAT), .B(n408), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n410), .B(n409), .ZN(n415) );
  XOR2_X1 U468 ( .A(G106GAT), .B(n411), .Z(n413) );
  NAND2_X1 U469 ( .A1(G232GAT), .A2(G233GAT), .ZN(n412) );
  XNOR2_X1 U470 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U471 ( .A(n415), .B(n414), .Z(n421) );
  XOR2_X1 U472 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n417) );
  XNOR2_X1 U473 ( .A(G134GAT), .B(KEYINPUT77), .ZN(n416) );
  XNOR2_X1 U474 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U476 ( .A(n421), .B(n420), .ZN(n518) );
  XOR2_X1 U477 ( .A(KEYINPUT79), .B(G64GAT), .Z(n423) );
  XNOR2_X1 U478 ( .A(G8GAT), .B(G78GAT), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U480 ( .A(KEYINPUT78), .B(KEYINPUT12), .Z(n425) );
  XNOR2_X1 U481 ( .A(KEYINPUT80), .B(KEYINPUT14), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n440) );
  XOR2_X1 U484 ( .A(n428), .B(KEYINPUT15), .Z(n430) );
  NAND2_X1 U485 ( .A1(G231GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n438) );
  XOR2_X1 U488 ( .A(n433), .B(G211GAT), .Z(n436) );
  XNOR2_X1 U489 ( .A(G183GAT), .B(n434), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U491 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n440), .B(n439), .ZN(n499) );
  INV_X1 U493 ( .A(n499), .ZN(n573) );
  NAND2_X1 U494 ( .A1(n518), .A2(n573), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n443) );
  NOR2_X1 U496 ( .A1(n453), .A2(n443), .ZN(n473) );
  NAND2_X1 U497 ( .A1(n456), .A2(n473), .ZN(n450) );
  NOR2_X1 U498 ( .A1(n543), .A2(n450), .ZN(n445) );
  XNOR2_X1 U499 ( .A(KEYINPUT34), .B(KEYINPUT100), .ZN(n444) );
  XNOR2_X1 U500 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U501 ( .A(G1GAT), .B(n446), .Z(G1324GAT) );
  NOR2_X1 U502 ( .A1(n540), .A2(n450), .ZN(n447) );
  XOR2_X1 U503 ( .A(G8GAT), .B(n447), .Z(G1325GAT) );
  NOR2_X1 U504 ( .A1(n549), .A2(n450), .ZN(n449) );
  XNOR2_X1 U505 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n448) );
  XNOR2_X1 U506 ( .A(n449), .B(n448), .ZN(G1326GAT) );
  NOR2_X1 U507 ( .A1(n491), .A2(n450), .ZN(n451) );
  XOR2_X1 U508 ( .A(G22GAT), .B(n451), .Z(G1327GAT) );
  XOR2_X1 U509 ( .A(KEYINPUT103), .B(KEYINPUT39), .Z(n460) );
  XOR2_X1 U510 ( .A(KEYINPUT102), .B(KEYINPUT38), .Z(n458) );
  XOR2_X1 U511 ( .A(KEYINPUT36), .B(KEYINPUT101), .Z(n452) );
  XNOR2_X1 U512 ( .A(n518), .B(n452), .ZN(n577) );
  NOR2_X1 U513 ( .A1(n453), .A2(n577), .ZN(n454) );
  NAND2_X1 U514 ( .A1(n499), .A2(n454), .ZN(n455) );
  XNOR2_X1 U515 ( .A(KEYINPUT37), .B(n455), .ZN(n486) );
  NAND2_X1 U516 ( .A1(n456), .A2(n486), .ZN(n457) );
  XNOR2_X1 U517 ( .A(n458), .B(n457), .ZN(n468) );
  NAND2_X1 U518 ( .A1(n468), .A2(n523), .ZN(n459) );
  XNOR2_X1 U519 ( .A(n460), .B(n459), .ZN(n461) );
  XOR2_X1 U520 ( .A(G29GAT), .B(n461), .Z(G1328GAT) );
  XNOR2_X1 U521 ( .A(G36GAT), .B(KEYINPUT104), .ZN(n464) );
  NAND2_X1 U522 ( .A1(n462), .A2(n468), .ZN(n463) );
  XNOR2_X1 U523 ( .A(n464), .B(n463), .ZN(G1329GAT) );
  XOR2_X1 U524 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n466) );
  NAND2_X1 U525 ( .A1(n468), .A2(n508), .ZN(n465) );
  XNOR2_X1 U526 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U527 ( .A(G43GAT), .B(n467), .ZN(G1330GAT) );
  NAND2_X1 U528 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U529 ( .A(n470), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U530 ( .A(KEYINPUT65), .B(KEYINPUT41), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n569), .B(n471), .ZN(n531) );
  XOR2_X1 U532 ( .A(n531), .B(KEYINPUT107), .Z(n554) );
  AND2_X1 U533 ( .A1(n472), .A2(n554), .ZN(n485) );
  NAND2_X1 U534 ( .A1(n485), .A2(n473), .ZN(n481) );
  NOR2_X1 U535 ( .A1(n481), .A2(n543), .ZN(n477) );
  XOR2_X1 U536 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n475) );
  XNOR2_X1 U537 ( .A(G57GAT), .B(KEYINPUT108), .ZN(n474) );
  XNOR2_X1 U538 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U539 ( .A(n477), .B(n476), .ZN(G1332GAT) );
  NOR2_X1 U540 ( .A1(n540), .A2(n481), .ZN(n478) );
  XOR2_X1 U541 ( .A(G64GAT), .B(n478), .Z(G1333GAT) );
  NOR2_X1 U542 ( .A1(n549), .A2(n481), .ZN(n480) );
  XNOR2_X1 U543 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n479) );
  XNOR2_X1 U544 ( .A(n480), .B(n479), .ZN(G1334GAT) );
  NOR2_X1 U545 ( .A1(n491), .A2(n481), .ZN(n483) );
  XNOR2_X1 U546 ( .A(KEYINPUT43), .B(KEYINPUT110), .ZN(n482) );
  XNOR2_X1 U547 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U548 ( .A(G78GAT), .B(n484), .ZN(G1335GAT) );
  NAND2_X1 U549 ( .A1(n486), .A2(n485), .ZN(n490) );
  NOR2_X1 U550 ( .A1(n543), .A2(n490), .ZN(n487) );
  XOR2_X1 U551 ( .A(G85GAT), .B(n487), .Z(G1336GAT) );
  NOR2_X1 U552 ( .A1(n540), .A2(n490), .ZN(n488) );
  XOR2_X1 U553 ( .A(G92GAT), .B(n488), .Z(G1337GAT) );
  NOR2_X1 U554 ( .A1(n549), .A2(n490), .ZN(n489) );
  XOR2_X1 U555 ( .A(G99GAT), .B(n489), .Z(G1338GAT) );
  NOR2_X1 U556 ( .A1(n491), .A2(n490), .ZN(n492) );
  XOR2_X1 U557 ( .A(KEYINPUT44), .B(n492), .Z(n493) );
  XNOR2_X1 U558 ( .A(G106GAT), .B(n493), .ZN(G1339GAT) );
  NAND2_X1 U559 ( .A1(n566), .A2(n531), .ZN(n494) );
  XNOR2_X1 U560 ( .A(KEYINPUT46), .B(n494), .ZN(n495) );
  NAND2_X1 U561 ( .A1(n495), .A2(n499), .ZN(n496) );
  XNOR2_X1 U562 ( .A(KEYINPUT111), .B(n496), .ZN(n497) );
  NAND2_X1 U563 ( .A1(n497), .A2(n518), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n498), .B(KEYINPUT47), .ZN(n505) );
  NOR2_X1 U565 ( .A1(n499), .A2(n577), .ZN(n500) );
  XOR2_X1 U566 ( .A(KEYINPUT45), .B(n500), .Z(n501) );
  NOR2_X1 U567 ( .A1(n569), .A2(n501), .ZN(n502) );
  XOR2_X1 U568 ( .A(KEYINPUT112), .B(n502), .Z(n503) );
  NOR2_X1 U569 ( .A1(n503), .A2(n566), .ZN(n504) );
  NOR2_X1 U570 ( .A1(n505), .A2(n504), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n506), .B(KEYINPUT64), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n507), .B(KEYINPUT48), .ZN(n541) );
  NAND2_X1 U573 ( .A1(n509), .A2(n508), .ZN(n510) );
  NOR2_X1 U574 ( .A1(n541), .A2(n510), .ZN(n519) );
  NAND2_X1 U575 ( .A1(n519), .A2(n566), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n511), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT49), .B(KEYINPUT113), .Z(n513) );
  NAND2_X1 U578 ( .A1(n519), .A2(n554), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U580 ( .A(G120GAT), .B(n514), .Z(G1341GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n516) );
  NAND2_X1 U582 ( .A1(n519), .A2(n573), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U584 ( .A(G127GAT), .B(n517), .Z(G1342GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n521) );
  INV_X1 U586 ( .A(n518), .ZN(n558) );
  NAND2_X1 U587 ( .A1(n519), .A2(n558), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U589 ( .A(G134GAT), .B(n522), .Z(G1343GAT) );
  NAND2_X1 U590 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U591 ( .A1(n541), .A2(n525), .ZN(n536) );
  NAND2_X1 U592 ( .A1(n536), .A2(n566), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n526), .B(KEYINPUT116), .ZN(n527) );
  XNOR2_X1 U594 ( .A(G141GAT), .B(n527), .ZN(G1344GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n529) );
  XNOR2_X1 U596 ( .A(G148GAT), .B(KEYINPUT117), .ZN(n528) );
  XNOR2_X1 U597 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U598 ( .A(KEYINPUT52), .B(n530), .Z(n533) );
  NAND2_X1 U599 ( .A1(n536), .A2(n531), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n533), .B(n532), .ZN(G1345GAT) );
  XOR2_X1 U601 ( .A(G155GAT), .B(KEYINPUT119), .Z(n535) );
  NAND2_X1 U602 ( .A1(n536), .A2(n573), .ZN(n534) );
  XNOR2_X1 U603 ( .A(n535), .B(n534), .ZN(G1346GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n538) );
  NAND2_X1 U605 ( .A1(n536), .A2(n558), .ZN(n537) );
  XNOR2_X1 U606 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U607 ( .A(G162GAT), .B(n539), .ZN(G1347GAT) );
  NOR2_X1 U608 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U609 ( .A(KEYINPUT54), .B(n542), .ZN(n544) );
  NAND2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n565) );
  NOR2_X1 U611 ( .A1(n545), .A2(n565), .ZN(n547) );
  XNOR2_X1 U612 ( .A(KEYINPUT55), .B(KEYINPUT122), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(n548) );
  NOR2_X1 U614 ( .A1(n549), .A2(n548), .ZN(n559) );
  NAND2_X1 U615 ( .A1(n566), .A2(n559), .ZN(n550) );
  XNOR2_X1 U616 ( .A(G169GAT), .B(n550), .ZN(G1348GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n552) );
  XNOR2_X1 U618 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U620 ( .A(KEYINPUT56), .B(n553), .Z(n556) );
  NAND2_X1 U621 ( .A1(n554), .A2(n559), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1349GAT) );
  NAND2_X1 U623 ( .A1(n573), .A2(n559), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U625 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n561) );
  NAND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1351GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n563) );
  XNOR2_X1 U629 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n568) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n575) );
  NAND2_X1 U632 ( .A1(n575), .A2(n566), .ZN(n567) );
  XOR2_X1 U633 ( .A(n568), .B(n567), .Z(G1352GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n571) );
  NAND2_X1 U635 ( .A1(n575), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G204GAT), .B(n572), .ZN(G1353GAT) );
  NAND2_X1 U638 ( .A1(n573), .A2(n575), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U640 ( .A(n575), .ZN(n576) );
  NOR2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n579) );
  XNOR2_X1 U642 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(n580), .ZN(G1355GAT) );
endmodule

