//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 1 0 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  INV_X1    g0013(.A(new_n201), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n208), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(KEYINPUT65), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n222), .A2(KEYINPUT65), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n210), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n213), .B(new_n219), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n202), .A2(G68), .ZN(new_n243));
  INV_X1    g0043(.A(G68), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G50), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n242), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n253));
  AND2_X1   g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(G222), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G77), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n254), .A2(G1698), .ZN(new_n258));
  INV_X1    g0058(.A(G223), .ZN(new_n259));
  OAI221_X1 g0059(.A(new_n256), .B1(new_n257), .B2(new_n254), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  AND2_X1   g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(new_n217), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n264));
  INV_X1    g0064(.A(G274), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(KEYINPUT66), .B1(new_n261), .B2(new_n217), .ZN(new_n267));
  AND2_X1   g0067(.A1(G1), .A2(G13), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT66), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n266), .A2(new_n267), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT67), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT67), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n266), .A2(new_n267), .A3(new_n274), .A4(new_n271), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  AND3_X1   g0076(.A1(new_n267), .A2(new_n271), .A3(new_n264), .ZN(new_n277));
  XOR2_X1   g0077(.A(KEYINPUT68), .B(G226), .Z(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n263), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G200), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT8), .B(G58), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n208), .A2(G33), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n217), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G13), .ZN(new_n290));
  NOR3_X1   g0090(.A1(new_n290), .A2(new_n208), .A3(G1), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(new_n288), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n202), .B1(new_n207), .B2(G20), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n292), .A2(new_n293), .B1(new_n202), .B2(new_n291), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT9), .ZN(new_n296));
  INV_X1    g0096(.A(G190), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n281), .B(new_n296), .C1(new_n297), .C2(new_n280), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n298), .A2(KEYINPUT10), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(KEYINPUT10), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n295), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n302), .B1(new_n280), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(G179), .B2(new_n280), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n277), .A2(G244), .ZN(new_n306));
  INV_X1    g0106(.A(G238), .ZN(new_n307));
  INV_X1    g0107(.A(G107), .ZN(new_n308));
  OAI22_X1  g0108(.A1(new_n258), .A2(new_n307), .B1(new_n308), .B2(new_n254), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n251), .A2(new_n253), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n310), .A2(new_n232), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n309), .B1(new_n255), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n262), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n276), .B(new_n306), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G200), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n288), .B1(new_n207), .B2(G20), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G77), .ZN(new_n317));
  INV_X1    g0117(.A(new_n291), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n317), .B1(G77), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(G20), .A2(G77), .ZN(new_n320));
  INV_X1    g0120(.A(new_n282), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT15), .B(G87), .ZN(new_n322));
  OAI221_X1 g0122(.A(new_n320), .B1(new_n284), .B2(new_n321), .C1(new_n285), .C2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n319), .B1(new_n288), .B2(new_n323), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n315), .B(new_n324), .C1(new_n297), .C2(new_n314), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n324), .B1(new_n314), .B2(new_n303), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(G179), .B2(new_n314), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n301), .A2(new_n305), .A3(new_n325), .A4(new_n327), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n250), .A2(KEYINPUT70), .A3(G33), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT70), .B1(new_n250), .B2(G33), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n253), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT7), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n250), .A2(G33), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT70), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(new_n252), .B2(KEYINPUT3), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n250), .A2(KEYINPUT70), .A3(G33), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n334), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n333), .B1(new_n338), .B2(G20), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n332), .A2(new_n339), .A3(KEYINPUT71), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT71), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n341), .B(new_n333), .C1(new_n338), .C2(G20), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n340), .A2(G68), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G58), .A2(G68), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n214), .A2(new_n344), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n345), .A2(G20), .B1(G159), .B2(new_n282), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n343), .A2(KEYINPUT16), .A3(new_n346), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT73), .B1(new_n252), .B2(KEYINPUT3), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT73), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n350), .A2(new_n250), .A3(G33), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n349), .A2(new_n351), .A3(new_n253), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n333), .B1(new_n352), .B2(new_n208), .ZN(new_n353));
  AOI211_X1 g0153(.A(KEYINPUT7), .B(G20), .C1(new_n251), .C2(new_n253), .ZN(new_n354));
  NOR3_X1   g0154(.A1(new_n353), .A2(new_n354), .A3(new_n244), .ZN(new_n355));
  INV_X1    g0155(.A(new_n346), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n348), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n347), .A2(new_n357), .A3(new_n288), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n318), .A2(new_n284), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n316), .B2(new_n284), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n273), .A2(new_n275), .B1(new_n277), .B2(G232), .ZN(new_n362));
  INV_X1    g0162(.A(G179), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n259), .A2(new_n255), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(G226), .B2(new_n255), .ZN(new_n365));
  INV_X1    g0165(.A(G87), .ZN(new_n366));
  OAI22_X1  g0166(.A1(new_n331), .A2(new_n365), .B1(new_n252), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n262), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n362), .A2(new_n363), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT74), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT74), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n362), .A2(new_n371), .A3(new_n363), .A4(new_n368), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n362), .A2(new_n368), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n303), .ZN(new_n374));
  AND3_X1   g0174(.A1(new_n370), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n361), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT18), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT18), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n361), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G200), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n373), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n362), .A2(new_n297), .A3(new_n368), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n358), .A2(new_n360), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT17), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n358), .A2(new_n383), .A3(KEYINPUT17), .A4(new_n360), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n377), .A2(new_n379), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n316), .A2(G68), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n318), .A2(KEYINPUT12), .A3(G68), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT12), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n391), .B1(new_n291), .B2(new_n244), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n389), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n282), .A2(G50), .B1(G20), .B2(new_n244), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(new_n257), .B2(new_n285), .ZN(new_n395));
  AND3_X1   g0195(.A1(new_n395), .A2(KEYINPUT11), .A3(new_n288), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT11), .B1(new_n395), .B2(new_n288), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n393), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n251), .A2(new_n253), .A3(G226), .A4(new_n255), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT69), .ZN(new_n401));
  XNOR2_X1  g0201(.A(new_n400), .B(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(G97), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n252), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n404), .B1(new_n311), .B2(G1698), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n313), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT13), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n277), .A2(G238), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n407), .A2(new_n408), .A3(new_n276), .A4(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n276), .A2(new_n409), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT13), .B1(new_n411), .B2(new_n406), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n303), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT14), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n410), .A2(new_n412), .A3(G179), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(new_n413), .B2(new_n414), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n399), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n410), .A2(new_n412), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n399), .B1(new_n419), .B2(G190), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n380), .B2(new_n419), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n328), .A2(new_n388), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  OR2_X1    g0224(.A1(new_n255), .A2(G264), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n338), .B(new_n425), .C1(G257), .C2(G1698), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n310), .A2(G303), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n313), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT82), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n207), .A2(G45), .A3(G274), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT5), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G41), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT76), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n432), .B2(G41), .ZN(new_n435));
  INV_X1    g0235(.A(G41), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n436), .A2(KEYINPUT76), .A3(KEYINPUT5), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n431), .A2(new_n433), .A3(new_n435), .A4(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NOR3_X1   g0239(.A1(new_n261), .A2(KEYINPUT66), .A3(new_n217), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n269), .B1(new_n268), .B2(new_n270), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT77), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n439), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n267), .A2(new_n271), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT77), .B1(new_n445), .B2(new_n438), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(G45), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(G1), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n436), .A2(KEYINPUT5), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n449), .A2(new_n433), .A3(new_n450), .ZN(new_n451));
  AND4_X1   g0251(.A1(G270), .A2(new_n451), .A3(new_n267), .A4(new_n271), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n430), .B1(new_n447), .B2(new_n453), .ZN(new_n454));
  AOI211_X1 g0254(.A(KEYINPUT82), .B(new_n452), .C1(new_n444), .C2(new_n446), .ZN(new_n455));
  OAI211_X1 g0255(.A(G190), .B(new_n429), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n292), .B1(G1), .B2(new_n252), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G116), .ZN(new_n459));
  INV_X1    g0259(.A(G116), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n291), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT83), .ZN(new_n462));
  XNOR2_X1  g0262(.A(new_n461), .B(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(G33), .A2(G283), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT75), .ZN(new_n465));
  XNOR2_X1  g0265(.A(new_n464), .B(new_n465), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n466), .B(new_n208), .C1(G33), .C2(new_n403), .ZN(new_n467));
  INV_X1    g0267(.A(new_n288), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n468), .B1(G20), .B2(new_n460), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n467), .A2(KEYINPUT20), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT20), .B1(new_n467), .B2(new_n469), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n459), .B(new_n463), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n443), .B1(new_n439), .B2(new_n442), .ZN(new_n474));
  NOR3_X1   g0274(.A1(new_n445), .A2(new_n438), .A3(KEYINPUT77), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n453), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT82), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n447), .A2(new_n430), .A3(new_n453), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n428), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n456), .B(new_n473), .C1(new_n479), .C2(new_n380), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT21), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n472), .A2(G169), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n481), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n479), .A2(G179), .A3(new_n472), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n429), .B1(new_n454), .B2(new_n455), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n485), .A2(KEYINPUT21), .A3(G169), .A4(new_n472), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n480), .A2(new_n483), .A3(new_n484), .A4(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT19), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n285), .B2(new_n403), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n366), .A2(new_n403), .A3(new_n308), .ZN(new_n490));
  XNOR2_X1  g0290(.A(new_n490), .B(KEYINPUT80), .ZN(new_n491));
  AOI21_X1  g0291(.A(G20), .B1(new_n404), .B2(KEYINPUT19), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NOR3_X1   g0293(.A1(new_n331), .A2(G20), .A3(new_n244), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n288), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n322), .A2(new_n291), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n458), .A2(G87), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n336), .A2(new_n337), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n499), .A2(G244), .A3(G1698), .A4(new_n253), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G33), .A2(G116), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n307), .A2(G1698), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n499), .A2(new_n253), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n500), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT79), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n500), .A2(new_n503), .A3(KEYINPUT79), .A4(new_n501), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n506), .A2(new_n262), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n431), .ZN(new_n509));
  OAI21_X1  g0309(.A(G250), .B1(new_n448), .B2(G1), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n445), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n508), .A2(G190), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n313), .B1(new_n504), .B2(new_n505), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n511), .B1(new_n514), .B2(new_n507), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n498), .B(new_n513), .C1(new_n380), .C2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n508), .A2(new_n363), .A3(new_n512), .ZN(new_n517));
  XOR2_X1   g0317(.A(new_n322), .B(KEYINPUT81), .Z(new_n518));
  OAI211_X1 g0318(.A(new_n495), .B(new_n496), .C1(new_n457), .C2(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n517), .B(new_n519), .C1(G169), .C2(new_n515), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n499), .A2(G244), .A3(new_n255), .A4(new_n253), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT4), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n251), .A2(new_n253), .A3(G250), .A4(G1698), .ZN(new_n525));
  AND2_X1   g0325(.A1(KEYINPUT4), .A2(G244), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n251), .A2(new_n253), .A3(new_n526), .A4(new_n255), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n466), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n262), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT78), .ZN(new_n531));
  AND4_X1   g0331(.A1(G257), .A2(new_n451), .A3(new_n267), .A4(new_n271), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n531), .B1(new_n447), .B2(new_n533), .ZN(new_n534));
  AOI211_X1 g0334(.A(KEYINPUT78), .B(new_n532), .C1(new_n444), .C2(new_n446), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n530), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G200), .ZN(new_n537));
  NOR3_X1   g0337(.A1(new_n353), .A2(new_n354), .A3(new_n308), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT6), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n539), .A2(new_n403), .A3(G107), .ZN(new_n540));
  XNOR2_X1  g0340(.A(G97), .B(G107), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n540), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  OAI22_X1  g0342(.A1(new_n542), .A2(new_n208), .B1(new_n257), .B2(new_n321), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n288), .B1(new_n538), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n318), .A2(G97), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n545), .B1(new_n458), .B2(G97), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n533), .B1(new_n474), .B2(new_n475), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n313), .B1(new_n524), .B2(new_n528), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n547), .B1(G190), .B2(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n363), .B(new_n530), .C1(new_n534), .C2(new_n535), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n532), .B1(new_n444), .B2(new_n446), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n530), .A2(new_n553), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n554), .A2(new_n303), .B1(new_n544), .B2(new_n546), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n537), .A2(new_n551), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(KEYINPUT23), .B1(new_n208), .B2(G107), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT23), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n558), .A2(new_n308), .A3(G20), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n208), .A2(G33), .A3(G116), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n557), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT84), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT84), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n557), .A2(new_n559), .A3(new_n560), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n338), .A2(KEYINPUT22), .A3(new_n208), .A4(G87), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT22), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n208), .A2(G87), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n567), .B1(new_n310), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n565), .A2(new_n566), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT24), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT24), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n565), .A2(new_n572), .A3(new_n566), .A4(new_n569), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n468), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT25), .B1(new_n291), .B2(new_n308), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n291), .A2(KEYINPUT25), .A3(new_n308), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  OAI22_X1  g0377(.A1(new_n457), .A2(new_n308), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  OR2_X1    g0379(.A1(G250), .A2(G1698), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(G257), .B2(new_n255), .ZN(new_n581));
  INV_X1    g0381(.A(G294), .ZN(new_n582));
  OAI22_X1  g0382(.A1(new_n331), .A2(new_n581), .B1(new_n252), .B2(new_n582), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n451), .A2(new_n267), .A3(new_n271), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n583), .A2(new_n262), .B1(G264), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(G200), .B1(new_n585), .B2(new_n447), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT85), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n447), .ZN(new_n588));
  OAI22_X1  g0388(.A1(new_n586), .A2(new_n587), .B1(new_n588), .B2(G190), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n586), .A2(new_n587), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n579), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n585), .A2(new_n447), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n363), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n588), .A2(new_n303), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n593), .B(new_n594), .C1(new_n574), .C2(new_n578), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n521), .A2(new_n556), .A3(new_n591), .A4(new_n595), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n424), .A2(new_n487), .A3(new_n596), .ZN(G372));
  INV_X1    g0397(.A(new_n305), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n361), .A2(new_n375), .A3(new_n378), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n378), .B1(new_n361), .B2(new_n375), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n418), .A2(new_n327), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n421), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n386), .A2(new_n387), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n601), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT86), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n301), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n299), .A2(KEYINPUT86), .A3(new_n300), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n598), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n520), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n516), .A2(new_n520), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n552), .A2(new_n555), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT26), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n611), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n483), .A2(new_n486), .A3(new_n484), .A4(new_n595), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n617), .A2(new_n521), .A3(new_n556), .A4(new_n591), .ZN(new_n618));
  OAI21_X1  g0418(.A(KEYINPUT26), .B1(new_n612), .B2(new_n613), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n616), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n423), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n610), .A2(new_n621), .ZN(G369));
  NAND3_X1  g0422(.A1(new_n483), .A2(new_n486), .A3(new_n484), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n624));
  OR2_X1    g0424(.A1(new_n624), .A2(KEYINPUT27), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(KEYINPUT27), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(G213), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(G343), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n473), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n623), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n487), .B2(new_n631), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n633), .A2(G330), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n629), .B1(new_n574), .B2(new_n578), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n591), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n595), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n595), .A2(new_n629), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n634), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n636), .A2(new_n623), .A3(new_n595), .A4(new_n630), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n642), .B1(new_n595), .B2(new_n629), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n641), .A2(new_n643), .ZN(G399));
  INV_X1    g0444(.A(new_n211), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n645), .A2(G41), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n491), .A2(new_n460), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n646), .A2(new_n647), .A3(new_n207), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n648), .B1(new_n216), .B2(new_n646), .ZN(new_n649));
  XOR2_X1   g0449(.A(new_n649), .B(KEYINPUT28), .Z(new_n650));
  INV_X1    g0450(.A(KEYINPUT29), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n620), .A2(new_n651), .A3(new_n630), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n651), .B1(new_n620), .B2(new_n630), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(G330), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT30), .ZN(new_n656));
  OAI211_X1 g0456(.A(G179), .B(new_n429), .C1(new_n454), .C2(new_n455), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n550), .A2(new_n515), .A3(new_n585), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n508), .A2(new_n512), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n530), .A2(new_n553), .A3(new_n585), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n662), .A2(new_n479), .A3(KEYINPUT30), .A4(G179), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n592), .A2(G179), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n485), .A2(new_n536), .A3(new_n664), .A4(new_n660), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n659), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n666), .A2(KEYINPUT31), .A3(new_n629), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(KEYINPUT31), .B1(new_n666), .B2(new_n629), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n521), .A2(new_n556), .A3(new_n591), .ZN(new_n671));
  INV_X1    g0471(.A(new_n487), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n671), .A2(new_n672), .A3(new_n595), .A4(new_n630), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n655), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n654), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n650), .B1(new_n677), .B2(G1), .ZN(G364));
  NOR2_X1   g0478(.A1(new_n290), .A2(G20), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n207), .B1(new_n679), .B2(G45), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n646), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n634), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(G330), .B2(new_n633), .ZN(new_n684));
  INV_X1    g0484(.A(new_n682), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n217), .B1(G20), .B2(new_n303), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(G20), .A2(G179), .ZN(new_n688));
  XOR2_X1   g0488(.A(new_n688), .B(KEYINPUT88), .Z(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G190), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G200), .ZN(new_n691));
  XOR2_X1   g0491(.A(new_n691), .B(KEYINPUT89), .Z(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n689), .A2(new_n297), .A3(new_n380), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT90), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  AOI22_X1  g0499(.A1(new_n693), .A2(G58), .B1(G77), .B2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n208), .A2(G190), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(new_n363), .A3(G200), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT93), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G107), .ZN(new_n708));
  NOR4_X1   g0508(.A1(new_n208), .A2(new_n297), .A3(new_n380), .A4(G179), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(G87), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n708), .A2(new_n254), .A3(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n690), .A2(new_n380), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n711), .B1(G50), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(KEYINPUT91), .B1(G179), .B2(G200), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR3_X1   g0515(.A1(KEYINPUT91), .A2(G179), .A3(G200), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n701), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(G159), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g0519(.A(KEYINPUT92), .B(KEYINPUT32), .Z(new_n720));
  XOR2_X1   g0520(.A(new_n719), .B(new_n720), .Z(new_n721));
  NAND3_X1  g0521(.A1(new_n689), .A2(new_n297), .A3(G200), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n715), .A2(new_n716), .ZN(new_n724));
  OAI21_X1  g0524(.A(G20), .B1(new_n724), .B2(new_n297), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n723), .A2(G68), .B1(new_n725), .B2(G97), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n700), .A2(new_n713), .A3(new_n721), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n699), .A2(G311), .ZN(new_n728));
  INV_X1    g0528(.A(G303), .ZN(new_n729));
  INV_X1    g0529(.A(new_n709), .ZN(new_n730));
  INV_X1    g0530(.A(G283), .ZN(new_n731));
  OAI221_X1 g0531(.A(new_n310), .B1(new_n729), .B2(new_n730), .C1(new_n706), .C2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n717), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n732), .B1(G329), .B2(new_n733), .ZN(new_n734));
  AOI22_X1  g0534(.A1(G322), .A2(new_n691), .B1(new_n712), .B2(G326), .ZN(new_n735));
  XNOR2_X1  g0535(.A(KEYINPUT33), .B(G317), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n723), .A2(new_n736), .B1(new_n725), .B2(G294), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n728), .A2(new_n734), .A3(new_n735), .A4(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n687), .B1(new_n727), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G13), .A2(G33), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G20), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n686), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n645), .A2(new_n310), .ZN(new_n744));
  AOI22_X1  g0544(.A1(new_n744), .A2(G355), .B1(new_n460), .B2(new_n645), .ZN(new_n745));
  XOR2_X1   g0545(.A(new_n745), .B(KEYINPUT87), .Z(new_n746));
  NOR2_X1   g0546(.A1(new_n248), .A2(new_n448), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n645), .A2(new_n338), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(G45), .B2(new_n215), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n746), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  AOI211_X1 g0550(.A(new_n685), .B(new_n739), .C1(new_n743), .C2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n742), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n751), .B1(new_n633), .B2(new_n752), .ZN(new_n753));
  AND2_X1   g0553(.A1(new_n684), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(G396));
  NOR2_X1   g0555(.A1(new_n706), .A2(new_n244), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n331), .B(new_n756), .C1(G50), .C2(new_n709), .ZN(new_n757));
  INV_X1    g0557(.A(G58), .ZN(new_n758));
  INV_X1    g0558(.A(new_n725), .ZN(new_n759));
  INV_X1    g0559(.A(G132), .ZN(new_n760));
  OAI221_X1 g0560(.A(new_n757), .B1(new_n758), .B2(new_n759), .C1(new_n760), .C2(new_n717), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT95), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT34), .ZN(new_n763));
  AOI22_X1  g0563(.A1(G137), .A2(new_n712), .B1(new_n723), .B2(G150), .ZN(new_n764));
  INV_X1    g0564(.A(G143), .ZN(new_n765));
  OAI221_X1 g0565(.A(new_n764), .B1(new_n718), .B2(new_n698), .C1(new_n692), .C2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n762), .B1(new_n763), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(new_n763), .B2(new_n766), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n699), .A2(G116), .ZN(new_n769));
  INV_X1    g0569(.A(G311), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n310), .B1(new_n717), .B2(new_n770), .C1(new_n730), .C2(new_n308), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(G87), .B2(new_n707), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n691), .A2(G294), .B1(G97), .B2(new_n725), .ZN(new_n773));
  AOI22_X1  g0573(.A1(G303), .A2(new_n712), .B1(new_n723), .B2(G283), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n769), .A2(new_n772), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT94), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n686), .B1(new_n768), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n686), .A2(new_n740), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n777), .B(new_n682), .C1(G77), .C2(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n325), .B1(new_n324), .B2(new_n630), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n327), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n327), .A2(new_n629), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n780), .B1(new_n740), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n620), .A2(new_n630), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(new_n784), .ZN(new_n787));
  INV_X1    g0587(.A(new_n784), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n620), .A2(new_n788), .A3(new_n630), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n787), .A2(new_n674), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n787), .A2(new_n789), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n682), .B1(new_n791), .B2(new_n675), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n785), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(G384));
  INV_X1    g0594(.A(new_n542), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n795), .A2(KEYINPUT35), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(KEYINPUT35), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n796), .A2(G116), .A3(new_n218), .A4(new_n797), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT36), .Z(new_n799));
  NAND3_X1  g0599(.A1(new_n216), .A2(G77), .A3(new_n344), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n207), .B(G13), .C1(new_n800), .C2(new_n243), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n398), .A2(new_n630), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n418), .A2(new_n421), .A3(new_n804), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n415), .A2(new_n417), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(new_n803), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(new_n789), .B2(new_n783), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n370), .A2(new_n372), .A3(new_n374), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(new_n358), .B2(new_n360), .ZN(new_n811));
  AND3_X1   g0611(.A1(new_n358), .A2(new_n360), .A3(new_n383), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT98), .ZN(new_n814));
  XNOR2_X1  g0614(.A(KEYINPUT97), .B(KEYINPUT37), .ZN(new_n815));
  INV_X1    g0615(.A(new_n627), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n361), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n813), .A2(new_n814), .A3(new_n815), .A4(new_n817), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n376), .A2(new_n817), .A3(new_n384), .A4(new_n815), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(KEYINPUT98), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n347), .A2(new_n288), .ZN(new_n821));
  INV_X1    g0621(.A(new_n348), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(new_n343), .B2(new_n346), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n360), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n816), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(KEYINPUT96), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT96), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n824), .A2(new_n827), .A3(new_n816), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n824), .A2(new_n375), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n826), .A2(new_n384), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n818), .A2(new_n820), .B1(new_n830), .B2(KEYINPUT37), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n826), .A2(new_n828), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n388), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT38), .ZN(new_n835));
  NOR3_X1   g0635(.A1(new_n831), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n818), .A2(new_n820), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n830), .A2(KEYINPUT37), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(KEYINPUT38), .B1(new_n839), .B2(new_n833), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n809), .B1(new_n836), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n627), .B1(new_n599), .B2(new_n600), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(KEYINPUT99), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT99), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n841), .A2(new_n845), .A3(new_n842), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT39), .ZN(new_n847));
  INV_X1    g0647(.A(new_n817), .ZN(new_n848));
  AND3_X1   g0648(.A1(new_n388), .A2(KEYINPUT100), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(KEYINPUT100), .B1(new_n388), .B2(new_n848), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n813), .A2(new_n817), .ZN(new_n852));
  INV_X1    g0652(.A(new_n815), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n818), .A2(new_n820), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT38), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n847), .B1(new_n856), .B2(new_n836), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n806), .A2(new_n399), .A3(new_n630), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n835), .B1(new_n831), .B2(new_n834), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n839), .A2(KEYINPUT38), .A3(new_n833), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n860), .A2(new_n861), .A3(KEYINPUT39), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n857), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n844), .A2(new_n846), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n423), .B1(new_n652), .B2(new_n653), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n610), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n864), .B(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n670), .A2(new_n673), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n784), .B1(new_n805), .B2(new_n807), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT40), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n870), .B(new_n871), .C1(new_n836), .C2(new_n840), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n868), .A2(new_n869), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT100), .ZN(new_n874));
  NOR3_X1   g0674(.A1(new_n604), .A2(new_n599), .A3(new_n600), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n874), .B1(new_n875), .B2(new_n817), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n388), .A2(KEYINPUT100), .A3(new_n848), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n835), .B1(new_n878), .B2(new_n854), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n873), .B1(new_n879), .B2(new_n861), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n872), .B1(new_n880), .B2(new_n871), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(new_n423), .A3(new_n868), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n868), .A2(new_n869), .A3(new_n871), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(new_n861), .B2(new_n860), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n870), .B1(new_n856), .B2(new_n836), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n884), .B1(new_n885), .B2(KEYINPUT40), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n423), .A2(new_n868), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n882), .A2(new_n888), .A3(G330), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n867), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n679), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n890), .B1(G1), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT101), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n867), .A2(new_n889), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n892), .B2(new_n893), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n802), .B1(new_n894), .B2(new_n896), .ZN(G367));
  XOR2_X1   g0697(.A(new_n646), .B(KEYINPUT41), .Z(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n623), .A2(new_n630), .ZN(new_n900));
  XOR2_X1   g0700(.A(new_n640), .B(new_n900), .Z(new_n901));
  XOR2_X1   g0701(.A(new_n901), .B(new_n634), .Z(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n677), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n547), .A2(new_n629), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n556), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n552), .A2(new_n555), .A3(new_n629), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n643), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT104), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT44), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n911), .A2(KEYINPUT103), .ZN(new_n912));
  OR3_X1    g0712(.A1(new_n909), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n910), .B1(new_n909), .B2(new_n912), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n913), .A2(new_n914), .B1(KEYINPUT103), .B2(new_n911), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT105), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n641), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n913), .A2(KEYINPUT103), .A3(new_n911), .A4(new_n914), .ZN(new_n920));
  OR3_X1    g0720(.A1(new_n643), .A2(KEYINPUT45), .A3(new_n908), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT45), .B1(new_n643), .B2(new_n908), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n917), .B2(new_n641), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n916), .A2(new_n919), .A3(new_n920), .A4(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n920), .A2(new_n924), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n918), .B1(new_n926), .B2(new_n915), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n904), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n899), .B1(new_n928), .B2(new_n676), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n680), .ZN(new_n930));
  INV_X1    g0730(.A(new_n908), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n641), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT102), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n908), .A2(new_n642), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n934), .A2(KEYINPUT42), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n537), .A2(new_n551), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n637), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n629), .B1(new_n937), .B2(new_n613), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n934), .B2(KEYINPUT42), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n498), .A2(new_n630), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n612), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n611), .A2(new_n940), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n935), .A2(new_n939), .B1(KEYINPUT43), .B2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n933), .B(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n945), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n930), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n712), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n949), .A2(new_n770), .B1(new_n582), .B2(new_n722), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n709), .A2(G116), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n951), .B(KEYINPUT46), .Z(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(G317), .B2(new_n733), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n707), .A2(G97), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n953), .A2(new_n331), .A3(new_n954), .ZN(new_n955));
  AOI211_X1 g0755(.A(new_n950), .B(new_n955), .C1(G107), .C2(new_n725), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n956), .B1(new_n731), .B2(new_n698), .C1(new_n729), .C2(new_n692), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n691), .A2(G150), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n244), .B2(new_n759), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n959), .A2(KEYINPUT106), .B1(new_n765), .B2(new_n949), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(KEYINPUT106), .B2(new_n959), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT107), .Z(new_n962));
  NAND2_X1  g0762(.A1(new_n707), .A2(G77), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n733), .A2(G137), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n310), .B1(new_n709), .B2(G58), .ZN(new_n965));
  AND3_X1   g0765(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n966), .B1(new_n202), .B2(new_n698), .C1(new_n718), .C2(new_n722), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n957), .B1(new_n962), .B2(new_n967), .ZN(new_n968));
  XOR2_X1   g0768(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n969));
  XNOR2_X1  g0769(.A(new_n968), .B(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n686), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n941), .A2(new_n742), .A3(new_n942), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n748), .A2(new_n238), .ZN(new_n973));
  INV_X1    g0773(.A(new_n743), .ZN(new_n974));
  INV_X1    g0774(.A(new_n322), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n974), .B1(new_n645), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n685), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n971), .A2(new_n972), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n948), .A2(new_n978), .ZN(G387));
  OAI21_X1  g0779(.A(new_n742), .B1(new_n638), .B2(new_n639), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n744), .A2(new_n647), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(G107), .B2(new_n211), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n235), .A2(new_n448), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT109), .Z(new_n984));
  INV_X1    g0784(.A(new_n748), .ZN(new_n985));
  AOI211_X1 g0785(.A(G45), .B(new_n647), .C1(G68), .C2(G77), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n284), .A2(G50), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT50), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n985), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n982), .B1(new_n984), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n682), .B1(new_n990), .B2(new_n974), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n709), .A2(G77), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n954), .A2(new_n338), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(G150), .B2(new_n733), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n699), .A2(G68), .ZN(new_n995));
  INV_X1    g0795(.A(new_n518), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n996), .A2(new_n725), .B1(new_n712), .B2(G159), .ZN(new_n997));
  INV_X1    g0797(.A(new_n284), .ZN(new_n998));
  AOI22_X1  g0798(.A1(G50), .A2(new_n691), .B1(new_n723), .B2(new_n998), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n994), .A2(new_n995), .A3(new_n997), .A4(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n338), .B1(new_n733), .B2(G326), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(G322), .A2(new_n712), .B1(new_n723), .B2(G311), .ZN(new_n1002));
  INV_X1    g0802(.A(G317), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1002), .B1(new_n729), .B2(new_n698), .C1(new_n692), .C2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT48), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n725), .A2(G283), .B1(G294), .B2(new_n709), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT49), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1001), .B1(new_n460), .B2(new_n706), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1000), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n991), .B1(new_n1013), .B2(new_n686), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n903), .A2(new_n681), .B1(new_n980), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n902), .A2(KEYINPUT111), .A3(new_n676), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n646), .B(KEYINPUT110), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n904), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(KEYINPUT111), .B1(new_n902), .B2(new_n676), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1015), .B1(new_n1018), .B2(new_n1019), .ZN(G393));
  INV_X1    g0820(.A(KEYINPUT113), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n927), .A2(new_n925), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1022), .A2(new_n677), .A3(new_n903), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n927), .A2(new_n904), .A3(new_n925), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1023), .A2(new_n1017), .A3(new_n1024), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n743), .B1(new_n403), .B2(new_n211), .C1(new_n985), .C2(new_n242), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G150), .A2(new_n712), .B1(new_n691), .B2(G159), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT112), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT51), .Z(new_n1029));
  AOI21_X1  g0829(.A(new_n331), .B1(G68), .B2(new_n709), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n765), .B2(new_n717), .C1(new_n706), .C2(new_n366), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n759), .A2(new_n257), .B1(new_n722), .B2(new_n202), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(new_n699), .C2(new_n998), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G311), .A2(new_n691), .B1(new_n712), .B2(G317), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT52), .Z(new_n1035));
  OAI22_X1  g0835(.A1(new_n759), .A2(new_n460), .B1(new_n722), .B2(new_n729), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n733), .A2(G322), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n254), .B1(new_n709), .B2(G283), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n708), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1036), .B(new_n1039), .C1(G294), .C2(new_n699), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n1029), .A2(new_n1033), .B1(new_n1035), .B2(new_n1040), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n682), .B(new_n1026), .C1(new_n1041), .C2(new_n687), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n908), .B2(new_n742), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n1022), .B2(new_n681), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1021), .B1(new_n1025), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1025), .A2(new_n1021), .A3(new_n1044), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(G390));
  NAND2_X1  g0848(.A1(new_n805), .A2(new_n807), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n674), .A2(new_n788), .A3(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1050), .A2(KEYINPUT115), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n809), .A2(new_n859), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n857), .B2(new_n862), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n879), .A2(new_n861), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT114), .ZN(new_n1055));
  AND3_X1   g0855(.A1(new_n805), .A2(new_n807), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1055), .B1(new_n805), .B2(new_n807), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n789), .A2(new_n783), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n859), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1054), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1051), .B1(new_n1053), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1051), .ZN(new_n1064));
  AOI21_X1  g0864(.A(KEYINPUT39), .B1(new_n879), .B2(new_n861), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n862), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1064), .B(new_n1061), .C1(new_n1067), .C2(new_n1052), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1063), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n681), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n682), .B1(new_n998), .B2(new_n779), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT118), .Z(new_n1072));
  NAND2_X1  g0872(.A1(new_n710), .A2(new_n310), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1073), .B(new_n756), .C1(G294), .C2(new_n733), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n699), .A2(G97), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n691), .A2(G116), .B1(G77), .B2(new_n725), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(G283), .A2(new_n712), .B1(new_n723), .B2(G107), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(KEYINPUT54), .B(G143), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n699), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n733), .A2(G125), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n706), .B2(new_n202), .ZN(new_n1083));
  INV_X1    g0883(.A(G150), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n730), .A2(KEYINPUT53), .A3(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(KEYINPUT53), .B1(new_n730), .B2(new_n1084), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n254), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n1083), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n723), .A2(G137), .B1(new_n725), .B2(G159), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G128), .A2(new_n712), .B1(new_n691), .B2(G132), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1081), .A2(new_n1088), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  AND2_X1   g0891(.A1(new_n1078), .A2(new_n1091), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1072), .B1(new_n687), .B2(new_n1092), .C1(new_n1067), .C2(new_n741), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1070), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n674), .A2(new_n423), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n865), .A2(new_n610), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1049), .B1(new_n674), .B2(new_n788), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n666), .A2(new_n629), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT31), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n667), .ZN(new_n1101));
  NOR3_X1   g0901(.A1(new_n596), .A2(new_n487), .A3(new_n629), .ZN(new_n1102));
  OAI211_X1 g0902(.A(G330), .B(new_n788), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1103), .A2(new_n808), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1059), .B1(new_n1097), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1103), .B1(new_n1057), .B2(new_n1056), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1059), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1106), .A2(new_n1107), .A3(new_n1050), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1096), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT116), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1109), .B(new_n1110), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1111), .A2(KEYINPUT117), .A3(new_n1068), .A4(new_n1063), .ZN(new_n1112));
  AOI211_X1 g0912(.A(KEYINPUT116), .B(new_n1096), .C1(new_n1105), .C2(new_n1108), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1096), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1110), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1063), .B(new_n1068), .C1(new_n1113), .C2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1112), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1017), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1063), .A2(new_n1068), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1094), .B1(new_n1120), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(G378));
  NOR2_X1   g0926(.A1(new_n302), .A2(new_n627), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n609), .A2(new_n305), .A3(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n607), .A2(new_n305), .A3(new_n608), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n1127), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n1129), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1132), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT121), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  NOR3_X1   g0936(.A1(new_n886), .A2(new_n655), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1134), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1129), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1138), .A2(KEYINPUT121), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n881), .B2(G330), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n864), .B1(new_n1137), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1136), .B1(new_n886), .B2(new_n655), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1067), .A2(new_n859), .B1(KEYINPUT99), .B2(new_n843), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n881), .A2(G330), .A3(new_n1140), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .A4(new_n846), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT122), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1142), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n1145), .A2(new_n1143), .B1(new_n1144), .B2(new_n846), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(KEYINPUT122), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n740), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n331), .A2(new_n436), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n706), .A2(new_n758), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n992), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1154), .B(new_n1157), .C1(G283), .C2(new_n733), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n699), .A2(new_n996), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n723), .A2(G97), .B1(new_n725), .B2(G68), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G107), .A2(new_n691), .B1(new_n712), .B2(G116), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT58), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1154), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n699), .A2(G137), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n723), .A2(G132), .B1(new_n709), .B2(new_n1080), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n691), .A2(G128), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n712), .A2(G125), .B1(G150), .B2(new_n725), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(KEYINPUT59), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n707), .A2(G159), .ZN(new_n1172));
  AOI211_X1 g0972(.A(G33), .B(G41), .C1(new_n733), .C2(G124), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1163), .B(new_n1164), .C1(new_n1170), .C2(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT119), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n686), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT120), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n685), .B(new_n1178), .C1(new_n202), .C2(new_n778), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1151), .A2(new_n681), .B1(new_n1153), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(KEYINPUT117), .B1(new_n1069), .B2(new_n1111), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1115), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT57), .B1(new_n1183), .B2(new_n1151), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1096), .B1(new_n1112), .B2(new_n1119), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1146), .ZN(new_n1186));
  OAI21_X1  g0986(.A(KEYINPUT57), .B1(new_n1186), .B2(new_n1149), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1017), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1180), .B1(new_n1184), .B2(new_n1188), .ZN(G375));
  NOR2_X1   g0989(.A1(new_n1058), .A2(new_n741), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT123), .Z(new_n1191));
  OAI22_X1  g0991(.A1(new_n759), .A2(new_n202), .B1(new_n722), .B2(new_n1079), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n733), .A2(G128), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n331), .B1(G159), .B2(new_n709), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1156), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n1192), .B(new_n1195), .C1(new_n693), .C2(G137), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT125), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n949), .B2(new_n760), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n712), .A2(KEYINPUT125), .A3(G132), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n699), .A2(G150), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n698), .A2(new_n308), .B1(new_n460), .B2(new_n722), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT124), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n996), .A2(new_n725), .B1(new_n691), .B2(G283), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n582), .B2(new_n949), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n254), .B1(new_n709), .B2(G97), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n963), .B(new_n1205), .C1(new_n729), .C2(new_n717), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1196), .A2(new_n1200), .B1(new_n1202), .B2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1208), .A2(new_n687), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n685), .B(new_n1209), .C1(new_n244), .C2(new_n778), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1114), .A2(new_n681), .B1(new_n1191), .B2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1105), .A2(new_n1096), .A3(new_n1108), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1122), .A2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1211), .B1(new_n1213), .B2(new_n898), .ZN(G381));
  NAND4_X1  g1014(.A1(new_n1046), .A2(new_n948), .A3(new_n978), .A4(new_n1047), .ZN(new_n1215));
  OR2_X1    g1015(.A1(G393), .A2(G396), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(new_n1215), .A2(G384), .A3(G381), .A4(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(G375), .A2(G378), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(G407));
  INV_X1    g1019(.A(G213), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1220), .A2(G343), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1218), .A2(new_n1221), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT126), .Z(new_n1223));
  NAND3_X1  g1023(.A1(new_n1223), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1024(.A(new_n1047), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n947), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n680), .B2(new_n929), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n978), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n1225), .A2(new_n1045), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(G393), .B(new_n754), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1229), .A2(new_n1215), .A3(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1230), .B1(new_n1229), .B2(new_n1215), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  OAI211_X1 g1033(.A(G378), .B(new_n1180), .C1(new_n1184), .C2(new_n1188), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1185), .A2(new_n1235), .A3(new_n898), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1179), .A2(new_n1153), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n681), .B1(new_n1186), .B2(new_n1149), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1125), .B1(new_n1236), .B2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1221), .B1(new_n1234), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1213), .A2(KEYINPUT60), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1242), .B(new_n1017), .C1(KEYINPUT60), .C2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1211), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n793), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1244), .A2(G384), .A3(new_n1211), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT62), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  AND2_X1   g1050(.A1(new_n1241), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1234), .A2(new_n1240), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT127), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1221), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1248), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1234), .A2(KEYINPUT127), .A3(new_n1240), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .A4(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1251), .B1(new_n1258), .B2(new_n1249), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT61), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1221), .A2(G2897), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1248), .B(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1260), .B1(new_n1263), .B2(new_n1241), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1233), .B1(new_n1259), .B2(new_n1264), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1241), .A2(KEYINPUT63), .A3(new_n1256), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n1266), .A2(new_n1233), .A3(KEYINPUT61), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT63), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1254), .A2(new_n1255), .A3(new_n1257), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1268), .B1(new_n1269), .B2(new_n1262), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1258), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1267), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1265), .A2(new_n1272), .ZN(G405));
  INV_X1    g1073(.A(new_n1218), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(G375), .A2(G378), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1256), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1274), .A2(new_n1248), .A3(new_n1275), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1233), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1279), .B(new_n1280), .ZN(G402));
endmodule


