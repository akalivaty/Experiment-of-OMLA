//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n528, new_n529, new_n530, new_n531, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n540, new_n542, new_n543, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n601, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1186, new_n1187, new_n1188;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  XNOR2_X1  g016(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n452), .B(new_n453), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT68), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n462), .B1(new_n454), .B2(G2106), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n468), .B1(new_n469), .B2(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n466), .B1(new_n470), .B2(new_n464), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  OAI211_X1 g048(.A(G137), .B(new_n464), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n469), .A2(KEYINPUT69), .A3(G137), .A4(new_n464), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n471), .A2(new_n478), .ZN(G160));
  OR2_X1    g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  AOI21_X1  g056(.A(G2105), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n464), .B1(new_n480), .B2(new_n481), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  MUX2_X1   g060(.A(G100), .B(G112), .S(G2105), .Z(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2104), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND2_X1  g064(.A1(G114), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G102), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  AOI22_X1  g067(.A1(new_n484), .A2(G126), .B1(G2104), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n482), .B2(G138), .ZN(new_n495));
  OAI211_X1 g070(.A(G138), .B(new_n464), .C1(new_n472), .C2(new_n473), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n493), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(KEYINPUT70), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(KEYINPUT6), .A3(G651), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n500), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G50), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n503), .A2(new_n505), .ZN(new_n508));
  OR2_X1    g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  OAI221_X1 g089(.A(new_n507), .B1(new_n512), .B2(new_n513), .C1(new_n514), .C2(new_n502), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  AOI22_X1  g091(.A1(new_n503), .A2(new_n505), .B1(new_n509), .B2(new_n510), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G89), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n506), .A2(G51), .ZN(new_n519));
  AND2_X1   g094(.A1(G63), .A2(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT7), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT7), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n523), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n511), .A2(new_n520), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n518), .A2(new_n519), .A3(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(G168));
  AOI22_X1  g102(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n502), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT71), .ZN(new_n530));
  AOI22_X1  g105(.A1(G90), .A2(new_n517), .B1(new_n506), .B2(G52), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(G171));
  AOI22_X1  g107(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(new_n502), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n517), .A2(G81), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n506), .A2(G43), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G860), .ZN(G153));
  AND3_X1   g114(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G36), .ZN(G176));
  NAND2_X1  g116(.A1(G1), .A2(G3), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT8), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n540), .A2(new_n543), .ZN(G188));
  NAND2_X1  g119(.A1(new_n506), .A2(G53), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(KEYINPUT9), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT72), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT9), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n506), .A2(new_n548), .A3(G53), .ZN(new_n549));
  AND3_X1   g124(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n547), .B1(new_n546), .B2(new_n549), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT73), .ZN(new_n553));
  INV_X1    g128(.A(G91), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n512), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n517), .A2(KEYINPUT73), .A3(G91), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n511), .A2(G65), .ZN(new_n557));
  INV_X1    g132(.A(G78), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n558), .B2(new_n500), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n555), .A2(new_n556), .B1(new_n559), .B2(G651), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n552), .A2(new_n560), .ZN(G299));
  INV_X1    g136(.A(G171), .ZN(G301));
  XOR2_X1   g137(.A(new_n526), .B(KEYINPUT74), .Z(G286));
  NAND2_X1  g138(.A1(new_n517), .A2(G87), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n506), .A2(G49), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(G288));
  NAND2_X1  g142(.A1(new_n511), .A2(G61), .ZN(new_n568));
  NAND2_X1  g143(.A1(G73), .A2(G543), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G651), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n570), .A2(KEYINPUT75), .A3(G651), .ZN(new_n574));
  AOI22_X1  g149(.A1(G86), .A2(new_n517), .B1(new_n506), .B2(G48), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G305));
  AOI22_X1  g151(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(new_n502), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n517), .A2(G85), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n506), .A2(G47), .ZN(new_n580));
  AND3_X1   g155(.A1(new_n579), .A2(new_n580), .A3(KEYINPUT76), .ZN(new_n581));
  AOI21_X1  g156(.A(KEYINPUT76), .B1(new_n579), .B2(new_n580), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n578), .B1(new_n581), .B2(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G171), .A2(G868), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n517), .A2(G92), .ZN(new_n585));
  XOR2_X1   g160(.A(new_n585), .B(KEYINPUT10), .Z(new_n586));
  AOI22_X1  g161(.A1(new_n511), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT77), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n502), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n589), .B1(new_n588), .B2(new_n587), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n506), .A2(G54), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n586), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n584), .B1(G868), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G284));
  XNOR2_X1  g169(.A(new_n593), .B(KEYINPUT78), .ZN(G321));
  NAND2_X1  g170(.A1(G286), .A2(G868), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n552), .A2(new_n560), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(G297));
  XOR2_X1   g173(.A(G297), .B(KEYINPUT79), .Z(G280));
  AND3_X1   g174(.A1(new_n586), .A2(new_n590), .A3(new_n591), .ZN(new_n600));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(G860), .ZN(G148));
  NAND2_X1  g177(.A1(new_n600), .A2(new_n601), .ZN(new_n603));
  MUX2_X1   g178(.A(new_n537), .B(new_n603), .S(G868), .Z(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g180(.A1(new_n482), .A2(G2104), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT12), .Z(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT80), .ZN(new_n609));
  INV_X1    g184(.A(G2100), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n608), .A2(KEYINPUT13), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(KEYINPUT13), .B2(new_n608), .ZN(new_n612));
  OR3_X1    g187(.A1(new_n612), .A2(new_n609), .A3(new_n610), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n609), .B2(new_n610), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n484), .A2(G123), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT81), .Z(new_n616));
  NAND2_X1  g191(.A1(new_n482), .A2(G135), .ZN(new_n617));
  OAI21_X1  g192(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n618));
  AND2_X1   g193(.A1(new_n618), .A2(KEYINPUT82), .ZN(new_n619));
  OAI22_X1  g194(.A1(new_n618), .A2(KEYINPUT82), .B1(G111), .B2(new_n464), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n616), .B(new_n617), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT83), .B(G2096), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n613), .A2(new_n614), .A3(new_n623), .ZN(G156));
  INV_X1    g199(.A(KEYINPUT14), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT15), .B(G2435), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2438), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2427), .ZN(new_n628));
  INV_X1    g203(.A(G2430), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n625), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(new_n629), .B2(new_n628), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(KEYINPUT84), .B(KEYINPUT16), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G1341), .B(G1348), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n631), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n631), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(G14), .A3(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(G401));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  NOR3_X1   g222(.A1(new_n644), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT18), .ZN(new_n649));
  INV_X1    g224(.A(new_n645), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n650), .A2(KEYINPUT17), .A3(new_n643), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n643), .B1(new_n650), .B2(KEYINPUT17), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n651), .B1(new_n652), .B2(new_n647), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n644), .A2(new_n647), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n650), .B1(new_n654), .B2(KEYINPUT17), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n649), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2096), .ZN(new_n657));
  XOR2_X1   g232(.A(KEYINPUT85), .B(G2100), .Z(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(G1971), .B(G1976), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  XOR2_X1   g238(.A(G1956), .B(G2474), .Z(new_n664));
  XOR2_X1   g239(.A(G1961), .B(G1966), .Z(new_n665));
  AND2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT20), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n664), .A2(new_n665), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n663), .A2(new_n666), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(new_n663), .B2(new_n669), .ZN(new_n671));
  AND2_X1   g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT86), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(G229));
  MUX2_X1   g255(.A(G6), .B(G305), .S(G16), .Z(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT32), .B(G1981), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(G16), .A2(G22), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(G166), .B2(G16), .ZN(new_n685));
  INV_X1    g260(.A(G1971), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G23), .ZN(new_n689));
  INV_X1    g264(.A(G288), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n689), .B1(new_n690), .B2(new_n688), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT33), .B(G1976), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n687), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n683), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(KEYINPUT34), .ZN(new_n697));
  MUX2_X1   g272(.A(G95), .B(G107), .S(G2105), .Z(new_n698));
  AOI22_X1  g273(.A1(G119), .A2(new_n484), .B1(new_n698), .B2(G2104), .ZN(new_n699));
  INV_X1    g274(.A(G131), .ZN(new_n700));
  INV_X1    g275(.A(new_n482), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  MUX2_X1   g277(.A(G25), .B(new_n702), .S(G29), .Z(new_n703));
  XOR2_X1   g278(.A(KEYINPUT35), .B(G1991), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G290), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G16), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G16), .B2(G24), .ZN(new_n708));
  INV_X1    g283(.A(G1986), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n705), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n709), .B2(new_n708), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n696), .B2(KEYINPUT34), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n712), .A2(KEYINPUT87), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(KEYINPUT87), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n697), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n715), .A2(KEYINPUT36), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(KEYINPUT36), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n688), .A2(G21), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G168), .B2(new_n688), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n720), .A2(G1966), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT94), .ZN(new_n722));
  NOR2_X1   g297(.A1(G29), .A2(G33), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT89), .Z(new_n724));
  AND3_X1   g299(.A1(new_n465), .A2(KEYINPUT25), .A3(G103), .ZN(new_n725));
  AOI21_X1  g300(.A(KEYINPUT25), .B1(new_n465), .B2(G103), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n469), .A2(G127), .ZN(new_n728));
  NAND2_X1  g303(.A1(G115), .A2(G2104), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n464), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI211_X1 g305(.A(new_n727), .B(new_n730), .C1(G139), .C2(new_n482), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n724), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT90), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(G2072), .Z(new_n736));
  INV_X1    g311(.A(G1348), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n600), .A2(G16), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G4), .B2(G16), .ZN(new_n739));
  AOI211_X1 g314(.A(new_n722), .B(new_n736), .C1(new_n737), .C2(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(G16), .A2(G19), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n538), .B2(G16), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1341), .ZN(new_n743));
  NOR2_X1   g318(.A1(G171), .A2(new_n688), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G5), .B2(new_n688), .ZN(new_n745));
  INV_X1    g320(.A(G1961), .ZN(new_n746));
  NOR2_X1   g321(.A1(G29), .A2(G35), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G162), .B2(G29), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G2090), .ZN(new_n751));
  OAI22_X1  g326(.A1(new_n745), .A2(new_n746), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AOI211_X1 g327(.A(new_n743), .B(new_n752), .C1(new_n751), .C2(new_n750), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n745), .A2(new_n746), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n733), .A2(G26), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT28), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n482), .A2(G140), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n484), .A2(G128), .ZN(new_n758));
  MUX2_X1   g333(.A(G104), .B(G116), .S(G2105), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G2104), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n756), .B1(new_n762), .B2(new_n733), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT88), .B(G2067), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n621), .A2(new_n733), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n763), .A2(new_n764), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT30), .B(G28), .Z(new_n768));
  NOR2_X1   g343(.A1(new_n768), .A2(G29), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT31), .B(G11), .Z(new_n770));
  NOR4_X1   g345(.A1(new_n766), .A2(new_n767), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n754), .A2(new_n765), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(G27), .A2(G29), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G164), .B2(G29), .ZN(new_n774));
  INV_X1    g349(.A(G2078), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G2084), .ZN(new_n777));
  NAND2_X1  g352(.A1(G160), .A2(G29), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT24), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n733), .B1(new_n779), .B2(G34), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n780), .A2(KEYINPUT91), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n779), .A2(G34), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n780), .B2(KEYINPUT91), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n778), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n733), .A2(G32), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT92), .B(KEYINPUT26), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT93), .ZN(new_n787));
  NAND3_X1  g362(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n787), .B(new_n788), .Z(new_n789));
  AOI22_X1  g364(.A1(new_n482), .A2(G141), .B1(G105), .B2(new_n465), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n484), .A2(G129), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n785), .B1(new_n794), .B2(new_n733), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT27), .B(G1996), .Z(new_n796));
  OAI221_X1 g371(.A(new_n776), .B1(new_n777), .B2(new_n784), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n784), .A2(new_n777), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n720), .A2(G1966), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n739), .A2(new_n737), .ZN(new_n802));
  NOR4_X1   g377(.A1(new_n772), .A2(new_n797), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n688), .A2(G20), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT96), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT23), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G299), .B2(G16), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1956), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n740), .A2(new_n753), .A3(new_n803), .A4(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n718), .A2(new_n809), .ZN(G311));
  OR2_X1    g385(.A1(new_n718), .A2(new_n809), .ZN(G150));
  XOR2_X1   g386(.A(KEYINPUT98), .B(G55), .Z(new_n812));
  AOI22_X1  g387(.A1(G93), .A2(new_n517), .B1(new_n506), .B2(new_n812), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n502), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(G860), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT37), .Z(new_n817));
  XOR2_X1   g392(.A(new_n537), .B(new_n815), .Z(new_n818));
  NOR2_X1   g393(.A1(new_n592), .A2(new_n601), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n818), .B(new_n819), .Z(new_n820));
  XOR2_X1   g395(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n823), .A2(KEYINPUT39), .ZN(new_n824));
  INV_X1    g399(.A(G860), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n823), .B2(KEYINPUT39), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n817), .B1(new_n824), .B2(new_n826), .ZN(G145));
  XNOR2_X1  g402(.A(G160), .B(G162), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(new_n621), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT99), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n495), .B2(new_n497), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n469), .A2(new_n494), .A3(G138), .A4(new_n464), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n832), .A2(new_n833), .A3(KEYINPUT99), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n831), .A2(new_n493), .A3(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(new_n762), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n836), .A2(new_n793), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n793), .ZN(new_n838));
  AOI22_X1  g413(.A1(new_n837), .A2(new_n838), .B1(KEYINPUT100), .B2(new_n732), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n732), .A2(KEYINPUT100), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n607), .B(new_n702), .Z(new_n842));
  NAND2_X1  g417(.A1(new_n484), .A2(G130), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT101), .ZN(new_n844));
  MUX2_X1   g419(.A(G106), .B(G118), .S(G2105), .Z(new_n845));
  AOI22_X1  g420(.A1(G142), .A2(new_n482), .B1(new_n845), .B2(G2104), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n842), .B(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(KEYINPUT102), .B1(new_n841), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n841), .A2(new_n848), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR3_X1   g426(.A1(new_n841), .A2(KEYINPUT102), .A3(new_n848), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n829), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT103), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n848), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n841), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n829), .B1(new_n841), .B2(new_n856), .ZN(new_n858));
  AOI21_X1  g433(.A(G37), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n853), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g436(.A1(new_n815), .A2(G868), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n597), .A2(new_n592), .ZN(new_n863));
  NAND2_X1  g438(.A1(G299), .A2(new_n600), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(KEYINPUT104), .ZN(new_n866));
  NOR2_X1   g441(.A1(G299), .A2(new_n600), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n592), .B1(new_n552), .B2(new_n560), .ZN(new_n868));
  OR3_X1    g443(.A1(new_n867), .A2(new_n868), .A3(KEYINPUT104), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n818), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n603), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT105), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n865), .A2(KEYINPUT41), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT106), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n597), .A2(new_n876), .A3(new_n592), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT41), .ZN(new_n878));
  OAI21_X1  g453(.A(KEYINPUT106), .B1(G299), .B2(new_n600), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .A4(new_n864), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n881), .A2(new_n872), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT105), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n870), .A2(new_n883), .A3(new_n872), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n874), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(KEYINPUT42), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT42), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n874), .A2(new_n887), .A3(new_n882), .A4(new_n884), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(G290), .B(G288), .ZN(new_n890));
  XNOR2_X1  g465(.A(G305), .B(G303), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT107), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n892), .B(new_n893), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n890), .A2(new_n891), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n889), .B(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n862), .B1(new_n897), .B2(G868), .ZN(G295));
  AOI21_X1  g473(.A(new_n862), .B1(new_n897), .B2(G868), .ZN(G331));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n878), .B1(new_n867), .B2(new_n868), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT108), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n877), .A2(KEYINPUT41), .A3(new_n879), .A4(new_n864), .ZN(new_n904));
  OAI211_X1 g479(.A(KEYINPUT108), .B(new_n878), .C1(new_n867), .C2(new_n868), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(G171), .A2(G286), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n907), .B1(new_n526), .B2(G171), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(new_n818), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n906), .A2(KEYINPUT109), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT109), .B1(new_n906), .B2(new_n909), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n866), .A2(new_n869), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n912), .A2(new_n909), .ZN(new_n913));
  NOR3_X1   g488(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n914), .A2(new_n896), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n909), .A2(new_n875), .A3(new_n880), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n908), .B(new_n871), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n865), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n916), .A2(new_n896), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(G37), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT43), .B1(new_n915), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n916), .A2(new_n918), .ZN(new_n925));
  INV_X1    g500(.A(new_n896), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n921), .A2(new_n924), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n900), .B1(new_n923), .B2(new_n928), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n921), .B(new_n924), .C1(new_n914), .C2(new_n896), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT110), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n911), .A2(new_n913), .ZN(new_n933));
  INV_X1    g508(.A(new_n910), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n926), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n936), .A2(KEYINPUT110), .A3(new_n924), .A4(new_n921), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n921), .A2(new_n927), .ZN(new_n938));
  AOI22_X1  g513(.A1(new_n932), .A2(new_n937), .B1(KEYINPUT43), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n929), .B1(new_n939), .B2(new_n900), .ZN(G397));
  NAND3_X1  g515(.A1(new_n469), .A2(G126), .A3(G2105), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n492), .A2(G2104), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n832), .A2(new_n833), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n943), .B1(new_n944), .B2(new_n830), .ZN(new_n945));
  AOI21_X1  g520(.A(G1384), .B1(new_n945), .B2(new_n834), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n465), .A2(G101), .ZN(new_n947));
  OAI21_X1  g522(.A(G125), .B1(new_n472), .B2(new_n473), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n467), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n947), .B1(new_n949), .B2(G2105), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n950), .A2(G40), .A3(new_n476), .A4(new_n477), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n946), .A2(KEYINPUT45), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n761), .B(G2067), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  XOR2_X1   g529(.A(new_n954), .B(KEYINPUT112), .Z(new_n955));
  INV_X1    g530(.A(G1996), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n794), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n955), .B1(new_n952), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n952), .A2(new_n956), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n959), .B(KEYINPUT111), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n794), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n706), .A2(new_n709), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n706), .A2(new_n709), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n952), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n704), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n702), .B(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n952), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n963), .A2(new_n967), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(G303), .A2(G8), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT55), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n972), .B(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n975));
  INV_X1    g550(.A(G1384), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n835), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n498), .A2(new_n976), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n951), .B1(new_n978), .B2(KEYINPUT50), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n977), .A2(new_n979), .A3(new_n751), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n835), .A2(KEYINPUT45), .A3(new_n976), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n951), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(G1971), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  OAI211_X1 g559(.A(G8), .B(new_n974), .C1(new_n980), .C2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT113), .ZN(new_n986));
  AOI211_X1 g561(.A(new_n982), .B(G1384), .C1(new_n945), .C2(new_n834), .ZN(new_n987));
  INV_X1    g562(.A(G40), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n471), .A2(new_n478), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(G1384), .B1(new_n944), .B2(new_n493), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n989), .B1(KEYINPUT45), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n686), .B1(new_n987), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n977), .A2(new_n979), .A3(new_n751), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT113), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n994), .A2(new_n995), .A3(G8), .A4(new_n974), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n986), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n835), .A2(new_n989), .A3(new_n976), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n690), .A2(G1976), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n998), .A2(G8), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n1001));
  INV_X1    g576(.A(G1976), .ZN(new_n1002));
  NAND2_X1  g577(.A1(G288), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n1000), .A2(KEYINPUT114), .A3(new_n1001), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n506), .A2(G48), .ZN(new_n1005));
  XNOR2_X1  g580(.A(KEYINPUT115), .B(G86), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n571), .B(new_n1005), .C1(new_n512), .C2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(G1981), .ZN(new_n1008));
  INV_X1    g583(.A(G1981), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n573), .A2(new_n1009), .A3(new_n574), .A4(new_n575), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT116), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1012), .A2(KEYINPUT49), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G8), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1015), .B1(new_n946), .B2(new_n989), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1008), .B(new_n1010), .C1(new_n1012), .C2(KEYINPUT49), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1004), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n998), .A2(G8), .A3(new_n999), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT52), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT52), .B1(G288), .B2(new_n1002), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1021), .A2(KEYINPUT114), .B1(new_n1000), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1019), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n974), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n835), .A2(KEYINPUT50), .A3(new_n976), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n990), .A2(KEYINPUT50), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n951), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n984), .B1(new_n751), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1025), .B1(new_n1030), .B2(new_n1015), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n990), .A2(KEYINPUT45), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n989), .B(new_n1032), .C1(new_n946), .C2(KEYINPUT45), .ZN(new_n1033));
  INV_X1    g608(.A(G1966), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n977), .A2(new_n979), .A3(new_n777), .ZN(new_n1036));
  AOI211_X1 g611(.A(new_n1015), .B(G286), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n997), .A2(new_n1024), .A3(new_n1031), .A4(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT63), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n994), .A2(G8), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1039), .B1(new_n1041), .B2(new_n1025), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n997), .A2(new_n1024), .A3(new_n1037), .A4(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1018), .A2(new_n1002), .A3(new_n690), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n1010), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1016), .B(KEYINPUT117), .ZN(new_n1047));
  INV_X1    g622(.A(new_n997), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1046), .A2(new_n1047), .B1(new_n1048), .B2(new_n1024), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1044), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n977), .A2(new_n979), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n737), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n998), .A2(G2067), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n592), .A2(KEYINPUT60), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n981), .A2(new_n983), .A3(new_n956), .ZN(new_n1056));
  XOR2_X1   g631(.A(KEYINPUT58), .B(G1341), .Z(new_n1057));
  NAND2_X1  g632(.A1(new_n998), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n538), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT59), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT59), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(new_n1062), .A3(new_n538), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1055), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT61), .ZN(new_n1065));
  XNOR2_X1  g640(.A(KEYINPUT56), .B(G2072), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n981), .A2(new_n983), .A3(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(KEYINPUT57), .B(new_n560), .C1(new_n550), .C2(new_n551), .ZN(new_n1068));
  XOR2_X1   g643(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n1069));
  NAND2_X1  g644(.A1(new_n555), .A2(new_n556), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n559), .A2(G651), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n546), .A2(new_n549), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1069), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1068), .A2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1067), .B(new_n1075), .C1(new_n1029), .C2(G1956), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G1956), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1027), .B1(new_n946), .B2(KEYINPUT50), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1078), .B1(new_n1079), .B2(new_n951), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1075), .B1(new_n1080), .B2(new_n1067), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1065), .B1(new_n1077), .B2(new_n1081), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1052), .A2(new_n592), .A3(new_n1053), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n592), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT60), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n989), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n987), .A2(new_n991), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1087), .A2(new_n1078), .B1(new_n1088), .B2(new_n1066), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1068), .A2(new_n1074), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1090), .B1(new_n1068), .B2(new_n1074), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g668(.A(KEYINPUT61), .B(new_n1076), .C1(new_n1089), .C2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1064), .A2(new_n1082), .A3(new_n1085), .A4(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1089), .A2(new_n1093), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1096), .B1(new_n1084), .B2(new_n1076), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1095), .A2(KEYINPUT120), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT120), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n981), .A2(new_n983), .A3(new_n775), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1102), .A2(KEYINPUT124), .A3(new_n1103), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1106), .A2(new_n1107), .B1(new_n746), .B2(new_n1051), .ZN(new_n1108));
  INV_X1    g683(.A(new_n946), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n951), .B1(new_n1109), .B2(new_n982), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1110), .A2(KEYINPUT123), .A3(new_n775), .A4(new_n1032), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT123), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(new_n1033), .B2(G2078), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1111), .A2(KEYINPUT53), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(G301), .B1(new_n1108), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1051), .A2(new_n746), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1110), .A2(KEYINPUT53), .A3(new_n775), .A4(new_n981), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1102), .A2(KEYINPUT124), .A3(new_n1103), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT124), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1116), .B(new_n1117), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1120), .A2(G171), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1101), .B1(new_n1115), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1108), .A2(G301), .A3(new_n1114), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1120), .A2(G171), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1123), .A2(KEYINPUT54), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1127), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n526), .A2(G8), .ZN(new_n1130));
  XOR2_X1   g705(.A(new_n1130), .B(KEYINPUT122), .Z(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1035), .A2(new_n1127), .A3(new_n1036), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1129), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n1035), .A2(new_n1127), .A3(new_n1036), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1135), .A2(new_n1128), .A3(new_n1015), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1134), .B(KEYINPUT51), .C1(new_n1136), .C2(new_n1132), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n997), .A2(new_n1024), .A3(new_n1031), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1132), .A2(KEYINPUT51), .ZN(new_n1139));
  AND2_X1   g714(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1139), .B1(new_n1140), .B2(new_n1015), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1137), .A2(new_n1138), .A3(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1126), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1050), .B1(new_n1100), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1137), .A2(KEYINPUT62), .A3(new_n1141), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1138), .A2(new_n1115), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n971), .B1(new_n1144), .B2(new_n1150), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n962), .A2(new_n702), .A3(new_n968), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n761), .A2(G2067), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n952), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n960), .A2(KEYINPUT46), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n952), .B1(new_n793), .B2(new_n953), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n960), .A2(KEYINPUT46), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(KEYINPUT125), .B(KEYINPUT47), .Z(new_n1159));
  XNOR2_X1  g734(.A(new_n1158), .B(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n965), .A2(new_n952), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(KEYINPUT48), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n963), .A2(new_n970), .A3(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1154), .A2(new_n1160), .A3(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(KEYINPUT126), .B1(new_n1151), .B2(new_n1164), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1044), .A2(new_n1049), .ZN(new_n1166));
  OR2_X1    g741(.A1(new_n1126), .A2(new_n1142), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT120), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1095), .A2(KEYINPUT120), .A3(new_n1097), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1150), .B(new_n1166), .C1(new_n1167), .C2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(new_n971), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1164), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT126), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1165), .A2(new_n1178), .ZN(G329));
  assign    G231 = 1'b0;
  AND4_X1   g754(.A1(G319), .A2(new_n641), .A3(new_n659), .A4(new_n660), .ZN(new_n1181));
  NAND2_X1  g755(.A1(new_n679), .A2(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g756(.A(new_n1182), .B(KEYINPUT127), .ZN(new_n1183));
  NAND2_X1  g757(.A1(new_n1183), .A2(new_n860), .ZN(new_n1184));
  NOR2_X1   g758(.A1(new_n1184), .A2(new_n939), .ZN(G308));
  NAND2_X1  g759(.A1(new_n932), .A2(new_n937), .ZN(new_n1186));
  NAND2_X1  g760(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n1187));
  NAND2_X1  g761(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g762(.A1(new_n1188), .A2(new_n860), .A3(new_n1183), .ZN(G225));
endmodule


