//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 0 0 1 0 1 0 0 1 0 0 1 1 0 1 1 0 1 0 0 1 0 0 0 1 0 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT77), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT75), .B1(new_n189), .B2(G119), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT75), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G128), .ZN(new_n193));
  AND2_X1   g007(.A1(new_n190), .A2(new_n193), .ZN(new_n194));
  AND3_X1   g008(.A1(new_n189), .A2(KEYINPUT74), .A3(G119), .ZN(new_n195));
  AOI21_X1  g009(.A(KEYINPUT74), .B1(new_n189), .B2(G119), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT24), .B(G110), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT76), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  OR2_X1    g014(.A1(KEYINPUT24), .A2(G110), .ZN(new_n201));
  NAND2_X1  g015(.A1(KEYINPUT24), .A2(G110), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(KEYINPUT76), .A3(new_n202), .ZN(new_n203));
  AOI22_X1  g017(.A1(new_n194), .A2(new_n197), .B1(new_n200), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n189), .A2(G119), .ZN(new_n205));
  OR2_X1    g019(.A1(new_n205), .A2(KEYINPUT23), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n192), .A2(G128), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(new_n205), .A3(KEYINPUT23), .ZN(new_n208));
  AOI21_X1  g022(.A(G110), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n188), .B1(new_n204), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n195), .ZN(new_n211));
  INV_X1    g025(.A(new_n196), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n211), .A2(new_n212), .A3(new_n190), .A4(new_n193), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n200), .A2(new_n203), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n206), .A2(new_n208), .ZN(new_n216));
  INV_X1    g030(.A(G110), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n215), .A2(KEYINPUT77), .A3(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(G125), .A2(G140), .ZN(new_n220));
  NOR2_X1   g034(.A1(G125), .A2(G140), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT16), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT16), .ZN(new_n223));
  INV_X1    g037(.A(G140), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n224), .A3(G125), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n222), .A2(G146), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT78), .ZN(new_n227));
  XNOR2_X1  g041(.A(new_n226), .B(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G125), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(new_n224), .ZN(new_n230));
  NAND2_X1  g044(.A1(G125), .A2(G140), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n210), .A2(new_n219), .A3(new_n228), .A4(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n223), .B1(new_n230), .B2(new_n231), .ZN(new_n236));
  INV_X1    g050(.A(new_n225), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n233), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n226), .ZN(new_n239));
  OAI221_X1 g053(.A(new_n239), .B1(new_n217), .B2(new_n216), .C1(new_n214), .C2(new_n213), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n235), .A2(KEYINPUT79), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(KEYINPUT79), .B1(new_n235), .B2(new_n240), .ZN(new_n242));
  INV_X1    g056(.A(G953), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(G221), .A3(G234), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n244), .B(KEYINPUT22), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n245), .B(G137), .ZN(new_n246));
  NOR3_X1   g060(.A1(new_n241), .A2(new_n242), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n246), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n248), .B1(new_n235), .B2(new_n240), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n187), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT25), .ZN(new_n251));
  INV_X1    g065(.A(G217), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n252), .B1(G234), .B2(new_n187), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT25), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n254), .B(new_n187), .C1(new_n247), .C2(new_n249), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n251), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  OR2_X1    g070(.A1(new_n247), .A2(new_n249), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n253), .A2(G902), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G137), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT65), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT65), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G137), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(KEYINPUT11), .A3(G134), .ZN(new_n266));
  INV_X1    g080(.A(G131), .ZN(new_n267));
  INV_X1    g081(.A(G134), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n268), .A2(G137), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT11), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n270), .B1(new_n268), .B2(G137), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n266), .B(new_n267), .C1(new_n269), .C2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n265), .A2(G134), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n269), .A2(KEYINPUT66), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT66), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n275), .B1(new_n268), .B2(G137), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(G131), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n272), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G143), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G146), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n189), .A2(KEYINPUT1), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT64), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n283), .B1(G143), .B2(new_n233), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n280), .A2(KEYINPUT64), .A3(G146), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n281), .B(new_n282), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT67), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n233), .A2(G143), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT64), .B1(new_n280), .B2(G146), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n283), .A2(new_n233), .A3(G143), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT67), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n292), .A3(new_n282), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n287), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n233), .A2(G143), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT1), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n296), .A2(G128), .B1(new_n281), .B2(new_n295), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(KEYINPUT69), .B1(new_n294), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT69), .ZN(new_n300));
  AOI211_X1 g114(.A(new_n300), .B(new_n297), .C1(new_n287), .C2(new_n293), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n279), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  AOI211_X1 g116(.A(new_n270), .B(new_n268), .C1(new_n262), .C2(new_n264), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n271), .A2(new_n269), .ZN(new_n304));
  OAI21_X1  g118(.A(G131), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n272), .ZN(new_n306));
  NAND2_X1  g120(.A1(KEYINPUT0), .A2(G128), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(KEYINPUT0), .A2(G128), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n281), .A2(new_n295), .ZN(new_n311));
  AOI22_X1  g125(.A1(new_n291), .A2(new_n308), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n302), .A2(KEYINPUT30), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT2), .ZN(new_n315));
  INV_X1    g129(.A(G113), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT68), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT68), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(KEYINPUT2), .A3(G113), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n315), .A2(new_n316), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(G116), .B(G119), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n320), .A2(new_n321), .A3(new_n323), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n272), .A2(new_n278), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n297), .B1(new_n287), .B2(new_n293), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n313), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT30), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n314), .A2(new_n327), .A3(new_n332), .ZN(new_n333));
  NOR2_X1   g147(.A1(G237), .A2(G953), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G210), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n335), .B(KEYINPUT71), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT26), .B(G101), .Z(new_n337));
  XNOR2_X1  g151(.A(new_n336), .B(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n338), .B(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n313), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n289), .A2(new_n290), .ZN(new_n342));
  AND4_X1   g156(.A1(new_n292), .A2(new_n342), .A3(new_n281), .A4(new_n282), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n292), .B1(new_n291), .B2(new_n282), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n298), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n300), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n294), .A2(KEYINPUT69), .A3(new_n298), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n341), .B1(new_n348), .B2(new_n279), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n320), .A2(new_n321), .A3(new_n323), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n323), .B1(new_n320), .B2(new_n321), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n340), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n333), .A2(new_n353), .A3(KEYINPUT31), .ZN(new_n354));
  AOI21_X1  g168(.A(KEYINPUT31), .B1(new_n333), .B2(new_n353), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT28), .B1(new_n349), .B2(new_n352), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n302), .A2(new_n352), .A3(new_n313), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT72), .ZN(new_n358));
  AOI22_X1  g172(.A1(new_n279), .A2(new_n345), .B1(new_n306), .B2(new_n312), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n358), .B1(new_n359), .B2(new_n352), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n330), .A2(KEYINPUT72), .A3(new_n327), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n357), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n356), .B1(KEYINPUT28), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n340), .ZN(new_n364));
  OAI22_X1  g178(.A1(new_n354), .A2(new_n355), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(G472), .A2(G902), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(KEYINPUT32), .A3(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT73), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n366), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n333), .A2(new_n353), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT31), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n333), .A2(new_n353), .A3(KEYINPUT31), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n362), .A2(KEYINPUT28), .ZN(new_n376));
  INV_X1    g190(.A(new_n356), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n340), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n370), .B1(new_n375), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(KEYINPUT73), .A3(KEYINPUT32), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n369), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT29), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n333), .A2(new_n357), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n340), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n383), .B(new_n385), .C1(new_n378), .C2(new_n340), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n340), .A2(new_n383), .ZN(new_n387));
  OR2_X1    g201(.A1(new_n349), .A2(new_n352), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n388), .A2(new_n357), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT28), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n377), .B(new_n387), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n386), .A2(new_n391), .A3(new_n187), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n365), .A2(new_n366), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT32), .ZN(new_n394));
  AOI22_X1  g208(.A1(new_n392), .A2(G472), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n260), .B1(new_n382), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G469), .ZN(new_n397));
  INV_X1    g211(.A(new_n291), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n296), .A2(G128), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n400), .B1(new_n343), .B2(new_n344), .ZN(new_n401));
  INV_X1    g215(.A(G104), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G107), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n402), .A2(G107), .ZN(new_n405));
  OAI21_X1  g219(.A(G101), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT3), .B1(new_n402), .B2(G107), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT3), .ZN(new_n408));
  INV_X1    g222(.A(G107), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n409), .A3(G104), .ZN(new_n410));
  INV_X1    g224(.A(G101), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n407), .A2(new_n410), .A3(new_n411), .A4(new_n403), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n406), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n401), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT10), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n407), .A2(new_n410), .A3(new_n403), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G101), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(KEYINPUT4), .A3(new_n412), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT4), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n416), .A2(new_n419), .A3(G101), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n414), .A2(new_n415), .B1(new_n422), .B2(new_n312), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n406), .A2(new_n412), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n424), .A2(new_n415), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n425), .B1(new_n299), .B2(new_n301), .ZN(new_n426));
  INV_X1    g240(.A(new_n306), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n423), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(G110), .B(G140), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n243), .A2(G227), .ZN(new_n430));
  XOR2_X1   g244(.A(new_n429), .B(new_n430), .Z(new_n431));
  OAI211_X1 g245(.A(new_n298), .B(new_n424), .C1(new_n343), .C2(new_n344), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n287), .A2(new_n293), .B1(new_n398), .B2(new_n399), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n432), .B1(new_n433), .B2(new_n424), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n434), .A2(KEYINPUT12), .A3(new_n306), .ZN(new_n435));
  AOI21_X1  g249(.A(KEYINPUT12), .B1(new_n434), .B2(new_n306), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n428), .B(new_n431), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n425), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n439), .B1(new_n346), .B2(new_n347), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n424), .B1(new_n294), .B2(new_n400), .ZN(new_n441));
  INV_X1    g255(.A(new_n312), .ZN(new_n442));
  OAI22_X1  g256(.A1(new_n441), .A2(KEYINPUT10), .B1(new_n442), .B2(new_n421), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n306), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n431), .B1(new_n444), .B2(new_n428), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n397), .B(new_n187), .C1(new_n438), .C2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n431), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n435), .A2(new_n436), .ZN(new_n448));
  NOR3_X1   g262(.A1(new_n440), .A2(new_n443), .A3(new_n306), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n444), .A2(new_n428), .A3(new_n431), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n450), .A2(G469), .A3(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n397), .A2(new_n187), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n446), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  XOR2_X1   g269(.A(KEYINPUT9), .B(G234), .Z(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n187), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n457), .A2(G221), .ZN(new_n458));
  XOR2_X1   g272(.A(new_n458), .B(KEYINPUT80), .Z(new_n459));
  NAND2_X1  g273(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT5), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(new_n192), .A3(G116), .ZN(new_n462));
  OAI211_X1 g276(.A(G113), .B(new_n462), .C1(new_n324), .C2(new_n461), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n413), .A2(new_n326), .A3(new_n463), .ZN(new_n464));
  XOR2_X1   g278(.A(G110), .B(G122), .Z(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n464), .B(new_n466), .C1(new_n421), .C2(new_n352), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT81), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n327), .A2(new_n420), .A3(new_n418), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT81), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n469), .A2(new_n470), .A3(new_n464), .A4(new_n466), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n294), .A2(new_n229), .A3(new_n298), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n312), .A2(new_n229), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT82), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT82), .B1(new_n312), .B2(new_n229), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n473), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT7), .ZN(new_n479));
  INV_X1    g293(.A(G224), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n480), .A2(G953), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n478), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  AOI22_X1  g296(.A1(new_n329), .A2(new_n229), .B1(new_n474), .B2(new_n475), .ZN(new_n483));
  INV_X1    g297(.A(new_n481), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n483), .A2(KEYINPUT7), .A3(new_n484), .A4(new_n477), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n463), .A2(new_n326), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n424), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n464), .ZN(new_n488));
  XOR2_X1   g302(.A(new_n465), .B(KEYINPUT8), .Z(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n472), .A2(new_n482), .A3(new_n485), .A4(new_n490), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n491), .A2(new_n187), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n466), .B1(new_n469), .B2(new_n464), .ZN(new_n493));
  OR2_X1    g307(.A1(new_n493), .A2(KEYINPUT6), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n493), .B1(new_n468), .B2(new_n471), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT6), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n478), .B(new_n481), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n492), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(G210), .B1(G237), .B2(G902), .ZN(new_n501));
  XOR2_X1   g315(.A(new_n501), .B(KEYINPUT83), .Z(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(G214), .B1(G237), .B2(G902), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n492), .A2(new_n499), .A3(new_n502), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n460), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n334), .A2(G143), .A3(G214), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(G143), .B1(new_n334), .B2(G214), .ZN(new_n511));
  OAI211_X1 g325(.A(KEYINPUT17), .B(G131), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(new_n238), .A3(new_n226), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT87), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n334), .A2(G214), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n280), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n517), .A2(new_n267), .A3(new_n509), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT85), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n509), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G131), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT17), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT85), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n517), .A2(new_n523), .A3(new_n267), .A4(new_n509), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n519), .A2(new_n521), .A3(new_n522), .A4(new_n524), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n512), .A2(new_n238), .A3(KEYINPUT87), .A4(new_n226), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n515), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  XOR2_X1   g341(.A(G113), .B(G122), .Z(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(KEYINPUT86), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(G104), .ZN(new_n530));
  OAI211_X1 g344(.A(KEYINPUT18), .B(G131), .C1(new_n520), .C2(KEYINPUT84), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n520), .A2(KEYINPUT84), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n232), .B(new_n233), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n520), .A2(KEYINPUT84), .A3(KEYINPUT18), .A4(G131), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n527), .A2(new_n530), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n530), .B1(new_n527), .B2(new_n536), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n187), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(G475), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n243), .A2(G952), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n542), .B1(G234), .B2(G237), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  AOI211_X1 g358(.A(new_n187), .B(new_n243), .C1(G234), .C2(G237), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  XOR2_X1   g360(.A(KEYINPUT21), .B(G898), .Z(new_n547));
  OAI21_X1  g361(.A(new_n544), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(KEYINPUT95), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n541), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT88), .ZN(new_n552));
  INV_X1    g366(.A(G116), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n552), .B1(new_n553), .B2(G122), .ZN(new_n554));
  INV_X1    g368(.A(G122), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(KEYINPUT88), .A3(G116), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n553), .A2(G122), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT14), .ZN(new_n559));
  OR3_X1    g373(.A1(new_n555), .A2(KEYINPUT14), .A3(G116), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n557), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(G107), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n557), .A2(new_n409), .A3(new_n558), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT90), .ZN(new_n564));
  XNOR2_X1  g378(.A(G128), .B(G143), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(new_n268), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT90), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n557), .A2(new_n567), .A3(new_n409), .A4(new_n558), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n562), .A2(new_n564), .A3(new_n566), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n565), .A2(KEYINPUT13), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n280), .A2(G128), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n570), .B(G134), .C1(KEYINPUT13), .C2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n189), .A2(G143), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n571), .A2(new_n573), .A3(new_n268), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT89), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT89), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n565), .A2(new_n576), .A3(new_n268), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n563), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n409), .B1(new_n557), .B2(new_n558), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n572), .B(new_n578), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n569), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n456), .A2(G217), .A3(new_n243), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT91), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT91), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n583), .B(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n569), .A2(new_n587), .A3(new_n581), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n585), .A2(new_n187), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(KEYINPUT92), .ZN(new_n590));
  INV_X1    g404(.A(G478), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(KEYINPUT15), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT92), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n585), .A2(new_n593), .A3(new_n187), .A4(new_n588), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n590), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT93), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n596), .B1(new_n589), .B2(new_n592), .ZN(new_n597));
  INV_X1    g411(.A(new_n589), .ZN(new_n598));
  INV_X1    g412(.A(new_n592), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(KEYINPUT93), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n595), .A2(new_n597), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT94), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n595), .A2(new_n600), .A3(KEYINPUT94), .A4(new_n597), .ZN(new_n604));
  INV_X1    g418(.A(G475), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n519), .A2(new_n521), .A3(new_n524), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n232), .B(KEYINPUT19), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n233), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n228), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n530), .B1(new_n609), .B2(new_n536), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n605), .B(new_n187), .C1(new_n537), .C2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(KEYINPUT20), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n527), .A2(new_n530), .A3(new_n536), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n536), .A2(new_n609), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n613), .B1(new_n614), .B2(new_n530), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT20), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n615), .A2(new_n616), .A3(new_n605), .A4(new_n187), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  AND4_X1   g432(.A1(new_n551), .A2(new_n603), .A3(new_n604), .A4(new_n618), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n508), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n396), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G101), .ZN(G3));
  NAND3_X1  g436(.A1(new_n590), .A2(new_n591), .A3(new_n594), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT33), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT96), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n582), .A2(new_n625), .A3(new_n587), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n581), .B(new_n569), .C1(new_n584), .C2(KEYINPUT96), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n624), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT33), .B1(new_n585), .B2(new_n588), .ZN(new_n629));
  OAI211_X1 g443(.A(G478), .B(new_n187), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n618), .A2(new_n540), .B1(new_n623), .B2(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n631), .A2(new_n504), .A3(new_n505), .A4(new_n506), .ZN(new_n632));
  OAI21_X1  g446(.A(KEYINPUT97), .B1(new_n632), .B2(new_n550), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n492), .A2(new_n499), .A3(new_n502), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n502), .B1(new_n492), .B2(new_n499), .ZN(new_n635));
  INV_X1    g449(.A(new_n505), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT97), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n637), .A2(new_n638), .A3(new_n549), .A4(new_n631), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n633), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(G902), .B1(new_n375), .B2(new_n379), .ZN(new_n641));
  INV_X1    g455(.A(G472), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n393), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n455), .A2(new_n256), .A3(new_n259), .A4(new_n459), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n640), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT34), .B(G104), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  NAND3_X1  g462(.A1(new_n612), .A2(KEYINPUT98), .A3(new_n617), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n649), .B1(KEYINPUT98), .B2(new_n617), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n603), .B2(new_n604), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n651), .A2(new_n551), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n645), .A2(new_n652), .A3(new_n637), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT35), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  INV_X1    g469(.A(new_n459), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n427), .B1(new_n423), .B2(new_n426), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n447), .B1(new_n449), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(G902), .B1(new_n658), .B2(new_n437), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n453), .B1(new_n659), .B2(new_n397), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n656), .B1(new_n660), .B2(new_n452), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n241), .A2(new_n242), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n248), .A2(KEYINPUT36), .ZN(new_n663));
  XOR2_X1   g477(.A(new_n662), .B(new_n663), .Z(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n258), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n256), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n661), .A2(new_n637), .A3(new_n619), .A4(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n667), .A2(new_n643), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT37), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G110), .ZN(G12));
  NAND2_X1  g484(.A1(new_n393), .A2(new_n394), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n392), .A2(G472), .ZN(new_n672));
  AOI21_X1  g486(.A(KEYINPUT73), .B1(new_n380), .B2(KEYINPUT32), .ZN(new_n673));
  AND4_X1   g487(.A1(KEYINPUT73), .A2(new_n365), .A3(KEYINPUT32), .A4(new_n366), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n671), .B(new_n672), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT99), .B(G900), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n543), .B1(new_n545), .B2(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n541), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n651), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n675), .A2(new_n679), .A3(new_n508), .A4(new_n666), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G128), .ZN(G30));
  NAND2_X1  g495(.A1(new_n389), .A2(new_n340), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n187), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n340), .B1(new_n333), .B2(new_n357), .ZN(new_n684));
  OAI21_X1  g498(.A(G472), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n671), .B(new_n685), .C1(new_n673), .C2(new_n674), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n686), .A2(new_n256), .A3(new_n505), .A4(new_n665), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n677), .B(KEYINPUT39), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n661), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT40), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n603), .A2(new_n604), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n618), .A2(new_n540), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n634), .A2(new_n635), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n695), .B(KEYINPUT38), .Z(new_n696));
  NOR4_X1   g510(.A1(new_n687), .A2(new_n691), .A3(new_n694), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(new_n280), .ZN(G45));
  NAND2_X1  g512(.A1(new_n623), .A2(new_n630), .ZN(new_n699));
  INV_X1    g513(.A(new_n677), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n693), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n661), .A2(new_n637), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n675), .A2(new_n666), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  INV_X1    g518(.A(new_n260), .ZN(new_n705));
  INV_X1    g519(.A(new_n446), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n659), .A2(new_n397), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n706), .A2(new_n707), .A3(new_n458), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n675), .A2(new_n640), .A3(new_n705), .A4(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT100), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT100), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n396), .A2(new_n711), .A3(new_n640), .A4(new_n708), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT41), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G113), .ZN(G15));
  NAND2_X1  g529(.A1(new_n708), .A2(new_n637), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n675), .A2(new_n652), .A3(new_n705), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G116), .ZN(G18));
  NAND4_X1  g533(.A1(new_n675), .A2(new_n619), .A3(new_n666), .A4(new_n717), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G119), .ZN(G21));
  AND2_X1   g535(.A1(new_n692), .A2(new_n693), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n708), .A2(new_n637), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n365), .A2(new_n187), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(G472), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n390), .B1(new_n388), .B2(new_n357), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n340), .B1(new_n726), .B2(new_n356), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n375), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n366), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n723), .A2(new_n705), .A3(new_n549), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  NAND4_X1  g546(.A1(new_n725), .A2(new_n666), .A3(new_n701), .A4(new_n729), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n716), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n229), .ZN(G27));
  INV_X1    g549(.A(new_n458), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n636), .B1(new_n504), .B2(new_n506), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT101), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n452), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n450), .A2(KEYINPUT101), .A3(G469), .A4(new_n451), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n739), .A2(new_n446), .A3(new_n454), .A4(new_n740), .ZN(new_n741));
  AND4_X1   g555(.A1(new_n736), .A2(new_n737), .A3(new_n701), .A4(new_n741), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n673), .A2(new_n674), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n672), .A2(new_n671), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n705), .B(new_n742), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT102), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT42), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n396), .A2(KEYINPUT102), .A3(new_n742), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n260), .B1(new_n395), .B2(new_n367), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(KEYINPUT42), .A3(new_n742), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G131), .ZN(G33));
  NAND2_X1  g568(.A1(new_n737), .A2(new_n736), .ZN(new_n755));
  INV_X1    g569(.A(new_n741), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n396), .A2(new_n679), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G134), .ZN(G36));
  NAND2_X1  g573(.A1(new_n450), .A2(new_n451), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT45), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(G469), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(KEYINPUT46), .A3(new_n454), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n763), .A2(KEYINPUT103), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(KEYINPUT103), .ZN(new_n765));
  AOI21_X1  g579(.A(KEYINPUT46), .B1(new_n762), .B2(new_n454), .ZN(new_n766));
  OR4_X1    g580(.A1(new_n706), .A2(new_n764), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n736), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n688), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(KEYINPUT104), .ZN(new_n770));
  INV_X1    g584(.A(new_n693), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n699), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT43), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n774), .A2(KEYINPUT105), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(KEYINPUT105), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n775), .A2(new_n643), .A3(new_n666), .A4(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT44), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n770), .A2(new_n737), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G137), .ZN(G39));
  XOR2_X1   g594(.A(new_n768), .B(KEYINPUT47), .Z(new_n781));
  NOR2_X1   g595(.A1(new_n675), .A2(new_n705), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n781), .A2(new_n701), .A3(new_n737), .A4(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G140), .ZN(G42));
  INV_X1    g598(.A(new_n696), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n260), .A2(new_n656), .A3(new_n636), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT106), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n686), .ZN(new_n789));
  INV_X1    g603(.A(new_n786), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n772), .B1(new_n790), .B2(KEYINPUT106), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n706), .A2(new_n707), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT49), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n788), .A2(new_n789), .A3(new_n791), .A4(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n792), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n755), .A2(new_n795), .A3(new_n544), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n774), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n751), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(KEYINPUT113), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT48), .ZN(new_n800));
  AND4_X1   g614(.A1(new_n705), .A2(new_n774), .A3(new_n543), .A4(new_n730), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n717), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n542), .B(KEYINPUT112), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n789), .A2(new_n705), .A3(new_n796), .ZN(new_n804));
  INV_X1    g618(.A(new_n631), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n800), .A2(new_n802), .A3(new_n803), .A4(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT114), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n795), .A2(new_n459), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n737), .B(new_n801), .C1(new_n781), .C2(new_n809), .ZN(new_n810));
  OR3_X1    g624(.A1(new_n804), .A2(new_n693), .A3(new_n699), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n801), .A2(new_n636), .A3(new_n696), .A4(new_n708), .ZN(new_n812));
  XOR2_X1   g626(.A(new_n812), .B(KEYINPUT50), .Z(new_n813));
  NAND3_X1  g627(.A1(new_n797), .A2(new_n666), .A3(new_n730), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n810), .A2(new_n811), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT51), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n637), .A2(new_n549), .A3(new_n631), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n818), .A2(new_n643), .A3(new_n644), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n396), .B2(new_n620), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT107), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n771), .A2(new_n549), .A3(new_n601), .ZN(new_n822));
  NOR4_X1   g636(.A1(new_n643), .A2(new_n644), .A3(new_n507), .A4(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n821), .B1(new_n823), .B2(new_n668), .ZN(new_n824));
  INV_X1    g638(.A(new_n822), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n645), .A2(new_n637), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n643), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(new_n508), .A3(new_n619), .A4(new_n666), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n826), .A2(new_n828), .A3(KEYINPUT107), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n820), .A2(new_n824), .A3(new_n829), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n460), .A2(new_n541), .A3(new_n650), .A4(new_n677), .ZN(new_n831));
  INV_X1    g645(.A(new_n737), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n601), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n675), .A2(new_n666), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n742), .A2(new_n730), .A3(new_n666), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n758), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n830), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n817), .B1(new_n837), .B2(KEYINPUT109), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n718), .A2(new_n720), .A3(new_n731), .ZN(new_n839));
  AOI221_X4 g653(.A(new_n839), .B1(new_n710), .B2(new_n712), .C1(new_n750), .C2(new_n752), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT109), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n841), .B1(new_n830), .B2(new_n836), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n838), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n694), .A2(new_n507), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n756), .A2(new_n666), .A3(new_n677), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n686), .A2(new_n736), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n734), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n680), .A2(new_n846), .A3(new_n703), .A4(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n679), .A2(new_n508), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n382), .A2(new_n395), .B1(new_n256), .B2(new_n665), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n734), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n853), .A2(KEYINPUT52), .A3(new_n703), .A4(new_n846), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT108), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n850), .A2(new_n854), .A3(KEYINPUT108), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(KEYINPUT110), .B1(new_n843), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n850), .A2(KEYINPUT108), .A3(new_n854), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT108), .B1(new_n850), .B2(new_n854), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT110), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n839), .B1(new_n712), .B2(new_n710), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n842), .A2(new_n753), .A3(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n864), .A2(new_n865), .A3(new_n838), .A4(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n840), .A2(new_n855), .A3(new_n837), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n817), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n860), .A2(new_n861), .A3(new_n868), .A4(new_n870), .ZN(new_n871));
  OR2_X1    g685(.A1(new_n871), .A2(KEYINPUT111), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n869), .A2(KEYINPUT53), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n840), .A2(new_n817), .A3(new_n837), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n873), .B1(new_n874), .B2(new_n859), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  AOI22_X1  g690(.A1(KEYINPUT111), .A2(new_n871), .B1(new_n876), .B2(KEYINPUT54), .ZN(new_n877));
  AND4_X1   g691(.A1(new_n808), .A2(new_n816), .A3(new_n872), .A4(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(G952), .A2(G953), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT115), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n794), .B1(new_n878), .B2(new_n880), .ZN(G75));
  NAND3_X1  g695(.A1(new_n860), .A2(new_n870), .A3(new_n868), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n882), .A2(G902), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n502), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT117), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n497), .B(new_n498), .ZN(new_n887));
  XOR2_X1   g701(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n888));
  XNOR2_X1  g702(.A(new_n887), .B(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT56), .ZN(new_n890));
  AOI22_X1  g704(.A1(new_n886), .A2(new_n889), .B1(new_n890), .B2(new_n884), .ZN(new_n891));
  AND4_X1   g705(.A1(KEYINPUT117), .A2(new_n884), .A3(new_n890), .A4(new_n889), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n243), .A2(G952), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(G51));
  NAND2_X1  g708(.A1(new_n882), .A2(KEYINPUT54), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n895), .A2(KEYINPUT118), .A3(new_n871), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT118), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n882), .A2(new_n897), .A3(KEYINPUT54), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n453), .B(KEYINPUT57), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT119), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n658), .A2(new_n437), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n896), .A2(KEYINPUT119), .A3(new_n898), .A4(new_n899), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n883), .A2(G469), .A3(new_n761), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n893), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT120), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT120), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n907), .A2(new_n911), .A3(new_n908), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n910), .A2(new_n912), .ZN(G54));
  NAND3_X1  g727(.A1(new_n883), .A2(KEYINPUT58), .A3(G475), .ZN(new_n914));
  INV_X1    g728(.A(new_n615), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT121), .ZN(new_n917));
  AOI211_X1 g731(.A(new_n893), .B(new_n917), .C1(new_n915), .C2(new_n914), .ZN(G60));
  OR2_X1    g732(.A1(new_n628), .A2(new_n629), .ZN(new_n919));
  NAND2_X1  g733(.A1(G478), .A2(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT59), .Z(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n896), .A2(new_n919), .A3(new_n898), .A4(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n921), .B1(new_n877), .B2(new_n872), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n908), .B(new_n923), .C1(new_n924), .C2(new_n919), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(G63));
  NAND2_X1  g740(.A1(G217), .A2(G902), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT60), .Z(new_n928));
  NAND2_X1  g742(.A1(new_n882), .A2(new_n928), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n257), .B(KEYINPUT123), .Z(new_n930));
  AOI21_X1  g744(.A(new_n893), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n882), .A2(new_n664), .A3(new_n928), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n931), .A2(KEYINPUT61), .A3(new_n932), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n932), .A2(KEYINPUT122), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(KEYINPUT122), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n934), .A2(new_n931), .A3(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT124), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n937), .B1(new_n936), .B2(new_n938), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n933), .B1(new_n939), .B2(new_n940), .ZN(G66));
  INV_X1    g755(.A(new_n830), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n866), .A2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT125), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n243), .B1(new_n547), .B2(G224), .ZN(new_n945));
  AOI22_X1  g759(.A1(new_n943), .A2(new_n243), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n946), .B1(new_n944), .B2(new_n945), .ZN(new_n947));
  INV_X1    g761(.A(new_n497), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n948), .B1(G898), .B2(new_n243), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n947), .B(new_n949), .ZN(G69));
  AND3_X1   g764(.A1(new_n779), .A2(new_n783), .A3(new_n758), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n853), .A2(new_n703), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n753), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n770), .A2(new_n844), .A3(new_n751), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n951), .A2(KEYINPUT126), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n779), .A2(new_n956), .A3(new_n783), .A4(new_n758), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n958), .B1(new_n959), .B2(new_n954), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n957), .A2(new_n960), .A3(new_n243), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n314), .A2(new_n332), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(new_n607), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(G900), .A2(G953), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n961), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n697), .A2(new_n952), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT62), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n690), .A2(new_n832), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n771), .A2(new_n601), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n396), .B(new_n969), .C1(new_n631), .C2(new_n970), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n779), .A2(new_n783), .A3(new_n968), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n243), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n963), .ZN(new_n974));
  AOI21_X1  g788(.A(KEYINPUT127), .B1(new_n966), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(G227), .B1(new_n964), .B2(KEYINPUT127), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n243), .B1(new_n977), .B2(G900), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n975), .B(new_n978), .ZN(G72));
  NAND2_X1  g793(.A1(G472), .A2(G902), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT63), .Z(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(new_n972), .B2(new_n943), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n684), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n385), .A2(new_n371), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n876), .A2(new_n981), .A3(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n983), .A2(new_n908), .A3(new_n985), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n957), .A2(new_n960), .A3(new_n866), .A4(new_n942), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n384), .B1(new_n987), .B2(new_n981), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n986), .B1(new_n988), .B2(new_n340), .ZN(G57));
endmodule


