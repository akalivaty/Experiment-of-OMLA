//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n823, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932;
  INV_X1    g000(.A(G218gat), .ZN(new_n202));
  INV_X1    g001(.A(G43gat), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT15), .B1(new_n203), .B2(G50gat), .ZN(new_n204));
  AOI21_X1  g003(.A(new_n204), .B1(new_n203), .B2(G50gat), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n203), .A2(G50gat), .ZN(new_n206));
  XOR2_X1   g005(.A(KEYINPUT91), .B(G50gat), .Z(new_n207));
  OAI21_X1  g006(.A(new_n206), .B1(new_n207), .B2(G43gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT15), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n205), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G29gat), .ZN(new_n211));
  INV_X1    g010(.A(G36gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  OR4_X1    g013(.A1(KEYINPUT92), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(G29gat), .A2(G36gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n216), .B(KEYINPUT14), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT92), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n210), .A2(new_n214), .A3(new_n215), .A4(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n205), .B1(new_n217), .B2(new_n213), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(KEYINPUT17), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT99), .B(G85gat), .ZN(new_n223));
  INV_X1    g022(.A(G92gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G85gat), .A2(G92gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n226), .B(KEYINPUT7), .ZN(new_n227));
  INV_X1    g026(.A(G99gat), .ZN(new_n228));
  INV_X1    g027(.A(G106gat), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT8), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n225), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G99gat), .B(G106gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n231), .B(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n222), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n233), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G190gat), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n238), .A2(G190gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n202), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n241), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n243), .A2(G218gat), .A3(new_n239), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT98), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n242), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G134gat), .B(G162gat), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n247), .B(new_n248), .Z(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n242), .A2(new_n244), .A3(new_n245), .A4(new_n249), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G8gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(G15gat), .B(G22gat), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT16), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n256), .B1(new_n257), .B2(G1gat), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT93), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n255), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n258), .B1(G1gat), .B2(new_n256), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(KEYINPUT96), .B1(G71gat), .B2(G78gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(G57gat), .B(G64gat), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  XOR2_X1   g065(.A(G71gat), .B(G78gat), .Z(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n262), .B1(KEYINPUT21), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(KEYINPUT97), .ZN(new_n270));
  NAND2_X1  g069(.A1(G231gat), .A2(G233gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n268), .A2(KEYINPUT21), .ZN(new_n273));
  XOR2_X1   g072(.A(G127gat), .B(G155gat), .Z(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n272), .B(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n277));
  XNOR2_X1  g076(.A(G183gat), .B(G211gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n276), .B(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n254), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT100), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n231), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(new_n233), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT10), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n233), .A2(KEYINPUT10), .A3(new_n268), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G230gat), .A2(G233gat), .ZN(new_n290));
  AND2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n285), .A2(new_n290), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT101), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n292), .A2(KEYINPUT101), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G176gat), .B(G204gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(G148gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n297), .B(KEYINPUT102), .ZN(new_n298));
  INV_X1    g097(.A(G120gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n293), .A2(new_n300), .A3(new_n294), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n281), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(G141gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n306), .A2(G148gat), .ZN(new_n307));
  INV_X1    g106(.A(G148gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n308), .A2(G141gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(G155gat), .A2(G162gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312));
  OAI22_X1  g111(.A1(new_n307), .A2(new_n309), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT77), .ZN(new_n314));
  INV_X1    g113(.A(G155gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(KEYINPUT77), .A2(G155gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(G162gat), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n313), .B1(KEYINPUT2), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(KEYINPUT76), .A2(KEYINPUT2), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n308), .A2(G141gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n306), .A2(G148gat), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT76), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n310), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(KEYINPUT76), .A2(G155gat), .A3(G162gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NOR3_X1   g127(.A1(new_n324), .A2(new_n328), .A3(new_n312), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT3), .B1(new_n319), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n299), .A2(G113gat), .ZN(new_n331));
  INV_X1    g130(.A(G113gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G120gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  AND2_X1   g133(.A1(G127gat), .A2(G134gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(G127gat), .A2(G134gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NOR3_X1   g136(.A1(KEYINPUT66), .A2(KEYINPUT67), .A3(KEYINPUT1), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n334), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(G127gat), .ZN(new_n340));
  INV_X1    g139(.A(G134gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT1), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT66), .ZN(new_n344));
  NAND2_X1  g143(.A1(G127gat), .A2(G134gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n342), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G113gat), .B(G120gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI22_X1  g147(.A1(new_n335), .A2(new_n336), .B1(KEYINPUT67), .B2(KEYINPUT1), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n339), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n318), .A2(KEYINPUT2), .ZN(new_n351));
  INV_X1    g150(.A(G162gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n315), .A2(new_n352), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n322), .A2(new_n323), .B1(new_n353), .B2(new_n310), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT3), .ZN(new_n356));
  AND3_X1   g155(.A1(KEYINPUT76), .A2(G155gat), .A3(G162gat), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT76), .B1(G155gat), .B2(G162gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G141gat), .B(G148gat), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n359), .B(new_n353), .C1(new_n360), .C2(new_n321), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n355), .A2(new_n356), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n330), .A2(new_n350), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G225gat), .A2(G233gat), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n339), .A2(new_n348), .A3(new_n349), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n365), .A2(new_n355), .A3(new_n361), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT4), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n322), .A2(new_n323), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n312), .B1(new_n369), .B2(new_n320), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n370), .A2(new_n359), .B1(new_n351), .B2(new_n354), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n371), .A2(KEYINPUT4), .A3(new_n365), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n363), .A2(new_n364), .A3(new_n368), .A4(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(KEYINPUT78), .A2(KEYINPUT5), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AND3_X1   g174(.A1(new_n371), .A2(KEYINPUT4), .A3(new_n365), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT4), .B1(new_n371), .B2(new_n365), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n374), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n378), .A2(new_n364), .A3(new_n363), .A4(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT79), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n355), .A2(new_n361), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n350), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n366), .ZN(new_n385));
  INV_X1    g184(.A(new_n364), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n382), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI211_X1 g186(.A(KEYINPUT79), .B(new_n364), .C1(new_n384), .C2(new_n366), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT5), .ZN(new_n389));
  NOR3_X1   g188(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n381), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT86), .ZN(new_n392));
  XNOR2_X1  g191(.A(KEYINPUT0), .B(G57gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(G85gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(G1gat), .B(G29gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n391), .A2(new_n392), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n366), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n365), .B1(new_n355), .B2(new_n361), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n386), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT79), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n382), .A3(new_n386), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(KEYINPUT5), .A3(new_n402), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n403), .A2(new_n396), .A3(new_n375), .A4(new_n380), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT86), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n397), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n403), .A2(new_n375), .A3(new_n380), .ZN(new_n408));
  INV_X1    g207(.A(new_n396), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(G211gat), .A2(G218gat), .ZN(new_n412));
  OR2_X1    g211(.A1(G211gat), .A2(G218gat), .ZN(new_n413));
  AND2_X1   g212(.A1(G197gat), .A2(G204gat), .ZN(new_n414));
  NOR2_X1   g213(.A1(G197gat), .A2(G204gat), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT22), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n412), .B(new_n413), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G211gat), .B(G218gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n412), .A2(new_n417), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n419), .B(new_n420), .C1(new_n415), .C2(new_n414), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(G226gat), .A2(G233gat), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(G183gat), .A2(G190gat), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT64), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(G183gat), .A2(G190gat), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT24), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n428), .A2(new_n431), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  AND2_X1   g233(.A1(G169gat), .A2(G176gat), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT23), .ZN(new_n436));
  INV_X1    g235(.A(G169gat), .ZN(new_n437));
  INV_X1    g236(.A(G176gat), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n435), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n434), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT25), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AND3_X1   g243(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n426), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n443), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n441), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n444), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n437), .A2(new_n438), .A3(KEYINPUT26), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT26), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n453), .B1(G169gat), .B2(G176gat), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n452), .B(new_n429), .C1(new_n454), .C2(new_n435), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(G183gat), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n457), .A2(KEYINPUT27), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT27), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n459), .A2(G183gat), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT65), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n459), .A2(G183gat), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT65), .ZN(new_n463));
  AOI21_X1  g262(.A(G190gat), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT28), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT28), .ZN(new_n466));
  NOR4_X1   g265(.A1(new_n458), .A2(new_n460), .A3(new_n466), .A4(G190gat), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n456), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(KEYINPUT73), .B(KEYINPUT29), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n425), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n424), .B1(new_n451), .B2(new_n468), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n423), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n472), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT29), .B1(new_n451), .B2(new_n468), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n474), .B(new_n422), .C1(new_n425), .C2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G8gat), .B(G36gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(G92gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n479), .B(KEYINPUT74), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n480), .B(G64gat), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n477), .A2(KEYINPUT37), .ZN(new_n484));
  XOR2_X1   g283(.A(KEYINPUT89), .B(KEYINPUT37), .Z(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n484), .B(new_n482), .C1(new_n477), .C2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n483), .B1(new_n487), .B2(KEYINPUT38), .ZN(new_n488));
  INV_X1    g287(.A(new_n407), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n404), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n469), .A2(new_n470), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n472), .B1(new_n492), .B2(new_n424), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n422), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT88), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n475), .A2(new_n425), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n423), .B1(new_n496), .B2(new_n472), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT88), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n493), .A2(new_n498), .A3(new_n422), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n495), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT37), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT38), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n477), .A2(new_n486), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n503), .A2(new_n481), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n501), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n411), .A2(new_n488), .A3(new_n491), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(G228gat), .A2(G233gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n422), .A2(new_n470), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n371), .B1(new_n508), .B2(new_n356), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n422), .B1(new_n362), .B2(new_n470), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n507), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT29), .B1(new_n418), .B2(new_n421), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n383), .B1(new_n513), .B2(KEYINPUT3), .ZN(new_n514));
  INV_X1    g313(.A(new_n470), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n515), .B1(new_n371), .B2(new_n356), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n512), .B(new_n514), .C1(new_n516), .C2(new_n422), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT84), .ZN(new_n518));
  INV_X1    g317(.A(G22gat), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n511), .B(new_n517), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(KEYINPUT31), .B(G50gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT82), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(G78gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(new_n229), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n511), .A2(new_n517), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(G22gat), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n520), .B(new_n525), .C1(new_n527), .C2(new_n518), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n511), .A2(new_n517), .A3(new_n519), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT83), .B1(new_n530), .B2(new_n524), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n511), .A2(new_n519), .A3(new_n517), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n519), .B1(new_n511), .B2(new_n517), .ZN(new_n533));
  OAI211_X1 g332(.A(KEYINPUT83), .B(new_n524), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n528), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n363), .A2(new_n368), .A3(new_n372), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n386), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT85), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT85), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n537), .A2(new_n540), .A3(new_n386), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT39), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n384), .A2(new_n364), .A3(new_n366), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n539), .A2(KEYINPUT39), .A3(new_n541), .A4(new_n545), .ZN(new_n546));
  OR2_X1    g345(.A1(KEYINPUT87), .A2(KEYINPUT40), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n544), .A2(new_n409), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(KEYINPUT87), .A2(KEYINPUT40), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n396), .B1(new_n542), .B2(new_n543), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n551), .A2(KEYINPUT87), .A3(KEYINPUT40), .A4(new_n546), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT30), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n553), .B1(new_n477), .B2(new_n482), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n473), .A2(new_n476), .A3(new_n481), .A4(KEYINPUT30), .ZN(new_n555));
  AOI211_X1 g354(.A(KEYINPUT75), .B(new_n481), .C1(new_n473), .C2(new_n476), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT75), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n557), .B1(new_n477), .B2(new_n482), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n554), .B(new_n555), .C1(new_n556), .C2(new_n558), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n550), .A2(new_n552), .A3(new_n406), .A4(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n506), .A2(new_n536), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n536), .ZN(new_n562));
  INV_X1    g361(.A(new_n404), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n563), .B1(new_n410), .B2(KEYINPUT81), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n409), .B1(new_n381), .B2(new_n390), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(new_n489), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT81), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n490), .B1(new_n564), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n562), .B1(new_n569), .B2(new_n559), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n339), .A2(new_n348), .A3(KEYINPUT68), .A4(new_n349), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT68), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n365), .A2(new_n572), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n443), .A2(new_n442), .B1(new_n449), .B2(new_n441), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n457), .A2(KEYINPUT27), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n463), .B1(new_n462), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n463), .B1(new_n457), .B2(KEYINPUT27), .ZN(new_n577));
  INV_X1    g376(.A(G190gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n466), .B1(new_n576), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n458), .A2(new_n460), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n581), .A2(KEYINPUT28), .A3(new_n578), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n455), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n571), .B(new_n573), .C1(new_n574), .C2(new_n583), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n451), .A2(new_n468), .A3(KEYINPUT68), .A4(new_n350), .ZN(new_n585));
  INV_X1    g384(.A(G227gat), .ZN(new_n586));
  INV_X1    g385(.A(G233gat), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n584), .A2(new_n585), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT32), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT69), .B(KEYINPUT33), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n593));
  XNOR2_X1  g392(.A(G15gat), .B(G43gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G71gat), .B(G99gat), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n590), .A2(new_n592), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n597), .ZN(new_n599));
  OAI211_X1 g398(.A(new_n589), .B(KEYINPUT32), .C1(new_n591), .C2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT72), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n584), .A2(new_n585), .ZN(new_n603));
  INV_X1    g402(.A(new_n588), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT34), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n603), .A2(KEYINPUT34), .A3(new_n604), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n601), .A2(new_n602), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n607), .A2(KEYINPUT72), .A3(new_n608), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT34), .B1(new_n603), .B2(new_n604), .ZN(new_n612));
  AOI211_X1 g411(.A(new_n606), .B(new_n588), .C1(new_n584), .C2(new_n585), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n602), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n611), .A2(new_n614), .A3(new_n600), .A4(new_n598), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT36), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n561), .A2(new_n570), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT35), .ZN(new_n619));
  INV_X1    g418(.A(new_n559), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n566), .B1(new_n405), .B2(new_n397), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n620), .B1(new_n621), .B2(new_n490), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n536), .A2(new_n616), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n619), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n564), .A2(new_n568), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n559), .B1(new_n625), .B2(new_n491), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT90), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n627), .B1(new_n536), .B2(new_n616), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n536), .A2(new_n627), .A3(new_n616), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n626), .B(KEYINPUT35), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n618), .A2(new_n624), .A3(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n221), .A2(new_n262), .ZN(new_n632));
  INV_X1    g431(.A(new_n262), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n632), .B1(new_n222), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G229gat), .A2(G233gat), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT18), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n221), .B(new_n262), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n635), .B(KEYINPUT94), .Z(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n641), .B(KEYINPUT95), .Z(new_n642));
  NAND2_X1  g441(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT11), .B(G169gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(G197gat), .ZN(new_n645));
  XOR2_X1   g444(.A(G113gat), .B(G141gat), .Z(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT12), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n643), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n637), .A2(new_n648), .A3(new_n642), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n631), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n305), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n569), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n559), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n658), .B1(new_n257), .B2(new_n255), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n659), .B1(new_n257), .B2(new_n255), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT42), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n658), .A2(G8gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT103), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(G1325gat));
  AOI21_X1  g463(.A(new_n654), .B1(new_n610), .B2(new_n615), .ZN(new_n665));
  INV_X1    g464(.A(new_n617), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n655), .A2(new_n666), .ZN(new_n667));
  MUX2_X1   g466(.A(new_n665), .B(new_n667), .S(G15gat), .Z(G1326gat));
  NOR2_X1   g467(.A1(new_n654), .A2(new_n536), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT43), .B(G22gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT104), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n669), .B(new_n671), .ZN(G1327gat));
  INV_X1    g471(.A(KEYINPUT106), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT35), .B1(new_n629), .B2(new_n628), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n625), .A2(new_n491), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n620), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n624), .B(new_n673), .C1(new_n674), .C2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n673), .B1(new_n630), .B2(new_n624), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n618), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n680), .A2(new_n681), .A3(new_n253), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT107), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n631), .A2(new_n253), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n683), .B1(new_n684), .B2(KEYINPUT44), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n652), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n304), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n280), .B(KEYINPUT105), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n680), .A2(new_n683), .A3(new_n681), .A4(new_n253), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n686), .A2(new_n688), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT108), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(new_n693));
  OR3_X1    g492(.A1(new_n693), .A2(KEYINPUT109), .A3(new_n675), .ZN(new_n694));
  OAI21_X1  g493(.A(KEYINPUT109), .B1(new_n693), .B2(new_n675), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(G29gat), .A3(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n280), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n254), .A2(new_n304), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n653), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n700), .A2(new_n211), .A3(new_n569), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT45), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n696), .A2(new_n702), .ZN(G1328gat));
  OAI21_X1  g502(.A(G36gat), .B1(new_n693), .B2(new_n620), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n699), .A2(G36gat), .A3(new_n620), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT46), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(G1329gat));
  OR3_X1    g506(.A1(new_n691), .A2(KEYINPUT112), .A3(new_n617), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT112), .B1(new_n691), .B2(new_n617), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n708), .A2(G43gat), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n700), .A2(new_n203), .A3(new_n616), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(KEYINPUT47), .A3(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT111), .ZN(new_n713));
  OR2_X1    g512(.A1(new_n691), .A2(KEYINPUT108), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n691), .A2(KEYINPUT108), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n617), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n713), .B1(new_n716), .B2(new_n203), .ZN(new_n717));
  OAI211_X1 g516(.A(KEYINPUT111), .B(G43gat), .C1(new_n693), .C2(new_n617), .ZN(new_n718));
  AND3_X1   g517(.A1(new_n717), .A2(new_n711), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n712), .B1(new_n719), .B2(new_n720), .ZN(G1330gat));
  INV_X1    g520(.A(new_n207), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(new_n691), .B2(new_n536), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n699), .A2(new_n536), .A3(new_n722), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n723), .A2(KEYINPUT48), .A3(new_n725), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n693), .A2(new_n536), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n724), .B1(new_n727), .B2(new_n722), .ZN(new_n728));
  XNOR2_X1  g527(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n726), .B1(new_n728), .B2(new_n729), .ZN(G1331gat));
  NOR2_X1   g529(.A1(new_n281), .A2(new_n652), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n731), .A2(new_n304), .A3(new_n680), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT114), .Z(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n569), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n559), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n737));
  XOR2_X1   g536(.A(KEYINPUT49), .B(G64gat), .Z(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n736), .B2(new_n738), .ZN(G1333gat));
  NAND3_X1  g538(.A1(new_n733), .A2(G71gat), .A3(new_n666), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n733), .A2(new_n616), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n741), .B2(G71gat), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g542(.A1(new_n733), .A2(new_n562), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(G78gat), .ZN(G1335gat));
  INV_X1    g544(.A(new_n304), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n280), .A2(new_n652), .A3(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n686), .A2(new_n690), .A3(new_n747), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n748), .A2(new_n675), .A3(new_n223), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n280), .A2(new_n652), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n680), .A2(new_n253), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT51), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT51), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n680), .A2(new_n753), .A3(new_n253), .A4(new_n750), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n304), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n569), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n749), .B1(new_n758), .B2(new_n223), .ZN(G1336gat));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n757), .A2(new_n224), .A3(new_n559), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(G92gat), .B1(new_n748), .B2(new_n620), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n763), .B(new_n765), .ZN(G1337gat));
  OAI21_X1  g565(.A(G99gat), .B1(new_n748), .B2(new_n617), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n616), .A2(new_n228), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n767), .B1(new_n756), .B2(new_n768), .ZN(G1338gat));
  NAND4_X1  g568(.A1(new_n686), .A2(new_n562), .A3(new_n690), .A4(new_n747), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(G106gat), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n752), .A2(new_n229), .A3(new_n304), .A4(new_n754), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n771), .B(new_n772), .C1(new_n536), .C2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT116), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n770), .A2(new_n775), .A3(G106gat), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n776), .A2(KEYINPUT53), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n771), .B(KEYINPUT116), .C1(new_n536), .C2(new_n773), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT117), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n779), .B1(new_n777), .B2(new_n778), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n774), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT118), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  OAI211_X1 g583(.A(KEYINPUT118), .B(new_n774), .C1(new_n780), .C2(new_n781), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(G1339gat));
  NOR2_X1   g585(.A1(new_n629), .A2(new_n628), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n634), .A2(new_n635), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n638), .A2(new_n640), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n647), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n651), .A2(new_n790), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n253), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n300), .B1(new_n291), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(KEYINPUT54), .B1(new_n289), .B2(new_n290), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n291), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n794), .B(KEYINPUT55), .C1(new_n291), .C2(new_n795), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n798), .A2(new_n303), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT119), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n798), .A2(KEYINPUT119), .A3(new_n303), .A4(new_n799), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n792), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n802), .A2(new_n652), .A3(new_n803), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n304), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n253), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n689), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n281), .A2(new_n652), .A3(new_n304), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n787), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n569), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(new_n559), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n814), .A2(new_n332), .A3(new_n652), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n623), .B1(new_n809), .B2(new_n811), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n816), .A2(new_n569), .A3(new_n620), .ZN(new_n817));
  OAI21_X1  g616(.A(G113gat), .B1(new_n817), .B2(new_n687), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n815), .A2(new_n818), .ZN(G1340gat));
  INV_X1    g618(.A(new_n813), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n746), .A2(new_n559), .ZN(new_n821));
  AOI21_X1  g620(.A(G120gat), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n817), .A2(new_n299), .A3(new_n746), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n822), .A2(new_n823), .ZN(G1341gat));
  NOR3_X1   g623(.A1(new_n817), .A2(new_n340), .A3(new_n689), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n814), .A2(new_n280), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n825), .B1(new_n826), .B2(new_n340), .ZN(G1342gat));
  NOR4_X1   g626(.A1(new_n813), .A2(G134gat), .A3(new_n559), .A4(new_n254), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT56), .ZN(new_n829));
  OR2_X1    g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  OAI21_X1  g630(.A(G134gat), .B1(new_n817), .B2(new_n254), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(G1343gat));
  NAND2_X1  g632(.A1(new_n792), .A2(new_n804), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n807), .B1(new_n687), .B2(new_n800), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n254), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n280), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  OAI211_X1 g636(.A(KEYINPUT57), .B(new_n562), .C1(new_n837), .C2(new_n810), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n536), .B1(new_n809), .B2(new_n811), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n838), .B1(new_n839), .B2(KEYINPUT57), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n666), .A2(new_n675), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n842), .A2(new_n559), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n840), .A2(new_n652), .A3(new_n843), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n844), .A2(KEYINPUT121), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(KEYINPUT121), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n845), .A2(new_n846), .A3(G141gat), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT58), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n839), .A2(new_n843), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n306), .A3(new_n652), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n847), .A2(new_n848), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n844), .A2(G141gat), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n851), .ZN(new_n854));
  AOI21_X1  g653(.A(KEYINPUT120), .B1(new_n854), .B2(KEYINPUT58), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n854), .A2(KEYINPUT120), .A3(KEYINPUT58), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n852), .B1(new_n855), .B2(new_n856), .ZN(G1344gat));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n840), .A2(new_n843), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n858), .B(G148gat), .C1(new_n859), .C2(new_n746), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT122), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n809), .A2(new_n811), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT57), .B1(new_n862), .B2(new_n536), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864));
  INV_X1    g663(.A(new_n800), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n792), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n280), .B1(new_n866), .B2(new_n836), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n864), .B(new_n562), .C1(new_n867), .C2(new_n810), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n863), .A2(new_n304), .A3(new_n843), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(G148gat), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n861), .B1(new_n870), .B2(KEYINPUT59), .ZN(new_n871));
  AOI211_X1 g670(.A(KEYINPUT122), .B(new_n858), .C1(new_n869), .C2(G148gat), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n860), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n839), .A2(new_n308), .A3(new_n821), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(new_n842), .B2(new_n874), .ZN(G1345gat));
  NAND2_X1  g674(.A1(new_n316), .A2(new_n317), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n859), .A2(new_n876), .A3(new_n689), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n850), .A2(new_n280), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n876), .B2(new_n878), .ZN(G1346gat));
  NOR3_X1   g678(.A1(new_n859), .A2(new_n352), .A3(new_n254), .ZN(new_n880));
  AOI21_X1  g679(.A(G162gat), .B1(new_n850), .B2(new_n253), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n880), .A2(new_n881), .ZN(G1347gat));
  NOR2_X1   g681(.A1(new_n569), .A2(new_n620), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n812), .A2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n437), .A3(new_n652), .ZN(new_n886));
  XOR2_X1   g685(.A(new_n883), .B(KEYINPUT123), .Z(new_n887));
  NAND2_X1  g686(.A1(new_n816), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(G169gat), .B1(new_n888), .B2(new_n687), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n886), .A2(new_n889), .ZN(G1348gat));
  NOR3_X1   g689(.A1(new_n888), .A2(new_n438), .A3(new_n746), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n438), .B1(new_n884), .B2(new_n746), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT124), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n893), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n891), .B1(new_n894), .B2(new_n895), .ZN(G1349gat));
  OAI21_X1  g695(.A(G183gat), .B1(new_n888), .B2(new_n689), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n280), .A2(new_n581), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n884), .B2(new_n898), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g699(.A1(new_n885), .A2(new_n578), .A3(new_n253), .ZN(new_n901));
  OAI21_X1  g700(.A(G190gat), .B1(new_n888), .B2(new_n254), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n902), .A2(KEYINPUT61), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n902), .A2(KEYINPUT61), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n901), .B1(new_n903), .B2(new_n904), .ZN(G1351gat));
  NAND2_X1  g704(.A1(new_n887), .A2(new_n617), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n868), .B(new_n907), .C1(new_n839), .C2(new_n864), .ZN(new_n908));
  OAI21_X1  g707(.A(G197gat), .B1(new_n908), .B2(new_n687), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n839), .A2(new_n617), .A3(new_n883), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n910), .A2(G197gat), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n909), .B1(new_n911), .B2(new_n687), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT125), .ZN(G1352gat));
  NOR3_X1   g712(.A1(new_n910), .A2(G204gat), .A3(new_n746), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT62), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n863), .A2(new_n304), .A3(new_n868), .ZN(new_n916));
  OAI21_X1  g715(.A(G204gat), .B1(new_n916), .B2(new_n906), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(G1353gat));
  OAI21_X1  g717(.A(G211gat), .B1(new_n908), .B2(new_n697), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT126), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT63), .ZN(new_n921));
  OR3_X1    g720(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n919), .A2(new_n921), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(KEYINPUT127), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n920), .B1(new_n919), .B2(new_n921), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT127), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n919), .A2(new_n926), .A3(new_n921), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n922), .A2(new_n924), .A3(new_n925), .A4(new_n927), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n697), .A2(G211gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n928), .B1(new_n910), .B2(new_n929), .ZN(G1354gat));
  OAI21_X1  g729(.A(G218gat), .B1(new_n908), .B2(new_n254), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n253), .A2(new_n202), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n910), .B2(new_n932), .ZN(G1355gat));
endmodule


