//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT75), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT22), .B(G137), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  OR2_X1    g005(.A1(KEYINPUT66), .A2(G128), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT66), .A2(G128), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n192), .A2(KEYINPUT23), .A3(G119), .A4(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n195));
  INV_X1    g009(.A(G119), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n195), .B1(new_n196), .B2(G128), .ZN(new_n197));
  AOI21_X1  g011(.A(KEYINPUT72), .B1(new_n196), .B2(G128), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n194), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT66), .A2(G128), .ZN(new_n200));
  NOR2_X1   g014(.A1(KEYINPUT66), .A2(G128), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n202), .A2(KEYINPUT72), .A3(KEYINPUT23), .A4(G119), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n199), .A2(G110), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(G119), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n196), .A2(G128), .ZN(new_n206));
  XOR2_X1   g020(.A(KEYINPUT24), .B(G110), .Z(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  INV_X1    g023(.A(G140), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G125), .ZN(new_n211));
  INV_X1    g025(.A(G125), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G140), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n211), .A2(new_n213), .A3(KEYINPUT73), .A4(KEYINPUT16), .ZN(new_n214));
  AND3_X1   g028(.A1(new_n211), .A2(new_n213), .A3(KEYINPUT16), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT73), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n216), .B1(new_n211), .B2(KEYINPUT16), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n209), .B(new_n214), .C1(new_n215), .C2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n211), .A2(new_n213), .A3(KEYINPUT16), .ZN(new_n220));
  OR3_X1    g034(.A1(new_n212), .A2(KEYINPUT16), .A3(G140), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(new_n216), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n209), .B1(new_n222), .B2(new_n214), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n204), .B(new_n208), .C1(new_n219), .C2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n214), .B1(new_n215), .B2(new_n217), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G146), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n211), .A2(new_n213), .A3(new_n209), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT74), .B(G110), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n228), .B1(new_n199), .B2(new_n203), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n207), .B1(new_n205), .B2(new_n206), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n226), .B(new_n227), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT76), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n224), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n232), .B1(new_n224), .B2(new_n231), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n191), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G902), .ZN(new_n236));
  INV_X1    g050(.A(new_n191), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n224), .A2(new_n231), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n237), .B1(new_n238), .B2(KEYINPUT76), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n235), .A2(new_n236), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT25), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n235), .A2(KEYINPUT25), .A3(new_n236), .A4(new_n239), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G217), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n245), .B1(G234), .B2(new_n236), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(G902), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n235), .A2(new_n239), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(G472), .A2(G902), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT2), .B(G113), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(G116), .B(G119), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G116), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(G119), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n196), .A2(G116), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n252), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G128), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(KEYINPUT1), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n209), .A2(G143), .ZN(new_n263));
  INV_X1    g077(.A(G143), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G146), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n262), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n192), .A2(new_n193), .B1(new_n263), .B2(KEYINPUT1), .ZN(new_n267));
  XNOR2_X1  g081(.A(G143), .B(G146), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G137), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT64), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT64), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G137), .ZN(new_n273));
  INV_X1    g087(.A(G134), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n271), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G131), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n276), .B1(G134), .B2(G137), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT65), .ZN(new_n279));
  AND2_X1   g093(.A1(KEYINPUT11), .A2(G134), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n271), .A2(new_n273), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(KEYINPUT11), .A2(G134), .ZN(new_n282));
  NOR2_X1   g096(.A1(KEYINPUT11), .A2(G134), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n282), .B1(new_n283), .B2(G137), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n281), .A2(new_n276), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT65), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n275), .A2(new_n286), .A3(new_n277), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n269), .A2(new_n279), .A3(new_n285), .A4(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT30), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT0), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n263), .B(new_n265), .C1(new_n290), .C2(new_n261), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n290), .A2(new_n261), .ZN(new_n292));
  NOR2_X1   g106(.A1(KEYINPUT0), .A2(G128), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n291), .B1(new_n294), .B2(new_n268), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n281), .A2(new_n276), .A3(new_n284), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n276), .B1(new_n281), .B2(new_n284), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n288), .A2(new_n289), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n289), .B1(new_n288), .B2(new_n298), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n260), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n260), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n288), .A2(new_n302), .A3(new_n298), .ZN(new_n303));
  XOR2_X1   g117(.A(KEYINPUT67), .B(KEYINPUT27), .Z(new_n304));
  NOR2_X1   g118(.A1(G237), .A2(G953), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G210), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n304), .B(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT26), .B(G101), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n307), .B(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n301), .A2(new_n303), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT68), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n301), .A2(KEYINPUT68), .A3(new_n303), .A4(new_n309), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n312), .A2(KEYINPUT31), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT31), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n301), .A2(new_n315), .A3(new_n303), .A4(new_n309), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n288), .A2(new_n298), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n260), .B1(new_n317), .B2(KEYINPUT70), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT70), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n288), .A2(new_n319), .A3(new_n298), .ZN(new_n320));
  AOI21_X1  g134(.A(KEYINPUT28), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n288), .A2(new_n302), .A3(new_n298), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n302), .B1(new_n288), .B2(new_n298), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT28), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT69), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI211_X1 g140(.A(KEYINPUT69), .B(KEYINPUT28), .C1(new_n322), .C2(new_n323), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n321), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n316), .B1(new_n328), .B2(new_n309), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n251), .B1(new_n314), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT32), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n318), .A2(new_n320), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n317), .A2(new_n260), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n303), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT69), .B1(new_n336), .B2(KEYINPUT28), .ZN(new_n337));
  INV_X1    g151(.A(new_n327), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n334), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n309), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n312), .A2(KEYINPUT31), .A3(new_n313), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n342), .A3(new_n316), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT32), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n344), .A3(new_n251), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n331), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n301), .A2(new_n303), .ZN(new_n347));
  AOI21_X1  g161(.A(KEYINPUT29), .B1(new_n347), .B2(new_n340), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n348), .B1(new_n339), .B2(new_n340), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT71), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n324), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n336), .A2(KEYINPUT71), .A3(KEYINPUT28), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n334), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n309), .A2(KEYINPUT29), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n349), .B(new_n236), .C1(new_n354), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G472), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n250), .B1(new_n346), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(G210), .B1(G237), .B2(G902), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n192), .A2(new_n193), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n263), .A2(KEYINPUT1), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n268), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n266), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n212), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n295), .A2(G125), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G224), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(G953), .ZN(new_n370));
  XOR2_X1   g184(.A(new_n368), .B(new_n370), .Z(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G122), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G110), .ZN(new_n374));
  INV_X1    g188(.A(G110), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G122), .ZN(new_n376));
  AOI21_X1  g190(.A(KEYINPUT85), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n374), .A2(new_n376), .A3(KEYINPUT85), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XOR2_X1   g194(.A(new_n380), .B(KEYINPUT86), .Z(new_n381));
  INV_X1    g195(.A(G104), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT3), .B1(new_n382), .B2(G107), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT3), .ZN(new_n384));
  INV_X1    g198(.A(G107), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(G104), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n382), .A2(G107), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n383), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT4), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n389), .A3(G101), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n260), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT77), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n388), .A2(G101), .ZN(new_n393));
  INV_X1    g207(.A(G101), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n383), .A2(new_n386), .A3(new_n394), .A4(new_n387), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT4), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n392), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n388), .A2(G101), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n398), .A2(KEYINPUT77), .A3(KEYINPUT4), .A4(new_n395), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n391), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n254), .A2(KEYINPUT5), .ZN(new_n401));
  INV_X1    g215(.A(G113), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT5), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n402), .B1(new_n257), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n255), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n382), .A2(G107), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n385), .A2(G104), .ZN(new_n408));
  OAI21_X1  g222(.A(G101), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n395), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT84), .B1(new_n406), .B2(new_n410), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n401), .A2(new_n404), .B1(new_n253), .B2(new_n254), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n395), .A2(new_n409), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT84), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n381), .B1(new_n400), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n380), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n400), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT6), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n417), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  OAI211_X1 g235(.A(KEYINPUT6), .B(new_n381), .C1(new_n400), .C2(new_n416), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n372), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n406), .A2(new_n410), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n412), .A2(new_n413), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n378), .A2(new_n379), .A3(KEYINPUT8), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT8), .ZN(new_n428));
  INV_X1    g242(.A(new_n379), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n428), .B1(new_n429), .B2(new_n377), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n426), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT88), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT7), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n370), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n435), .A2(KEYINPUT87), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n437), .B1(new_n368), .B2(new_n439), .ZN(new_n440));
  AOI211_X1 g254(.A(new_n436), .B(new_n438), .C1(new_n366), .C2(new_n367), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n433), .B(new_n434), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n411), .A2(new_n415), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n397), .A2(new_n399), .ZN(new_n444));
  INV_X1    g258(.A(new_n391), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n443), .A2(new_n446), .A3(new_n380), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n263), .A2(new_n265), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT1), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n450), .B1(G143), .B2(new_n209), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n449), .B1(new_n202), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(G125), .B1(new_n452), .B2(new_n266), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n449), .B1(new_n292), .B2(new_n293), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n212), .B1(new_n454), .B2(new_n291), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n439), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n436), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n368), .A2(new_n437), .A3(new_n439), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n457), .A2(new_n458), .B1(new_n426), .B2(new_n432), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n459), .A2(new_n434), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n236), .B1(new_n448), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n361), .B1(new_n423), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n443), .A2(new_n446), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n447), .A2(KEYINPUT6), .B1(new_n463), .B2(new_n381), .ZN(new_n464));
  INV_X1    g278(.A(new_n422), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n371), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n400), .A2(new_n416), .ZN(new_n467));
  AOI22_X1  g281(.A1(new_n459), .A2(new_n434), .B1(new_n467), .B2(new_n380), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n433), .B1(new_n440), .B2(new_n441), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT88), .ZN(new_n470));
  AOI21_X1  g284(.A(G902), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n466), .A2(new_n471), .A3(new_n360), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT89), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n462), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n466), .A2(new_n471), .A3(KEYINPUT89), .A4(new_n360), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT20), .ZN(new_n477));
  INV_X1    g291(.A(G237), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(new_n187), .A3(G214), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n264), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n305), .A2(G143), .A3(G214), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(KEYINPUT91), .B1(new_n482), .B2(G131), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(G131), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT91), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n480), .A2(new_n485), .A3(new_n276), .A4(new_n481), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n211), .A2(new_n213), .A3(KEYINPUT19), .ZN(new_n488));
  AOI21_X1  g302(.A(KEYINPUT19), .B1(new_n211), .B2(new_n213), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n209), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n487), .A2(new_n226), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(KEYINPUT18), .A2(G131), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n480), .A2(new_n481), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n482), .A2(KEYINPUT18), .A3(G131), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n211), .A2(new_n213), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G146), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n496), .A2(KEYINPUT90), .A3(new_n227), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT90), .B1(new_n496), .B2(new_n227), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n493), .B(new_n494), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n491), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(G113), .B(G122), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(new_n382), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n487), .A2(KEYINPUT17), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT17), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n226), .B(new_n218), .C1(new_n506), .C2(new_n484), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n502), .B(new_n499), .C1(new_n505), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(G475), .A2(G902), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n477), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n510), .ZN(new_n512));
  AOI211_X1 g326(.A(KEYINPUT20), .B(new_n512), .C1(new_n504), .C2(new_n508), .ZN(new_n513));
  INV_X1    g327(.A(G475), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n499), .B1(new_n505), .B2(new_n507), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n503), .ZN(new_n516));
  AOI21_X1  g330(.A(G902), .B1(new_n516), .B2(new_n508), .ZN(new_n517));
  OAI22_X1  g331(.A1(new_n511), .A2(new_n513), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n256), .A2(G122), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n373), .A2(G116), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n519), .A2(new_n520), .A3(G107), .ZN(new_n521));
  AOI21_X1  g335(.A(KEYINPUT14), .B1(new_n373), .B2(G116), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT93), .B1(new_n522), .B2(new_n520), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT93), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n256), .A2(G122), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n524), .B(new_n525), .C1(new_n519), .C2(KEYINPUT14), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT94), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT14), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n520), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT94), .B1(new_n525), .B2(KEYINPUT14), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n523), .A2(new_n526), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n521), .B1(new_n531), .B2(G107), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n192), .A2(G143), .A3(new_n193), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT92), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n192), .A2(KEYINPUT92), .A3(G143), .A4(new_n193), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n261), .A2(G143), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n274), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  AOI211_X1 g354(.A(G134), .B(new_n538), .C1(new_n535), .C2(new_n536), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n532), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n537), .A2(new_n274), .A3(new_n539), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n519), .A2(new_n520), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n544), .B(new_n385), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n538), .B(KEYINPUT13), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n535), .B2(new_n536), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n543), .B(new_n545), .C1(new_n547), .C2(new_n274), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT9), .B(G234), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n549), .A2(new_n245), .A3(G953), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n542), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n550), .B1(new_n542), .B2(new_n548), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n236), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(G478), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n554), .A2(KEYINPUT15), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n553), .B(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n518), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(G952), .ZN(new_n558));
  OR2_X1    g372(.A1(new_n558), .A2(KEYINPUT95), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(KEYINPUT95), .ZN(new_n560));
  AOI21_X1  g374(.A(G953), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(G234), .A2(G237), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(KEYINPUT96), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n562), .A2(G902), .A3(G953), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT21), .B(G898), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n557), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(G214), .B1(G237), .B2(G902), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n476), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(G221), .B1(new_n549), .B2(G902), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT79), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n266), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n449), .B1(new_n451), .B2(new_n261), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n266), .A2(new_n576), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n413), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT10), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n582), .B1(new_n452), .B2(new_n266), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n581), .A2(new_n582), .B1(new_n413), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT78), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n295), .A2(new_n390), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n585), .B1(new_n444), .B2(new_n587), .ZN(new_n588));
  AOI211_X1 g402(.A(KEYINPUT78), .B(new_n586), .C1(new_n397), .C2(new_n399), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n584), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n296), .A2(new_n297), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n591), .B(new_n584), .C1(new_n588), .C2(new_n589), .ZN(new_n595));
  XNOR2_X1  g409(.A(G110), .B(G140), .ZN(new_n596));
  INV_X1    g410(.A(G227), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(G953), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n596), .B(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n594), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT12), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(KEYINPUT81), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT80), .B1(new_n413), .B2(new_n269), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT80), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n410), .A2(new_n606), .A3(new_n266), .A4(new_n452), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n605), .A2(new_n581), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n604), .B1(new_n608), .B2(new_n592), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n603), .A2(KEYINPUT81), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n608), .A2(KEYINPUT81), .A3(new_n603), .A4(new_n592), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n595), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT82), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n610), .ZN(new_n616));
  AOI211_X1 g430(.A(new_n604), .B(new_n616), .C1(new_n608), .C2(new_n592), .ZN(new_n617));
  AND4_X1   g431(.A1(KEYINPUT81), .A2(new_n608), .A3(new_n603), .A4(new_n592), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n619), .A2(KEYINPUT82), .A3(new_n595), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n602), .B1(new_n621), .B2(new_n599), .ZN(new_n622));
  OAI21_X1  g436(.A(G469), .B1(new_n622), .B2(G902), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT83), .B(G469), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n619), .A2(new_n600), .A3(new_n595), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n600), .B1(new_n593), .B2(new_n595), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n236), .B(new_n625), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n575), .B1(new_n623), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n359), .A2(new_n573), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G101), .ZN(G3));
  NAND2_X1  g446(.A1(new_n623), .A2(new_n629), .ZN(new_n633));
  INV_X1    g447(.A(G472), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n343), .B2(new_n236), .ZN(new_n635));
  INV_X1    g449(.A(new_n330), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n250), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n633), .A2(new_n637), .A3(new_n574), .A4(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n572), .B1(new_n462), .B2(new_n472), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n569), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT33), .B1(new_n551), .B2(new_n552), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n542), .A2(new_n548), .ZN(new_n644));
  INV_X1    g458(.A(new_n550), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT33), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n542), .A2(new_n548), .A3(new_n550), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n643), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n554), .A2(G902), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(KEYINPUT97), .B1(new_n553), .B2(new_n554), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n650), .A2(KEYINPUT97), .A3(new_n651), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n518), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n642), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n640), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n659), .B(KEYINPUT98), .Z(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT34), .B(G104), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G6));
  INV_X1    g476(.A(new_n518), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n556), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n642), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n640), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT35), .B(G107), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  NOR2_X1   g482(.A1(new_n237), .A2(KEYINPUT36), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(new_n238), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n248), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n247), .A2(KEYINPUT99), .A3(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT99), .ZN(new_n673));
  INV_X1    g487(.A(new_n246), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n242), .B2(new_n243), .ZN(new_n675));
  INV_X1    g489(.A(new_n671), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n673), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n672), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n630), .A2(new_n573), .A3(new_n637), .A4(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT37), .B(G110), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G12));
  AND3_X1   g495(.A1(new_n672), .A2(new_n641), .A3(new_n677), .ZN(new_n682));
  INV_X1    g496(.A(new_n251), .ZN(new_n683));
  INV_X1    g497(.A(new_n316), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n684), .B1(new_n339), .B2(new_n340), .ZN(new_n685));
  AOI211_X1 g499(.A(KEYINPUT32), .B(new_n683), .C1(new_n685), .C2(new_n342), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n344), .B1(new_n343), .B2(new_n251), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n358), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(G900), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n565), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n564), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n663), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n556), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n630), .A2(new_n682), .A3(new_n688), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G128), .ZN(G30));
  NAND2_X1  g511(.A1(new_n312), .A2(new_n313), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n698), .B1(new_n340), .B2(new_n336), .ZN(new_n699));
  OAI21_X1  g513(.A(G472), .B1(new_n699), .B2(G902), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n346), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT101), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n346), .A2(KEYINPUT101), .A3(new_n700), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n691), .B(new_n706), .Z(new_n707));
  NAND2_X1  g521(.A1(new_n630), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(KEYINPUT40), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n476), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n474), .A2(new_n475), .A3(new_n710), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n675), .A2(new_n676), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n518), .A2(new_n571), .A3(new_n556), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(KEYINPUT102), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT102), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n715), .B2(new_n716), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n714), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT40), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n630), .A2(new_n722), .A3(new_n707), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n705), .A2(new_n709), .A3(new_n721), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G143), .ZN(G45));
  NAND4_X1  g539(.A1(new_n654), .A2(new_n518), .A3(new_n655), .A4(new_n692), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT104), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n630), .A2(new_n728), .A3(new_n682), .A4(new_n688), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G146), .ZN(G48));
  INV_X1    g544(.A(new_n628), .ZN(new_n731));
  AOI21_X1  g545(.A(G902), .B1(new_n731), .B2(new_n626), .ZN(new_n732));
  INV_X1    g546(.A(G469), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n629), .B(new_n574), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n658), .A2(new_n688), .A3(new_n638), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT41), .B(G113), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G15));
  NAND4_X1  g552(.A1(new_n665), .A2(new_n688), .A3(new_n638), .A4(new_n735), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G116), .ZN(G18));
  NOR2_X1   g554(.A1(new_n734), .A2(new_n568), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n682), .A2(new_n741), .A3(new_n557), .A4(new_n688), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G119), .ZN(G21));
  AOI21_X1  g557(.A(new_n684), .B1(new_n354), .B2(new_n340), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n683), .B1(new_n744), .B2(new_n342), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n635), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n462), .A2(new_n472), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n716), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n741), .A2(new_n638), .A3(new_n746), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G122), .ZN(G24));
  INV_X1    g564(.A(new_n641), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n734), .A2(new_n751), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n635), .A2(new_n715), .A3(new_n745), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n728), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(KEYINPUT105), .B(G125), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n754), .B(new_n755), .ZN(G27));
  INV_X1    g570(.A(KEYINPUT107), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT106), .B1(new_n686), .B2(new_n687), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT106), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n331), .A2(new_n759), .A3(new_n345), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n758), .A2(new_n358), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n638), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n572), .B1(new_n474), .B2(new_n475), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n630), .A2(new_n728), .A3(KEYINPUT42), .A4(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n757), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(KEYINPUT82), .B1(new_n619), .B2(new_n595), .ZN(new_n766));
  AND4_X1   g580(.A1(KEYINPUT82), .A2(new_n595), .A3(new_n611), .A4(new_n612), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n599), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n602), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n733), .B1(new_n770), .B2(new_n236), .ZN(new_n771));
  INV_X1    g585(.A(new_n629), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n763), .B(new_n574), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n656), .A2(new_n727), .A3(new_n518), .A4(new_n692), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n726), .A2(KEYINPUT104), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(KEYINPUT42), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n777), .A2(KEYINPUT107), .A3(new_n638), .A4(new_n761), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT42), .ZN(new_n779));
  INV_X1    g593(.A(new_n773), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(new_n359), .A3(new_n728), .ZN(new_n781));
  AOI22_X1  g595(.A1(new_n765), .A2(new_n778), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(new_n276), .ZN(G33));
  NAND3_X1  g597(.A1(new_n780), .A2(new_n359), .A3(new_n695), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G134), .ZN(G36));
  INV_X1    g599(.A(new_n656), .ZN(new_n786));
  OAI21_X1  g600(.A(KEYINPUT43), .B1(new_n786), .B2(new_n518), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT43), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n656), .A2(new_n788), .A3(new_n663), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n790), .A2(new_n637), .A3(new_n715), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n791), .A2(KEYINPUT44), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(KEYINPUT44), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(new_n763), .A3(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT109), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n600), .B1(new_n615), .B2(new_n620), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n796), .B1(new_n797), .B2(new_n602), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n768), .A2(KEYINPUT45), .A3(new_n769), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n799), .A3(G469), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(KEYINPUT108), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT108), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n798), .A2(new_n799), .A3(new_n802), .A4(G469), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n733), .A2(new_n236), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT46), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n795), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n807), .ZN(new_n810));
  AOI211_X1 g624(.A(KEYINPUT109), .B(new_n810), .C1(new_n801), .C2(new_n803), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n805), .B1(new_n801), .B2(new_n803), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n629), .B1(new_n814), .B2(KEYINPUT46), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n574), .B(new_n707), .C1(new_n813), .C2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT110), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n808), .A2(new_n811), .ZN(new_n819));
  INV_X1    g633(.A(new_n815), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n575), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n821), .A2(KEYINPUT110), .A3(new_n707), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n794), .B1(new_n818), .B2(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(new_n270), .ZN(G39));
  INV_X1    g638(.A(new_n728), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n476), .A2(new_n571), .ZN(new_n826));
  NOR4_X1   g640(.A1(new_n825), .A2(new_n688), .A3(new_n826), .A4(new_n638), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n821), .A2(KEYINPUT47), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT47), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n815), .A2(new_n808), .A3(new_n811), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n830), .B1(new_n831), .B2(new_n575), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n828), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(new_n210), .ZN(G42));
  NOR4_X1   g648(.A1(new_n786), .A2(new_n572), .A3(new_n518), .A4(new_n575), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n629), .B1(new_n732), .B2(new_n733), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n836), .A2(KEYINPUT49), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(KEYINPUT49), .B2(new_n836), .ZN(new_n839));
  INV_X1    g653(.A(new_n705), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n839), .A2(new_n840), .A3(new_n638), .A4(new_n714), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n696), .A2(new_n754), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT52), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n747), .A2(new_n715), .A3(new_n716), .A4(new_n692), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n346), .A2(KEYINPUT101), .A3(new_n700), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT101), .B1(new_n346), .B2(new_n700), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n630), .B(new_n845), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n843), .A2(new_n844), .A3(new_n729), .A4(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n729), .A2(new_n696), .A3(new_n754), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n630), .A2(new_n845), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n851), .B1(new_n703), .B2(new_n704), .ZN(new_n852));
  OAI21_X1  g666(.A(KEYINPUT52), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT112), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n849), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n854), .B1(new_n849), .B2(new_n853), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n742), .A2(new_n736), .A3(new_n749), .A4(new_n739), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n631), .A2(new_n679), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n694), .A2(KEYINPUT111), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT111), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n556), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n693), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n678), .A2(new_n688), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n753), .A2(new_n774), .A3(new_n775), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n773), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n476), .A2(new_n572), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n860), .A2(new_n862), .A3(new_n663), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n657), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n867), .A2(new_n869), .A3(new_n569), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n639), .A2(new_n870), .ZN(new_n871));
  NOR4_X1   g685(.A1(new_n858), .A2(new_n859), .A3(new_n866), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n765), .A2(new_n778), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n781), .A2(new_n779), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n872), .A2(new_n875), .A3(new_n784), .ZN(new_n876));
  OAI211_X1 g690(.A(KEYINPUT113), .B(new_n842), .C1(new_n857), .C2(new_n876), .ZN(new_n877));
  AND4_X1   g691(.A1(new_n736), .A2(new_n742), .A3(new_n739), .A4(new_n749), .ZN(new_n878));
  INV_X1    g692(.A(new_n866), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n631), .A2(new_n679), .ZN(new_n880));
  INV_X1    g694(.A(new_n871), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n878), .A2(new_n879), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n784), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n882), .A2(new_n782), .A3(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n884), .A2(KEYINPUT53), .A3(new_n849), .A4(new_n853), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n877), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n884), .B1(new_n856), .B2(new_n855), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT113), .B1(new_n887), .B2(new_n842), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT54), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n849), .A2(new_n853), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n842), .B1(new_n876), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT114), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n884), .B(KEYINPUT53), .C1(new_n856), .C2(new_n855), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT114), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n895), .B(new_n842), .C1(new_n876), .C2(new_n890), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n892), .A2(new_n893), .A3(new_n894), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n889), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g712(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n899));
  OAI21_X1  g713(.A(KEYINPUT116), .B1(new_n790), .B2(new_n564), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT116), .ZN(new_n901));
  INV_X1    g715(.A(new_n564), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n787), .A2(new_n901), .A3(new_n902), .A4(new_n789), .ZN(new_n903));
  AOI211_X1 g717(.A(new_n734), .B(new_n826), .C1(new_n900), .C2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n762), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n899), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n746), .A2(new_n638), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n900), .B2(new_n903), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n752), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n561), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n904), .A2(new_n905), .A3(new_n899), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n826), .A2(new_n564), .A3(new_n734), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n840), .A2(new_n638), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT117), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n840), .A2(KEYINPUT117), .A3(new_n638), .A4(new_n913), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n911), .B(new_n912), .C1(new_n657), .C2(new_n918), .ZN(new_n919));
  AOI211_X1 g733(.A(new_n571), .B(new_n734), .C1(new_n712), .C2(new_n713), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT50), .B1(new_n908), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n908), .A2(KEYINPUT50), .A3(new_n920), .ZN(new_n923));
  AOI22_X1  g737(.A1(new_n922), .A2(new_n923), .B1(new_n753), .B2(new_n904), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n656), .A2(new_n518), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n916), .A2(new_n917), .A3(new_n925), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n924), .A2(KEYINPUT51), .A3(new_n926), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n829), .B(new_n832), .C1(new_n574), .C2(new_n836), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n928), .A2(new_n763), .A3(new_n908), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n919), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n904), .A2(new_n753), .ZN(new_n931));
  INV_X1    g745(.A(new_n923), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n931), .B1(new_n932), .B2(new_n921), .ZN(new_n933));
  INV_X1    g747(.A(new_n926), .ZN(new_n934));
  OAI21_X1  g748(.A(KEYINPUT118), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT118), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n924), .A2(new_n936), .A3(new_n926), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n929), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  XOR2_X1   g752(.A(KEYINPUT115), .B(KEYINPUT51), .Z(new_n939));
  OAI21_X1  g753(.A(new_n930), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n898), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(G952), .A2(G953), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n841), .B1(new_n941), .B2(new_n942), .ZN(G75));
  NAND3_X1  g757(.A1(new_n892), .A2(new_n894), .A3(new_n896), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n944), .A2(G210), .A3(G902), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT56), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n464), .A2(new_n371), .A3(new_n465), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n947), .A2(new_n423), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT55), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n945), .A2(new_n946), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n949), .B1(new_n945), .B2(new_n946), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n187), .A2(G952), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(G51));
  NAND2_X1  g767(.A1(new_n894), .A2(new_n896), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n782), .A2(new_n883), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n955), .A2(new_n872), .A3(new_n849), .A4(new_n853), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n895), .B1(new_n956), .B2(new_n842), .ZN(new_n957));
  OAI21_X1  g771(.A(KEYINPUT54), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n897), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n805), .B(KEYINPUT57), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n627), .A2(new_n628), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n944), .A2(G902), .A3(new_n803), .A4(new_n801), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n952), .B1(new_n964), .B2(new_n965), .ZN(G54));
  NAND2_X1  g780(.A1(KEYINPUT58), .A2(G475), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT120), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n944), .A2(G902), .A3(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n509), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n971), .A2(new_n972), .A3(new_n952), .ZN(G60));
  NAND2_X1  g787(.A1(G478), .A2(G902), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT59), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n650), .B1(new_n898), .B2(new_n975), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n650), .A2(new_n975), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n959), .A2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n952), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n976), .A2(new_n980), .ZN(G63));
  NAND2_X1  g795(.A1(G217), .A2(G902), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT121), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT60), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n954), .B2(new_n957), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n235), .A2(new_n239), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n944), .A2(new_n670), .A3(new_n984), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n987), .A2(new_n979), .A3(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT61), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n987), .A2(KEYINPUT61), .A3(new_n979), .A4(new_n988), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(G66));
  OAI21_X1  g807(.A(G953), .B1(new_n566), .B2(new_n369), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n878), .A2(new_n880), .A3(new_n881), .ZN(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n994), .B1(new_n996), .B2(G953), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n421), .B(new_n422), .C1(G898), .C2(new_n187), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n997), .B(new_n998), .ZN(G69));
  NOR2_X1   g813(.A1(new_n488), .A2(new_n489), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT122), .Z(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(KEYINPUT123), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n299), .A2(new_n300), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1002), .B(new_n1003), .Z(new_n1004));
  INV_X1    g818(.A(new_n850), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n724), .A2(new_n1005), .A3(KEYINPUT62), .ZN(new_n1006));
  AOI21_X1  g820(.A(KEYINPUT62), .B1(new_n724), .B2(new_n1005), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n359), .A2(new_n763), .A3(new_n869), .ZN(new_n1008));
  OAI22_X1  g822(.A1(new_n1006), .A2(new_n1007), .B1(new_n708), .B2(new_n1008), .ZN(new_n1009));
  NOR3_X1   g823(.A1(new_n823), .A2(new_n833), .A3(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1004), .B1(new_n1010), .B2(G953), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n689), .A2(G953), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1012), .B(KEYINPUT124), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT125), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1005), .B1(new_n955), .B2(new_n1015), .ZN(new_n1016));
  NOR3_X1   g830(.A1(new_n782), .A2(KEYINPUT125), .A3(new_n883), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n905), .A2(new_n748), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n794), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(new_n822), .ZN(new_n1021));
  AOI21_X1  g835(.A(KEYINPUT110), .B1(new_n821), .B2(new_n707), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n833), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1018), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1014), .B1(new_n1025), .B2(new_n187), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1011), .B1(new_n1026), .B2(new_n1004), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n597), .A2(new_n689), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n1028), .A2(new_n187), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  OAI221_X1 g844(.A(new_n1011), .B1(new_n187), .B2(new_n1028), .C1(new_n1026), .C2(new_n1004), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1030), .A2(new_n1031), .ZN(G72));
  INV_X1    g846(.A(KEYINPUT113), .ZN(new_n1033));
  INV_X1    g847(.A(new_n856), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n849), .A2(new_n853), .A3(new_n854), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n876), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1033), .B1(new_n1036), .B2(KEYINPUT53), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1037), .A2(new_n885), .A3(new_n877), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n698), .B1(new_n347), .B2(new_n340), .ZN(new_n1039));
  NAND2_X1  g853(.A1(G472), .A2(G902), .ZN(new_n1040));
  XOR2_X1   g854(.A(new_n1040), .B(KEYINPUT63), .Z(new_n1041));
  INV_X1    g855(.A(new_n1041), .ZN(new_n1042));
  NOR2_X1   g856(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1043));
  AND3_X1   g857(.A1(new_n1038), .A2(KEYINPUT127), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g858(.A(KEYINPUT127), .B1(new_n1038), .B2(new_n1043), .ZN(new_n1045));
  NOR2_X1   g859(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g860(.A(KEYINPUT126), .ZN(new_n1047));
  NOR4_X1   g861(.A1(new_n823), .A2(new_n833), .A3(new_n995), .A4(new_n1009), .ZN(new_n1048));
  OAI21_X1  g862(.A(new_n1047), .B1(new_n1048), .B2(new_n1042), .ZN(new_n1049));
  INV_X1    g863(.A(new_n823), .ZN(new_n1050));
  NOR2_X1   g864(.A1(new_n833), .A2(new_n1009), .ZN(new_n1051));
  NAND3_X1  g865(.A1(new_n1050), .A2(new_n1051), .A3(new_n996), .ZN(new_n1052));
  NAND3_X1  g866(.A1(new_n1052), .A2(KEYINPUT126), .A3(new_n1041), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n340), .B1(new_n301), .B2(new_n303), .ZN(new_n1054));
  NAND3_X1  g868(.A1(new_n1049), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  NAND4_X1  g869(.A1(new_n1018), .A2(new_n1023), .A3(new_n1024), .A4(new_n996), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n1056), .A2(new_n1041), .ZN(new_n1057));
  NOR2_X1   g871(.A1(new_n347), .A2(new_n309), .ZN(new_n1058));
  AOI21_X1  g872(.A(new_n952), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g873(.A1(new_n1055), .A2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g874(.A1(new_n1046), .A2(new_n1060), .ZN(G57));
endmodule


