

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594;

  XNOR2_X1 U324 ( .A(n433), .B(n432), .ZN(n434) );
  INV_X1 U325 ( .A(G99GAT), .ZN(n432) );
  XOR2_X1 U326 ( .A(n486), .B(KEYINPUT28), .Z(n540) );
  XNOR2_X1 U327 ( .A(n292), .B(n356), .ZN(n357) );
  XOR2_X1 U328 ( .A(n419), .B(n353), .Z(n292) );
  INV_X1 U329 ( .A(KEYINPUT99), .ZN(n399) );
  XNOR2_X1 U330 ( .A(n480), .B(KEYINPUT64), .ZN(n481) );
  XNOR2_X1 U331 ( .A(n482), .B(n481), .ZN(n535) );
  XNOR2_X1 U332 ( .A(n457), .B(KEYINPUT105), .ZN(n458) );
  NOR2_X1 U333 ( .A1(n524), .A2(n485), .ZN(n578) );
  XNOR2_X1 U334 ( .A(n435), .B(n434), .ZN(n438) );
  XNOR2_X1 U335 ( .A(n459), .B(n458), .ZN(n521) );
  XNOR2_X1 U336 ( .A(n358), .B(n357), .ZN(n363) );
  XNOR2_X1 U337 ( .A(n440), .B(n439), .ZN(n564) );
  XNOR2_X1 U338 ( .A(n461), .B(n460), .ZN(n509) );
  INV_X1 U339 ( .A(KEYINPUT39), .ZN(n465) );
  XNOR2_X1 U340 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U341 ( .A(n465), .B(KEYINPUT104), .ZN(n466) );
  XNOR2_X1 U342 ( .A(n492), .B(n491), .ZN(G1351GAT) );
  XNOR2_X1 U343 ( .A(n467), .B(n466), .ZN(G1328GAT) );
  XOR2_X1 U344 ( .A(G148GAT), .B(G120GAT), .Z(n294) );
  XNOR2_X1 U345 ( .A(G127GAT), .B(G155GAT), .ZN(n293) );
  XNOR2_X1 U346 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U347 ( .A(G162GAT), .B(G85GAT), .Z(n296) );
  XNOR2_X1 U348 ( .A(KEYINPUT75), .B(G134GAT), .ZN(n295) );
  XNOR2_X1 U349 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n298), .B(n297), .ZN(n316) );
  XOR2_X1 U351 ( .A(KEYINPUT92), .B(KEYINPUT4), .Z(n300) );
  XNOR2_X1 U352 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n299) );
  XNOR2_X1 U353 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U354 ( .A(KEYINPUT93), .B(KEYINPUT6), .Z(n302) );
  XNOR2_X1 U355 ( .A(G57GAT), .B(KEYINPUT1), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U357 ( .A(n304), .B(n303), .Z(n314) );
  XOR2_X1 U358 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n306) );
  XNOR2_X1 U359 ( .A(KEYINPUT2), .B(G141GAT), .ZN(n305) );
  XNOR2_X1 U360 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U361 ( .A(KEYINPUT3), .B(n307), .Z(n368) );
  XOR2_X1 U362 ( .A(G113GAT), .B(KEYINPUT80), .Z(n309) );
  XNOR2_X1 U363 ( .A(KEYINPUT79), .B(KEYINPUT0), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n309), .B(n308), .ZN(n385) );
  XOR2_X1 U365 ( .A(n385), .B(KEYINPUT94), .Z(n311) );
  NAND2_X1 U366 ( .A1(G225GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U367 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U368 ( .A(n368), .B(n312), .ZN(n313) );
  XNOR2_X1 U369 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U370 ( .A(n316), .B(n315), .Z(n462) );
  XNOR2_X1 U371 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n317) );
  XNOR2_X1 U372 ( .A(n317), .B(KEYINPUT7), .ZN(n436) );
  XNOR2_X1 U373 ( .A(G1GAT), .B(G8GAT), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n318), .B(KEYINPUT68), .ZN(n445) );
  XNOR2_X1 U375 ( .A(n436), .B(n445), .ZN(n331) );
  XOR2_X1 U376 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n320) );
  NAND2_X1 U377 ( .A1(G229GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U379 ( .A(G197GAT), .B(G141GAT), .Z(n322) );
  XNOR2_X1 U380 ( .A(G15GAT), .B(G113GAT), .ZN(n321) );
  XNOR2_X1 U381 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U382 ( .A(n324), .B(n323), .Z(n329) );
  XOR2_X1 U383 ( .A(G169GAT), .B(G50GAT), .Z(n326) );
  XNOR2_X1 U384 ( .A(G36GAT), .B(G43GAT), .ZN(n325) );
  XNOR2_X1 U385 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U386 ( .A(G22GAT), .B(n327), .ZN(n328) );
  XNOR2_X1 U387 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U388 ( .A(n331), .B(n330), .Z(n541) );
  INV_X1 U389 ( .A(n541), .ZN(n580) );
  XOR2_X1 U390 ( .A(KEYINPUT32), .B(KEYINPUT71), .Z(n333) );
  XOR2_X1 U391 ( .A(G99GAT), .B(G120GAT), .Z(n392) );
  XOR2_X1 U392 ( .A(G64GAT), .B(G176GAT), .Z(n353) );
  XNOR2_X1 U393 ( .A(n392), .B(n353), .ZN(n332) );
  XNOR2_X1 U394 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U395 ( .A(KEYINPUT74), .B(KEYINPUT31), .Z(n335) );
  NAND2_X1 U396 ( .A1(G230GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U397 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U398 ( .A(n337), .B(n336), .Z(n339) );
  XOR2_X1 U399 ( .A(G92GAT), .B(G85GAT), .Z(n426) );
  XNOR2_X1 U400 ( .A(n426), .B(KEYINPUT33), .ZN(n338) );
  XNOR2_X1 U401 ( .A(n339), .B(n338), .ZN(n343) );
  XOR2_X1 U402 ( .A(KEYINPUT69), .B(KEYINPUT72), .Z(n341) );
  XNOR2_X1 U403 ( .A(KEYINPUT73), .B(KEYINPUT70), .ZN(n340) );
  XNOR2_X1 U404 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U405 ( .A(n343), .B(n342), .Z(n348) );
  XOR2_X1 U406 ( .A(KEYINPUT13), .B(G57GAT), .Z(n345) );
  XNOR2_X1 U407 ( .A(G71GAT), .B(G78GAT), .ZN(n344) );
  XNOR2_X1 U408 ( .A(n345), .B(n344), .ZN(n444) );
  XNOR2_X1 U409 ( .A(G106GAT), .B(G148GAT), .ZN(n346) );
  XNOR2_X1 U410 ( .A(n346), .B(G204GAT), .ZN(n364) );
  XNOR2_X1 U411 ( .A(n444), .B(n364), .ZN(n347) );
  XNOR2_X1 U412 ( .A(n348), .B(n347), .ZN(n584) );
  NOR2_X1 U413 ( .A1(n580), .A2(n584), .ZN(n496) );
  XNOR2_X1 U414 ( .A(G29GAT), .B(n462), .ZN(n524) );
  XOR2_X1 U415 ( .A(G197GAT), .B(KEYINPUT21), .Z(n350) );
  XNOR2_X1 U416 ( .A(G218GAT), .B(G211GAT), .ZN(n349) );
  XNOR2_X1 U417 ( .A(n350), .B(n349), .ZN(n375) );
  XOR2_X1 U418 ( .A(n375), .B(G8GAT), .Z(n352) );
  NAND2_X1 U419 ( .A1(G226GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U420 ( .A(n352), .B(n351), .ZN(n358) );
  XOR2_X1 U421 ( .A(KEYINPUT76), .B(G36GAT), .Z(n419) );
  XOR2_X1 U422 ( .A(KEYINPUT95), .B(G204GAT), .Z(n355) );
  INV_X1 U423 ( .A(G190GAT), .ZN(n489) );
  XNOR2_X1 U424 ( .A(G190GAT), .B(G92GAT), .ZN(n354) );
  XNOR2_X1 U425 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U426 ( .A(G169GAT), .B(KEYINPUT17), .Z(n360) );
  XNOR2_X1 U427 ( .A(G183GAT), .B(KEYINPUT18), .ZN(n359) );
  XNOR2_X1 U428 ( .A(n360), .B(n359), .ZN(n362) );
  XOR2_X1 U429 ( .A(KEYINPUT83), .B(KEYINPUT19), .Z(n361) );
  XNOR2_X1 U430 ( .A(n362), .B(n361), .ZN(n395) );
  XNOR2_X1 U431 ( .A(n363), .B(n395), .ZN(n526) );
  XNOR2_X1 U432 ( .A(n526), .B(KEYINPUT27), .ZN(n408) );
  NAND2_X1 U433 ( .A1(n524), .A2(n408), .ZN(n534) );
  XOR2_X1 U434 ( .A(G162GAT), .B(G50GAT), .Z(n430) );
  XOR2_X1 U435 ( .A(n430), .B(n364), .Z(n366) );
  NAND2_X1 U436 ( .A1(G228GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U437 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U438 ( .A(n368), .B(n367), .ZN(n379) );
  XOR2_X1 U439 ( .A(KEYINPUT23), .B(KEYINPUT89), .Z(n370) );
  XNOR2_X1 U440 ( .A(KEYINPUT24), .B(KEYINPUT86), .ZN(n369) );
  XNOR2_X1 U441 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U442 ( .A(n371), .B(KEYINPUT90), .Z(n373) );
  XOR2_X1 U443 ( .A(G155GAT), .B(G22GAT), .Z(n452) );
  XNOR2_X1 U444 ( .A(n452), .B(G78GAT), .ZN(n372) );
  XNOR2_X1 U445 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U446 ( .A(n374), .B(KEYINPUT22), .Z(n377) );
  XNOR2_X1 U447 ( .A(n375), .B(KEYINPUT91), .ZN(n376) );
  XNOR2_X1 U448 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U449 ( .A(n379), .B(n378), .ZN(n404) );
  INV_X1 U450 ( .A(n404), .ZN(n486) );
  NOR2_X1 U451 ( .A1(n534), .A2(n540), .ZN(n380) );
  XOR2_X1 U452 ( .A(KEYINPUT96), .B(n380), .Z(n398) );
  XOR2_X1 U453 ( .A(KEYINPUT81), .B(KEYINPUT84), .Z(n382) );
  NAND2_X1 U454 ( .A1(G227GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U455 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U456 ( .A(n383), .B(KEYINPUT65), .Z(n387) );
  XNOR2_X1 U457 ( .A(G43GAT), .B(G190GAT), .ZN(n384) );
  XNOR2_X1 U458 ( .A(n384), .B(G134GAT), .ZN(n420) );
  XNOR2_X1 U459 ( .A(n420), .B(n385), .ZN(n386) );
  XNOR2_X1 U460 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U461 ( .A(G176GAT), .B(KEYINPUT82), .Z(n389) );
  XNOR2_X1 U462 ( .A(G71GAT), .B(KEYINPUT20), .ZN(n388) );
  XNOR2_X1 U463 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U464 ( .A(n391), .B(n390), .Z(n394) );
  XOR2_X1 U465 ( .A(G127GAT), .B(G15GAT), .Z(n453) );
  XNOR2_X1 U466 ( .A(n453), .B(n392), .ZN(n393) );
  XNOR2_X1 U467 ( .A(n394), .B(n393), .ZN(n396) );
  XOR2_X1 U468 ( .A(n396), .B(n395), .Z(n403) );
  INV_X1 U469 ( .A(n403), .ZN(n538) );
  XNOR2_X1 U470 ( .A(n403), .B(KEYINPUT85), .ZN(n397) );
  NOR2_X1 U471 ( .A1(n398), .A2(n397), .ZN(n414) );
  NAND2_X1 U472 ( .A1(n538), .A2(n526), .ZN(n400) );
  XNOR2_X1 U473 ( .A(n400), .B(n399), .ZN(n401) );
  NAND2_X1 U474 ( .A1(n401), .A2(n486), .ZN(n402) );
  XNOR2_X1 U475 ( .A(n402), .B(KEYINPUT25), .ZN(n410) );
  XOR2_X1 U476 ( .A(KEYINPUT98), .B(KEYINPUT26), .Z(n406) );
  NAND2_X1 U477 ( .A1(n404), .A2(n403), .ZN(n405) );
  XNOR2_X1 U478 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U479 ( .A(KEYINPUT97), .B(n407), .Z(n579) );
  AND2_X1 U480 ( .A1(n579), .A2(n408), .ZN(n409) );
  NOR2_X1 U481 ( .A1(n410), .A2(n409), .ZN(n411) );
  NOR2_X1 U482 ( .A1(n411), .A2(n524), .ZN(n412) );
  XNOR2_X1 U483 ( .A(n412), .B(KEYINPUT100), .ZN(n413) );
  NOR2_X1 U484 ( .A1(n414), .A2(n413), .ZN(n415) );
  XNOR2_X1 U485 ( .A(n415), .B(KEYINPUT101), .ZN(n495) );
  XOR2_X1 U486 ( .A(KEYINPUT75), .B(KEYINPUT11), .Z(n417) );
  XNOR2_X1 U487 ( .A(KEYINPUT66), .B(KEYINPUT10), .ZN(n416) );
  XNOR2_X1 U488 ( .A(n417), .B(n416), .ZN(n440) );
  INV_X1 U489 ( .A(n420), .ZN(n418) );
  NAND2_X1 U490 ( .A1(n418), .A2(n419), .ZN(n423) );
  INV_X1 U491 ( .A(n419), .ZN(n421) );
  NAND2_X1 U492 ( .A1(n421), .A2(n420), .ZN(n422) );
  NAND2_X1 U493 ( .A1(n423), .A2(n422), .ZN(n425) );
  NAND2_X1 U494 ( .A1(G232GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U495 ( .A(n425), .B(n424), .ZN(n427) );
  XNOR2_X1 U496 ( .A(n427), .B(n426), .ZN(n435) );
  XOR2_X1 U497 ( .A(KEYINPUT9), .B(KEYINPUT77), .Z(n429) );
  XNOR2_X1 U498 ( .A(G218GAT), .B(KEYINPUT67), .ZN(n428) );
  XNOR2_X1 U499 ( .A(n429), .B(n428), .ZN(n431) );
  XOR2_X1 U500 ( .A(n431), .B(n430), .Z(n433) );
  XNOR2_X1 U501 ( .A(n436), .B(G106GAT), .ZN(n437) );
  XNOR2_X1 U502 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U503 ( .A(KEYINPUT36), .B(n564), .ZN(n592) );
  XOR2_X1 U504 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n442) );
  NAND2_X1 U505 ( .A1(G231GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U506 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U507 ( .A(n443), .B(KEYINPUT78), .Z(n447) );
  XNOR2_X1 U508 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U509 ( .A(n447), .B(n446), .ZN(n451) );
  XOR2_X1 U510 ( .A(KEYINPUT15), .B(G64GAT), .Z(n449) );
  XNOR2_X1 U511 ( .A(G183GAT), .B(G211GAT), .ZN(n448) );
  XNOR2_X1 U512 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U513 ( .A(n451), .B(n450), .Z(n455) );
  XNOR2_X1 U514 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U515 ( .A(n455), .B(n454), .Z(n561) );
  INV_X1 U516 ( .A(n561), .ZN(n587) );
  NOR2_X1 U517 ( .A1(n592), .A2(n587), .ZN(n456) );
  NAND2_X1 U518 ( .A1(n495), .A2(n456), .ZN(n459) );
  INV_X1 U519 ( .A(KEYINPUT37), .ZN(n457) );
  NAND2_X1 U520 ( .A1(n496), .A2(n521), .ZN(n461) );
  INV_X1 U521 ( .A(KEYINPUT38), .ZN(n460) );
  AND2_X1 U522 ( .A1(n462), .A2(n509), .ZN(n464) );
  NOR2_X1 U523 ( .A1(G29GAT), .A2(n509), .ZN(n463) );
  NOR2_X1 U524 ( .A1(n464), .A2(n463), .ZN(n467) );
  NOR2_X1 U525 ( .A1(n592), .A2(n561), .ZN(n468) );
  XOR2_X1 U526 ( .A(n468), .B(KEYINPUT45), .Z(n469) );
  NOR2_X1 U527 ( .A1(n584), .A2(n469), .ZN(n470) );
  XOR2_X1 U528 ( .A(KEYINPUT115), .B(n470), .Z(n471) );
  NAND2_X1 U529 ( .A1(n471), .A2(n580), .ZN(n479) );
  XOR2_X1 U530 ( .A(n561), .B(KEYINPUT112), .Z(n576) );
  XNOR2_X1 U531 ( .A(n584), .B(KEYINPUT41), .ZN(n555) );
  NOR2_X1 U532 ( .A1(n580), .A2(n555), .ZN(n473) );
  XNOR2_X1 U533 ( .A(KEYINPUT114), .B(KEYINPUT113), .ZN(n472) );
  XNOR2_X1 U534 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n474), .B(KEYINPUT46), .ZN(n475) );
  NAND2_X1 U536 ( .A1(n475), .A2(n564), .ZN(n476) );
  NOR2_X1 U537 ( .A1(n576), .A2(n476), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n477), .B(KEYINPUT47), .ZN(n478) );
  NAND2_X1 U539 ( .A1(n479), .A2(n478), .ZN(n482) );
  XNOR2_X1 U540 ( .A(KEYINPUT116), .B(KEYINPUT48), .ZN(n480) );
  NAND2_X1 U541 ( .A1(n535), .A2(n526), .ZN(n484) );
  XOR2_X1 U542 ( .A(KEYINPUT123), .B(KEYINPUT54), .Z(n483) );
  XNOR2_X1 U543 ( .A(n484), .B(n483), .ZN(n485) );
  NAND2_X1 U544 ( .A1(n578), .A2(n486), .ZN(n487) );
  XNOR2_X1 U545 ( .A(n487), .B(KEYINPUT55), .ZN(n488) );
  NAND2_X1 U546 ( .A1(n488), .A2(n538), .ZN(n574) );
  NOR2_X1 U547 ( .A1(n574), .A2(n564), .ZN(n492) );
  XNOR2_X1 U548 ( .A(KEYINPUT126), .B(KEYINPUT58), .ZN(n490) );
  XNOR2_X1 U549 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n499) );
  NAND2_X1 U550 ( .A1(n587), .A2(n564), .ZN(n493) );
  XOR2_X1 U551 ( .A(KEYINPUT16), .B(n493), .Z(n494) );
  AND2_X1 U552 ( .A1(n495), .A2(n494), .ZN(n511) );
  NAND2_X1 U553 ( .A1(n496), .A2(n511), .ZN(n497) );
  XOR2_X1 U554 ( .A(KEYINPUT102), .B(n497), .Z(n503) );
  NAND2_X1 U555 ( .A1(n524), .A2(n503), .ZN(n498) );
  XNOR2_X1 U556 ( .A(n499), .B(n498), .ZN(G1324GAT) );
  NAND2_X1 U557 ( .A1(n503), .A2(n526), .ZN(n500) );
  XNOR2_X1 U558 ( .A(n500), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U559 ( .A(G15GAT), .B(KEYINPUT35), .Z(n502) );
  NAND2_X1 U560 ( .A1(n538), .A2(n503), .ZN(n501) );
  XNOR2_X1 U561 ( .A(n502), .B(n501), .ZN(G1326GAT) );
  XOR2_X1 U562 ( .A(G22GAT), .B(KEYINPUT103), .Z(n505) );
  NAND2_X1 U563 ( .A1(n503), .A2(n540), .ZN(n504) );
  XNOR2_X1 U564 ( .A(n505), .B(n504), .ZN(G1327GAT) );
  NAND2_X1 U565 ( .A1(n509), .A2(n526), .ZN(n506) );
  XNOR2_X1 U566 ( .A(n506), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U567 ( .A1(n509), .A2(n538), .ZN(n507) );
  XNOR2_X1 U568 ( .A(n507), .B(KEYINPUT40), .ZN(n508) );
  XNOR2_X1 U569 ( .A(G43GAT), .B(n508), .ZN(G1330GAT) );
  NAND2_X1 U570 ( .A1(n509), .A2(n540), .ZN(n510) );
  XNOR2_X1 U571 ( .A(n510), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT107), .B(n555), .Z(n568) );
  NOR2_X1 U573 ( .A1(n541), .A2(n568), .ZN(n522) );
  AND2_X1 U574 ( .A1(n522), .A2(n511), .ZN(n517) );
  NAND2_X1 U575 ( .A1(n517), .A2(n524), .ZN(n514) );
  XNOR2_X1 U576 ( .A(G57GAT), .B(KEYINPUT106), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(KEYINPUT42), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n514), .B(n513), .ZN(G1332GAT) );
  NAND2_X1 U579 ( .A1(n517), .A2(n526), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n515), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U581 ( .A1(n517), .A2(n538), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n516), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n519) );
  NAND2_X1 U584 ( .A1(n517), .A2(n540), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U586 ( .A(G78GAT), .B(n520), .ZN(G1335GAT) );
  NAND2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n523), .B(KEYINPUT109), .ZN(n531) );
  NAND2_X1 U589 ( .A1(n531), .A2(n524), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n525), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U591 ( .A1(n531), .A2(n526), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n527), .B(KEYINPUT110), .ZN(n528) );
  XNOR2_X1 U593 ( .A(G92GAT), .B(n528), .ZN(G1337GAT) );
  XOR2_X1 U594 ( .A(G99GAT), .B(KEYINPUT111), .Z(n530) );
  NAND2_X1 U595 ( .A1(n531), .A2(n538), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n530), .B(n529), .ZN(G1338GAT) );
  NAND2_X1 U597 ( .A1(n540), .A2(n531), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n532), .B(KEYINPUT44), .ZN(n533) );
  XNOR2_X1 U599 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  INV_X1 U600 ( .A(n534), .ZN(n536) );
  NAND2_X1 U601 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U602 ( .A(KEYINPUT117), .B(n537), .ZN(n553) );
  NAND2_X1 U603 ( .A1(n538), .A2(n553), .ZN(n539) );
  NOR2_X1 U604 ( .A1(n540), .A2(n539), .ZN(n546) );
  NAND2_X1 U605 ( .A1(n546), .A2(n541), .ZN(n542) );
  XNOR2_X1 U606 ( .A(KEYINPUT118), .B(n542), .ZN(n543) );
  XNOR2_X1 U607 ( .A(G113GAT), .B(n543), .ZN(G1340GAT) );
  INV_X1 U608 ( .A(n546), .ZN(n550) );
  NOR2_X1 U609 ( .A1(n568), .A2(n550), .ZN(n545) );
  XNOR2_X1 U610 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n548) );
  NAND2_X1 U613 ( .A1(n546), .A2(n576), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U615 ( .A(G127GAT), .B(n549), .ZN(G1342GAT) );
  NOR2_X1 U616 ( .A1(n564), .A2(n550), .ZN(n552) );
  XNOR2_X1 U617 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1343GAT) );
  NAND2_X1 U619 ( .A1(n579), .A2(n553), .ZN(n563) );
  NOR2_X1 U620 ( .A1(n580), .A2(n563), .ZN(n554) );
  XOR2_X1 U621 ( .A(G141GAT), .B(n554), .Z(G1344GAT) );
  NOR2_X1 U622 ( .A1(n555), .A2(n563), .ZN(n560) );
  XOR2_X1 U623 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n557) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U626 ( .A(KEYINPUT52), .B(n558), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1345GAT) );
  NOR2_X1 U628 ( .A1(n561), .A2(n563), .ZN(n562) );
  XOR2_X1 U629 ( .A(G155GAT), .B(n562), .Z(G1346GAT) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U631 ( .A(KEYINPUT122), .B(n565), .Z(n566) );
  XNOR2_X1 U632 ( .A(G162GAT), .B(n566), .ZN(G1347GAT) );
  NOR2_X1 U633 ( .A1(n580), .A2(n574), .ZN(n567) );
  XOR2_X1 U634 ( .A(G169GAT), .B(n567), .Z(G1348GAT) );
  NOR2_X1 U635 ( .A1(n574), .A2(n568), .ZN(n573) );
  XOR2_X1 U636 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n570) );
  XNOR2_X1 U637 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n569) );
  XNOR2_X1 U638 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U639 ( .A(KEYINPUT124), .B(n571), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n573), .B(n572), .ZN(G1349GAT) );
  INV_X1 U641 ( .A(n574), .ZN(n575) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n577), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n591) );
  NOR2_X1 U645 ( .A1(n580), .A2(n591), .ZN(n582) );
  XNOR2_X1 U646 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(G197GAT), .B(n583), .ZN(G1352GAT) );
  XOR2_X1 U649 ( .A(G204GAT), .B(KEYINPUT61), .Z(n586) );
  INV_X1 U650 ( .A(n591), .ZN(n588) );
  NAND2_X1 U651 ( .A1(n588), .A2(n584), .ZN(n585) );
  XNOR2_X1 U652 ( .A(n586), .B(n585), .ZN(G1353GAT) );
  XOR2_X1 U653 ( .A(G211GAT), .B(KEYINPUT127), .Z(n590) );
  NAND2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U655 ( .A(n590), .B(n589), .ZN(G1354GAT) );
  NOR2_X1 U656 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U657 ( .A(KEYINPUT62), .B(n593), .Z(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

