//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 1 1 1 0 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n775, new_n777, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n859, new_n860, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G169gat), .B(G197gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(KEYINPUT90), .B(KEYINPUT12), .Z(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n206), .B(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G229gat), .A2(G233gat), .ZN(new_n210));
  XOR2_X1   g009(.A(new_n210), .B(KEYINPUT13), .Z(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G50gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G43gat), .ZN(new_n214));
  INV_X1    g013(.A(G43gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G50gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n216), .A3(KEYINPUT15), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT92), .ZN(new_n218));
  AND3_X1   g017(.A1(new_n214), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT15), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(new_n216), .B2(new_n218), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G29gat), .ZN(new_n223));
  INV_X1    g022(.A(G36gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT91), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT91), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(G29gat), .B2(G36gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n227), .A3(KEYINPUT14), .ZN(new_n228));
  NAND2_X1  g027(.A1(G29gat), .A2(G36gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT14), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n226), .B(new_n230), .C1(G29gat), .C2(G36gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n228), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n217), .B1(new_n222), .B2(new_n232), .ZN(new_n233));
  AND3_X1   g032(.A1(new_n225), .A2(new_n227), .A3(KEYINPUT14), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n231), .A2(new_n229), .ZN(new_n235));
  OR3_X1    g034(.A1(new_n234), .A2(new_n217), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G15gat), .B(G22gat), .ZN(new_n238));
  INV_X1    g037(.A(G1gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT16), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(G8gat), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n241), .B(new_n242), .C1(G1gat), .C2(new_n238), .ZN(new_n243));
  INV_X1    g042(.A(G15gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G22gat), .ZN(new_n245));
  INV_X1    g044(.A(G22gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G15gat), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n240), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(G1gat), .B1(new_n245), .B2(new_n247), .ZN(new_n249));
  OAI21_X1  g048(.A(G8gat), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n243), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n252), .ZN(new_n253));
  NOR3_X1   g052(.A1(new_n234), .A2(new_n217), .A3(new_n235), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n231), .A2(new_n229), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n255), .B(new_n228), .C1(new_n219), .C2(new_n221), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n254), .B1(new_n217), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(new_n251), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n212), .B1(new_n253), .B2(new_n258), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n233), .A2(new_n251), .A3(new_n236), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT17), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n251), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n261), .B1(new_n233), .B2(new_n236), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n260), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT18), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n266), .B1(G229gat), .B2(G233gat), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n259), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n233), .A2(new_n261), .A3(new_n236), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(new_n252), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n210), .B(new_n258), .C1(new_n270), .C2(new_n263), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(new_n266), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n209), .B1(new_n268), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n259), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n258), .B(new_n267), .C1(new_n270), .C2(new_n263), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n272), .A2(new_n274), .A3(new_n275), .A4(new_n209), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT93), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n268), .A2(KEYINPUT93), .A3(new_n272), .A4(new_n209), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n273), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT87), .ZN(new_n281));
  XNOR2_X1  g080(.A(G113gat), .B(G120gat), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT66), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G113gat), .ZN(new_n285));
  NOR3_X1   g084(.A1(new_n283), .A2(new_n285), .A3(G120gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT67), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G127gat), .B(G134gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT1), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n284), .A2(KEYINPUT67), .A3(new_n287), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT65), .ZN(new_n296));
  INV_X1    g095(.A(G127gat), .ZN(new_n297));
  NOR3_X1   g096(.A1(new_n296), .A2(new_n297), .A3(G134gat), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n298), .B1(new_n296), .B2(new_n289), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n282), .A2(KEYINPUT1), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G155gat), .B(G162gat), .ZN(new_n303));
  XOR2_X1   g102(.A(G141gat), .B(G148gat), .Z(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT74), .B(KEYINPUT2), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G155gat), .ZN(new_n307));
  INV_X1    g106(.A(G162gat), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT2), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n304), .A2(new_n303), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT75), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n304), .A2(KEYINPUT75), .A3(new_n303), .A4(new_n309), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n306), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n316));
  NOR3_X1   g115(.A1(new_n302), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT4), .ZN(new_n318));
  NOR3_X1   g117(.A1(new_n293), .A2(new_n288), .A3(new_n291), .ZN(new_n319));
  INV_X1    g118(.A(new_n301), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n314), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n317), .B1(new_n318), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G225gat), .A2(G233gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT76), .B1(new_n319), .B2(new_n320), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT76), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n286), .B1(new_n283), .B2(new_n282), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n290), .B(new_n289), .C1(new_n328), .C2(KEYINPUT67), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n327), .B(new_n301), .C1(new_n329), .C2(new_n293), .ZN(new_n330));
  AND2_X1   g129(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT3), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n314), .A2(new_n332), .ZN(new_n333));
  AOI211_X1 g132(.A(KEYINPUT3), .B(new_n306), .C1(new_n312), .C2(new_n313), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n325), .B1(new_n331), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT5), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n323), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n326), .A2(KEYINPUT78), .A3(new_n315), .A4(new_n330), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n339), .A2(new_n322), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n326), .A2(new_n315), .A3(new_n330), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT78), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n324), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n315), .A2(KEYINPUT3), .ZN(new_n345));
  INV_X1    g144(.A(new_n334), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n326), .A2(new_n345), .A3(new_n346), .A4(new_n330), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n324), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n316), .B1(new_n302), .B2(new_n315), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n321), .A2(KEYINPUT4), .A3(new_n314), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT5), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n338), .B1(new_n344), .B2(new_n352), .ZN(new_n353));
  XOR2_X1   g152(.A(G1gat), .B(G29gat), .Z(new_n354));
  XNOR2_X1  g153(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G57gat), .B(G85gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n353), .A2(KEYINPUT6), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n353), .A2(KEYINPUT86), .ZN(new_n361));
  AND2_X1   g160(.A1(new_n341), .A2(new_n342), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n339), .A2(new_n322), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n325), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n351), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n336), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n364), .A2(KEYINPUT5), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT86), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n367), .A2(new_n368), .A3(new_n338), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n361), .A2(new_n369), .A3(new_n359), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n358), .B(new_n338), .C1(new_n344), .C2(new_n352), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT6), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n360), .B1(new_n370), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G211gat), .B(G218gat), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  OR2_X1    g176(.A1(KEYINPUT70), .A2(G218gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(KEYINPUT70), .A2(G218gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT22), .B1(new_n380), .B2(G211gat), .ZN(new_n381));
  XOR2_X1   g180(.A(G197gat), .B(G204gat), .Z(new_n382));
  OAI21_X1  g181(.A(new_n377), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n382), .ZN(new_n384));
  INV_X1    g183(.A(G211gat), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n385), .B1(new_n378), .B2(new_n379), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n384), .B(new_n376), .C1(new_n386), .C2(KEYINPUT22), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(G226gat), .A2(G233gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(KEYINPUT72), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT27), .B(G183gat), .ZN(new_n391));
  INV_X1    g190(.A(G190gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT28), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n391), .A2(KEYINPUT28), .A3(new_n392), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G183gat), .A2(G190gat), .ZN(new_n398));
  NOR2_X1   g197(.A1(G169gat), .A2(G176gat), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT26), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n398), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n402), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n399), .A2(KEYINPUT23), .ZN(new_n405));
  NAND2_X1  g204(.A1(G169gat), .A2(G176gat), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT23), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n407), .B1(G169gat), .B2(G176gat), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n405), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  AND2_X1   g208(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT64), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n411), .A3(G190gat), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n398), .ZN(new_n414));
  NAND3_X1  g213(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT64), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n412), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n409), .A2(new_n417), .A3(KEYINPUT25), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT25), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n405), .A2(new_n406), .A3(new_n408), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n398), .A2(new_n413), .B1(new_n410), .B2(G190gat), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n397), .A2(new_n404), .B1(new_n418), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n390), .B1(new_n423), .B2(KEYINPUT29), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT73), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n397), .A2(new_n404), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n418), .A2(new_n422), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n390), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(new_n427), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT29), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n428), .B1(new_n431), .B2(new_n390), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n388), .B(new_n425), .C1(new_n432), .C2(KEYINPUT73), .ZN(new_n433));
  INV_X1    g232(.A(new_n428), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n424), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n383), .A2(new_n387), .A3(KEYINPUT71), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT71), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n388), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n435), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n433), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G8gat), .B(G36gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(G64gat), .B(G92gat), .ZN(new_n442));
  XOR2_X1   g241(.A(new_n441), .B(new_n442), .Z(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n433), .A2(new_n439), .A3(new_n443), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(KEYINPUT30), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n440), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT30), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n449), .A3(new_n443), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT83), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n447), .A2(KEYINPUT83), .A3(new_n450), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n281), .B1(new_n375), .B2(new_n455), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n447), .A2(KEYINPUT83), .A3(new_n450), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT83), .B1(new_n447), .B2(new_n450), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n358), .B1(new_n353), .B2(KEYINPUT86), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n373), .B1(new_n460), .B2(new_n369), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n459), .B(KEYINPUT87), .C1(new_n360), .C2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT35), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(G228gat), .ZN(new_n466));
  INV_X1    g265(.A(G233gat), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n388), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n469), .B1(new_n334), .B2(KEYINPUT29), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT29), .B1(new_n383), .B2(new_n387), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n315), .B1(KEYINPUT3), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n468), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT82), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n473), .B(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n438), .A2(new_n436), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT29), .B1(new_n314), .B2(new_n332), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n472), .B(new_n468), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n475), .A2(new_n246), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n470), .A2(new_n472), .ZN(new_n480));
  INV_X1    g279(.A(new_n468), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n474), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI211_X1 g281(.A(KEYINPUT82), .B(new_n468), .C1(new_n470), .C2(new_n472), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n478), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(G22gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(G78gat), .B(G106gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(new_n213), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n479), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n488), .B1(new_n479), .B2(new_n485), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n465), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n246), .B1(new_n475), .B2(new_n478), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n484), .A2(G22gat), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n487), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n479), .A2(new_n485), .A3(new_n488), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(new_n464), .A3(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G15gat), .B(G43gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(KEYINPUT68), .ZN(new_n498));
  XNOR2_X1  g297(.A(G71gat), .B(G99gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n498), .B(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n302), .B(new_n429), .ZN(new_n501));
  NAND2_X1  g300(.A1(G227gat), .A2(G233gat), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT33), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n500), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(KEYINPUT32), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT69), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n509), .B1(new_n501), .B2(new_n503), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n510), .A2(KEYINPUT34), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(KEYINPUT34), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n504), .B(KEYINPUT32), .C1(new_n505), .C2(new_n500), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n508), .A2(new_n511), .A3(new_n512), .A4(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n508), .A2(new_n513), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n510), .B(KEYINPUT34), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n491), .A2(new_n496), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n456), .A2(new_n462), .A3(new_n463), .A4(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT80), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n358), .B1(new_n367), .B2(new_n338), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n520), .B1(new_n373), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n360), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n353), .A2(new_n359), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n524), .A2(KEYINPUT80), .A3(new_n372), .A4(new_n371), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n522), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(new_n451), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n517), .A2(new_n514), .ZN(new_n528));
  NOR3_X1   g327(.A1(new_n489), .A2(new_n490), .A3(new_n465), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n464), .B1(new_n494), .B2(new_n495), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT35), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n519), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT85), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n343), .A2(new_n324), .A3(new_n322), .A4(new_n339), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n535), .A2(KEYINPUT84), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT39), .B1(new_n535), .B2(KEYINPUT84), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n535), .A2(KEYINPUT84), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT84), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n340), .A2(new_n540), .A3(new_n324), .A4(new_n343), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n539), .A2(new_n541), .A3(KEYINPUT85), .A4(KEYINPUT39), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n323), .A2(new_n347), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(new_n325), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n538), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(KEYINPUT39), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n546), .A2(new_n359), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT40), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n545), .A2(KEYINPUT40), .A3(new_n547), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n550), .A2(new_n551), .A3(new_n455), .A4(new_n370), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT38), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n444), .B1(new_n440), .B2(KEYINPUT37), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n440), .A2(KEYINPUT37), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n553), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n425), .B1(new_n432), .B2(KEYINPUT73), .ZN(new_n558));
  AOI22_X1  g357(.A1(new_n558), .A2(new_n469), .B1(new_n432), .B2(new_n476), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT37), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n553), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n446), .B1(new_n561), .B2(new_n554), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  AOI22_X1  g362(.A1(new_n375), .A2(new_n563), .B1(new_n491), .B2(new_n496), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n552), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT36), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n528), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n517), .A2(new_n514), .A3(KEYINPUT36), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n529), .A2(new_n530), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n569), .B1(new_n527), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n533), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT88), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n533), .A2(new_n572), .A3(KEYINPUT88), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n280), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G85gat), .A2(G92gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT7), .ZN(new_n579));
  XNOR2_X1  g378(.A(G99gat), .B(G106gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(G99gat), .A2(G106gat), .ZN(new_n581));
  INV_X1    g380(.A(G85gat), .ZN(new_n582));
  INV_X1    g381(.A(G92gat), .ZN(new_n583));
  AOI22_X1  g382(.A1(KEYINPUT8), .A2(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n579), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n580), .B1(new_n579), .B2(new_n584), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AND2_X1   g386(.A1(G232gat), .A2(G233gat), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n257), .A2(new_n587), .B1(KEYINPUT41), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n587), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n269), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n589), .B1(new_n591), .B2(new_n263), .ZN(new_n592));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n588), .A2(KEYINPUT41), .ZN(new_n595));
  XNOR2_X1  g394(.A(G134gat), .B(G162gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n594), .B(new_n597), .Z(new_n598));
  INV_X1    g397(.A(G57gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(G64gat), .ZN(new_n600));
  INV_X1    g399(.A(G64gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(G57gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G71gat), .A2(G78gat), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT9), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n604), .ZN(new_n607));
  NOR2_X1   g406(.A1(G71gat), .A2(G78gat), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n603), .B(new_n606), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n580), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT97), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n603), .A2(new_n606), .ZN(new_n612));
  INV_X1    g411(.A(G71gat), .ZN(new_n613));
  INV_X1    g412(.A(G78gat), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n613), .A2(new_n614), .A3(KEYINPUT94), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT94), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n616), .B1(G71gat), .B2(G78gat), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n607), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT95), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n612), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n619), .B1(new_n612), .B2(new_n618), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n609), .B(new_n611), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(new_n590), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n612), .A2(new_n618), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT95), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(new_n620), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n627), .A2(new_n587), .A3(new_n609), .A4(new_n611), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT10), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n624), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n627), .A2(new_n609), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n631), .A2(KEYINPUT10), .A3(new_n587), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G230gat), .A2(G233gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G120gat), .B(G148gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT98), .ZN(new_n637));
  XNOR2_X1  g436(.A(G176gat), .B(G204gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  AND2_X1   g438(.A1(new_n624), .A2(new_n628), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n635), .B(new_n639), .C1(new_n640), .C2(new_n634), .ZN(new_n641));
  INV_X1    g440(.A(new_n639), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n640), .A2(new_n634), .ZN(new_n643));
  INV_X1    g442(.A(new_n634), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n644), .B1(new_n630), .B2(new_n632), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n642), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n631), .A2(KEYINPUT21), .ZN(new_n648));
  NAND2_X1  g447(.A1(G231gat), .A2(G233gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G127gat), .B(G155gat), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n651), .B(KEYINPUT96), .Z(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n649), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n648), .B(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n652), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(G183gat), .B(G211gat), .Z(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n659), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n653), .A2(new_n657), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n631), .A2(KEYINPUT21), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n252), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n660), .A2(new_n667), .A3(new_n662), .ZN(new_n670));
  AOI211_X1 g469(.A(new_n598), .B(new_n647), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT99), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n577), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(new_n526), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(new_n239), .ZN(G1324gat));
  NOR2_X1   g476(.A1(new_n675), .A2(new_n459), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT16), .B(G8gat), .Z(new_n679));
  NAND3_X1  g478(.A1(new_n678), .A2(KEYINPUT42), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT101), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(KEYINPUT42), .B1(new_n678), .B2(new_n679), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT100), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(new_n678), .B2(new_n242), .ZN(new_n685));
  OAI211_X1 g484(.A(KEYINPUT100), .B(G8gat), .C1(new_n675), .C2(new_n459), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n683), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n682), .A2(new_n687), .ZN(G1325gat));
  INV_X1    g487(.A(new_n569), .ZN(new_n689));
  OAI21_X1  g488(.A(G15gat), .B1(new_n675), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n528), .A2(new_n244), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n690), .B1(new_n675), .B2(new_n691), .ZN(G1326gat));
  INV_X1    g491(.A(new_n570), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n675), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT43), .B(G22gat), .Z(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1327gat));
  NAND2_X1  g495(.A1(new_n278), .A2(new_n279), .ZN(new_n697));
  INV_X1    g496(.A(new_n273), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n669), .A2(new_n670), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n647), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n598), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT102), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n533), .A2(new_n572), .A3(KEYINPUT88), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT88), .B1(new_n533), .B2(new_n572), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n699), .B(new_n706), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(G29gat), .A3(new_n526), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n710), .B(KEYINPUT45), .Z(new_n711));
  AOI21_X1  g510(.A(KEYINPUT44), .B1(new_n573), .B2(new_n598), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n575), .A2(new_n576), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n704), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n712), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT103), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n699), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n280), .A2(KEYINPUT103), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n703), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n716), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(G29gat), .B1(new_n722), .B2(new_n526), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n711), .A2(new_n723), .ZN(G1328gat));
  NOR3_X1   g523(.A1(new_n709), .A2(G36gat), .A3(new_n459), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT46), .ZN(new_n726));
  OAI21_X1  g525(.A(G36gat), .B1(new_n722), .B2(new_n459), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(G1329gat));
  NAND2_X1  g527(.A1(new_n528), .A2(new_n215), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n709), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT104), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(G43gat), .B1(new_n722), .B2(new_n689), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT47), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1330gat));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n716), .A2(new_n737), .A3(new_n570), .A4(new_n721), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n715), .B1(new_n707), .B2(new_n708), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n573), .A2(new_n598), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n714), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n739), .A2(new_n570), .A3(new_n741), .A4(new_n721), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT107), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n738), .A2(new_n743), .A3(G50gat), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT48), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n570), .A2(new_n213), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT105), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT106), .B1(new_n709), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT106), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n577), .A2(new_n750), .A3(new_n706), .A4(new_n747), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n745), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n744), .A2(new_n752), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n742), .A2(G50gat), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n709), .A2(new_n748), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n745), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT108), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n753), .A2(new_n759), .A3(new_n756), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(G1331gat));
  INV_X1    g560(.A(new_n720), .ZN(new_n762));
  NOR4_X1   g561(.A1(new_n701), .A2(new_n762), .A3(new_n598), .A4(new_n702), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n573), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(new_n526), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(new_n599), .ZN(G1332gat));
  NOR2_X1   g565(.A1(new_n764), .A2(new_n459), .ZN(new_n767));
  NOR2_X1   g566(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n768));
  AND2_X1   g567(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(new_n767), .B2(new_n768), .ZN(G1333gat));
  OAI21_X1  g570(.A(G71gat), .B1(new_n764), .B2(new_n689), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n528), .A2(new_n613), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n764), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n774), .B(new_n775), .ZN(G1334gat));
  NOR2_X1   g575(.A1(new_n764), .A2(new_n693), .ZN(new_n777));
  XOR2_X1   g576(.A(KEYINPUT110), .B(G78gat), .Z(new_n778));
  XNOR2_X1  g577(.A(new_n777), .B(new_n778), .ZN(G1335gat));
  NOR2_X1   g578(.A1(new_n762), .A2(new_n700), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n573), .A2(new_n598), .A3(new_n780), .ZN(new_n781));
  XOR2_X1   g580(.A(new_n781), .B(KEYINPUT51), .Z(new_n782));
  AND2_X1   g581(.A1(new_n782), .A2(new_n647), .ZN(new_n783));
  INV_X1    g582(.A(new_n526), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(new_n582), .A3(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n716), .A2(new_n647), .A3(new_n780), .ZN(new_n786));
  OAI21_X1  g585(.A(G85gat), .B1(new_n786), .B2(new_n526), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(G1336gat));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n782), .A2(new_n583), .A3(new_n455), .A4(new_n647), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(G92gat), .B1(new_n786), .B2(new_n459), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n790), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n792), .B(new_n794), .ZN(G1337gat));
  INV_X1    g594(.A(G99gat), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n783), .A2(new_n796), .A3(new_n528), .ZN(new_n797));
  OAI21_X1  g596(.A(G99gat), .B1(new_n786), .B2(new_n689), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(G1338gat));
  OAI21_X1  g598(.A(G106gat), .B1(new_n786), .B2(new_n693), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n693), .A2(G106gat), .A3(new_n702), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(KEYINPUT112), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n782), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g604(.A1(new_n671), .A2(new_n720), .ZN(new_n806));
  XOR2_X1   g605(.A(new_n806), .B(KEYINPUT113), .Z(new_n807));
  NOR2_X1   g606(.A1(new_n265), .A2(new_n210), .ZN(new_n808));
  AND3_X1   g607(.A1(new_n253), .A2(new_n258), .A3(new_n212), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n206), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(KEYINPUT114), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n598), .A2(new_n697), .A3(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n630), .A2(new_n632), .A3(new_n644), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n814), .A2(new_n645), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n633), .A2(new_n815), .A3(new_n634), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n642), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n813), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n639), .B1(new_n645), .B2(new_n815), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n635), .A2(KEYINPUT54), .ZN(new_n821));
  OAI211_X1 g620(.A(KEYINPUT55), .B(new_n820), .C1(new_n821), .C2(new_n814), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n819), .A2(new_n641), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n812), .A2(new_n823), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n819), .A2(new_n641), .A3(new_n822), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n718), .A2(new_n719), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n647), .A3(new_n697), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n598), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n826), .A2(KEYINPUT115), .A3(new_n827), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n824), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n701), .B1(new_n832), .B2(KEYINPUT116), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n280), .A2(KEYINPUT103), .ZN(new_n834));
  AOI211_X1 g633(.A(new_n717), .B(new_n273), .C1(new_n278), .C2(new_n279), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n834), .A2(new_n835), .A3(new_n823), .ZN(new_n836));
  INV_X1    g635(.A(new_n827), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n829), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n838), .A2(new_n704), .A3(new_n831), .ZN(new_n839));
  INV_X1    g638(.A(new_n824), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n807), .B1(new_n833), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n531), .A2(new_n526), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n459), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n848), .A2(new_n285), .A3(new_n280), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n846), .B(new_n850), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n851), .A2(new_n459), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n762), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n849), .B1(new_n853), .B2(new_n285), .ZN(G1340gat));
  INV_X1    g653(.A(G120gat), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n848), .A2(new_n855), .A3(new_n702), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n852), .A2(new_n647), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n856), .B1(new_n857), .B2(new_n855), .ZN(G1341gat));
  NAND3_X1  g657(.A1(new_n852), .A2(new_n297), .A3(new_n700), .ZN(new_n859));
  OAI21_X1  g658(.A(G127gat), .B1(new_n848), .B2(new_n701), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(G1342gat));
  INV_X1    g660(.A(G134gat), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n455), .A2(new_n704), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n851), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(KEYINPUT56), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n862), .B1(new_n847), .B2(new_n863), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n864), .A2(KEYINPUT118), .A3(KEYINPUT56), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT118), .B1(new_n864), .B2(KEYINPUT56), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(G1343gat));
  NOR3_X1   g669(.A1(new_n569), .A2(new_n526), .A3(new_n455), .ZN(new_n871));
  XOR2_X1   g670(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n873), .B1(new_n844), .B2(new_n570), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n570), .A2(KEYINPUT57), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n806), .B(KEYINPUT113), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n827), .B1(new_n280), .B2(new_n823), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n877), .A2(new_n704), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n701), .B1(new_n878), .B2(new_n824), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n876), .B1(new_n879), .B2(KEYINPUT120), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n879), .A2(KEYINPUT120), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n875), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n871), .B1(new_n874), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(G141gat), .B1(new_n883), .B2(new_n280), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT58), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n700), .B1(new_n841), .B2(new_n842), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n832), .A2(KEYINPUT116), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n876), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(new_n693), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n889), .A2(new_n871), .ZN(new_n890));
  INV_X1    g689(.A(G141gat), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n890), .A2(new_n891), .A3(new_n699), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n884), .A2(new_n885), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(G141gat), .B1(new_n883), .B2(new_n720), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n892), .ZN(new_n895));
  AOI21_X1  g694(.A(KEYINPUT121), .B1(new_n895), .B2(KEYINPUT58), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n897));
  AOI211_X1 g696(.A(new_n897), .B(new_n885), .C1(new_n894), .C2(new_n892), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n893), .B1(new_n896), .B2(new_n898), .ZN(G1344gat));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n900), .B(G148gat), .C1(new_n883), .C2(new_n702), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT123), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n693), .A2(new_n872), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n903), .B1(new_n888), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n844), .A2(KEYINPUT122), .A3(new_n904), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT57), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n673), .A2(new_n280), .A3(new_n674), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n909), .A2(new_n879), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n908), .B1(new_n910), .B2(new_n693), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n906), .A2(new_n907), .A3(new_n911), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n871), .A2(new_n647), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(G148gat), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n902), .B1(new_n915), .B2(KEYINPUT59), .ZN(new_n916));
  INV_X1    g715(.A(G148gat), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n917), .B1(new_n912), .B2(new_n913), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n918), .A2(KEYINPUT123), .A3(new_n900), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n901), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n889), .A2(new_n917), .A3(new_n913), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1345gat));
  NOR3_X1   g721(.A1(new_n883), .A2(new_n307), .A3(new_n701), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n890), .A2(new_n700), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n924), .A2(KEYINPUT124), .ZN(new_n925));
  AOI21_X1  g724(.A(G155gat), .B1(new_n924), .B2(KEYINPUT124), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(G1346gat));
  OAI21_X1  g726(.A(G162gat), .B1(new_n883), .B2(new_n704), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n890), .A2(new_n308), .A3(new_n598), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(G1347gat));
  NOR2_X1   g729(.A1(new_n784), .A2(new_n459), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n844), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n518), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n934), .A2(G169gat), .A3(new_n699), .ZN(new_n935));
  AOI21_X1  g734(.A(G169gat), .B1(new_n934), .B2(new_n762), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n935), .A2(new_n936), .ZN(G1348gat));
  NAND2_X1  g736(.A1(new_n934), .A2(new_n647), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g738(.A1(new_n934), .A2(new_n391), .A3(new_n700), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(KEYINPUT60), .ZN(new_n942));
  OAI21_X1  g741(.A(G183gat), .B1(new_n933), .B2(new_n701), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n940), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n941), .A2(KEYINPUT60), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n944), .B(new_n945), .ZN(G1350gat));
  OAI22_X1  g745(.A1(new_n933), .A2(new_n704), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n947));
  NAND2_X1  g746(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n947), .B(new_n948), .ZN(G1351gat));
  NOR2_X1   g748(.A1(new_n693), .A2(new_n569), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n932), .A2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT126), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n932), .A2(KEYINPUT126), .A3(new_n950), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n720), .A2(G197gat), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT127), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n931), .A2(new_n689), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n912), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(new_n699), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(G197gat), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n957), .A2(new_n962), .ZN(G1352gat));
  NOR3_X1   g762(.A1(new_n951), .A2(G204gat), .A3(new_n702), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT62), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n960), .A2(new_n647), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(G204gat), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n965), .A2(new_n967), .ZN(G1353gat));
  AND2_X1   g767(.A1(new_n953), .A2(new_n954), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n969), .A2(new_n385), .A3(new_n700), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n912), .A2(new_n700), .A3(new_n959), .ZN(new_n971));
  AOI21_X1  g770(.A(KEYINPUT63), .B1(new_n971), .B2(G211gat), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n971), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(G1354gat));
  AOI21_X1  g773(.A(G218gat), .B1(new_n969), .B2(new_n598), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n598), .A2(new_n380), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n975), .B1(new_n960), .B2(new_n976), .ZN(G1355gat));
endmodule


