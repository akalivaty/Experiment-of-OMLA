//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 1 0 1 0 1 0 1 0 0 0 1 1 0 1 1 1 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n813, new_n814,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933;
  INV_X1    g000(.A(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT81), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT2), .ZN(new_n204));
  AOI22_X1  g003(.A1(new_n203), .A2(new_n204), .B1(G155gat), .B2(G162gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G155gat), .B2(G162gat), .ZN(new_n206));
  INV_X1    g005(.A(G155gat), .ZN(new_n207));
  INV_X1    g006(.A(G162gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT2), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210));
  INV_X1    g009(.A(G141gat), .ZN(new_n211));
  INV_X1    g010(.A(G148gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n209), .A2(new_n210), .A3(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(new_n206), .B(new_n214), .Z(new_n215));
  OAI21_X1  g014(.A(KEYINPUT82), .B1(new_n215), .B2(KEYINPUT3), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n206), .B(new_n214), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT82), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT29), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT22), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n222), .A2(KEYINPUT77), .B1(G211gat), .B2(G218gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(KEYINPUT77), .B2(new_n222), .ZN(new_n224));
  XNOR2_X1  g023(.A(G197gat), .B(G204gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G211gat), .B(G218gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n226), .B(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT29), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT3), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI22_X1  g030(.A1(new_n221), .A2(new_n229), .B1(new_n231), .B2(new_n217), .ZN(new_n232));
  NAND2_X1  g031(.A1(G228gat), .A2(G233gat), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n233), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G78gat), .B(G106gat), .ZN(new_n237));
  INV_X1    g036(.A(G50gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n239), .B(new_n240), .Z(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n236), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT85), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n202), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n241), .B1(new_n234), .B2(new_n235), .ZN(new_n246));
  NOR3_X1   g045(.A1(new_n246), .A2(KEYINPUT85), .A3(G22gat), .ZN(new_n247));
  OAI22_X1  g046(.A1(new_n245), .A2(new_n247), .B1(new_n236), .B2(new_n242), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n243), .A2(new_n244), .A3(new_n202), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n236), .A2(new_n242), .ZN(new_n250));
  OAI21_X1  g049(.A(G22gat), .B1(new_n246), .B2(KEYINPUT85), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT28), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT27), .B(G183gat), .ZN(new_n255));
  INV_X1    g054(.A(G190gat), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n257), .B1(G183gat), .B2(G190gat), .ZN(new_n258));
  INV_X1    g057(.A(G169gat), .ZN(new_n259));
  INV_X1    g058(.A(G176gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n260), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n261), .B1(KEYINPUT26), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT66), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(G169gat), .A2(G176gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT66), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n263), .B1(new_n268), .B2(KEYINPUT26), .ZN(new_n269));
  INV_X1    g068(.A(G183gat), .ZN(new_n270));
  NOR3_X1   g069(.A1(new_n270), .A2(KEYINPUT71), .A3(KEYINPUT27), .ZN(new_n271));
  OAI21_X1  g070(.A(KEYINPUT27), .B1(new_n270), .B2(KEYINPUT71), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(new_n254), .A3(new_n256), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n258), .B(new_n269), .C1(new_n271), .C2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n265), .A2(KEYINPUT23), .A3(new_n267), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT25), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n261), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT23), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT65), .B1(new_n262), .B2(new_n278), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n262), .A2(KEYINPUT65), .A3(new_n278), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n275), .B(new_n277), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n282));
  AOI22_X1  g081(.A1(new_n282), .A2(KEYINPUT67), .B1(new_n270), .B2(new_n256), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT68), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND4_X1  g086(.A1(KEYINPUT68), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n287), .B(new_n288), .C1(KEYINPUT67), .C2(new_n282), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT69), .B1(new_n284), .B2(new_n289), .ZN(new_n290));
  AND2_X1   g089(.A1(new_n287), .A2(new_n288), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT69), .ZN(new_n292));
  OR2_X1    g091(.A1(new_n282), .A2(KEYINPUT67), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n291), .A2(new_n292), .A3(new_n283), .A4(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n281), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT70), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT64), .ZN(new_n298));
  OAI221_X1 g097(.A(new_n285), .B1(G183gat), .B2(G190gat), .C1(new_n282), .C2(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n299), .B1(new_n298), .B2(new_n282), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n261), .B1(KEYINPUT23), .B2(new_n266), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n301), .B1(new_n280), .B2(new_n279), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n276), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n303), .B1(new_n295), .B2(new_n296), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n274), .B1(new_n297), .B2(new_n304), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n305), .A2(G226gat), .A3(G233gat), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n305), .A2(new_n230), .B1(G226gat), .B2(G233gat), .ZN(new_n307));
  OR3_X1    g106(.A1(new_n306), .A2(new_n307), .A3(new_n228), .ZN(new_n308));
  XNOR2_X1  g107(.A(G8gat), .B(G36gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(G64gat), .B(G92gat), .ZN(new_n310));
  XOR2_X1   g109(.A(new_n309), .B(new_n310), .Z(new_n311));
  OAI21_X1  g110(.A(new_n228), .B1(new_n306), .B2(new_n307), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n308), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT78), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT78), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n308), .A2(new_n315), .A3(new_n311), .A4(new_n312), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n308), .A2(new_n312), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n311), .B1(new_n318), .B2(KEYINPUT37), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT37), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n308), .A2(new_n320), .A3(new_n312), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT38), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT86), .ZN(new_n324));
  INV_X1    g123(.A(G120gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G113gat), .ZN(new_n326));
  INV_X1    g125(.A(G113gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G120gat), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT1), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G127gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(KEYINPUT72), .A2(G127gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n331), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n333), .A2(G134gat), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(G134gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(new_n217), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n335), .A2(new_n215), .A3(new_n336), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(KEYINPUT83), .A3(new_n339), .ZN(new_n340));
  OR3_X1    g139(.A1(new_n337), .A2(KEYINPUT83), .A3(new_n217), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(G225gat), .A2(G233gat), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT5), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n216), .A2(new_n220), .ZN(new_n345));
  INV_X1    g144(.A(new_n336), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n346), .A2(new_n334), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n345), .B(new_n347), .C1(new_n219), .C2(new_n217), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n337), .A2(KEYINPUT4), .A3(new_n217), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT4), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n338), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n348), .A2(new_n349), .A3(new_n343), .A4(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n344), .A2(new_n352), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n351), .A2(new_n349), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n354), .A2(KEYINPUT5), .A3(new_n348), .A4(new_n343), .ZN(new_n355));
  XNOR2_X1  g154(.A(G1gat), .B(G29gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n356), .B(KEYINPUT0), .ZN(new_n357));
  XNOR2_X1  g156(.A(G57gat), .B(G85gat), .ZN(new_n358));
  XOR2_X1   g157(.A(new_n357), .B(new_n358), .Z(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n353), .A2(new_n355), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT6), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n360), .B1(new_n353), .B2(new_n355), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n324), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n353), .A2(new_n355), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n359), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n367), .A2(KEYINPUT86), .A3(new_n362), .A4(new_n361), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n353), .A2(new_n355), .A3(KEYINPUT6), .A4(new_n360), .ZN(new_n370));
  XOR2_X1   g169(.A(new_n370), .B(KEYINPUT88), .Z(new_n371));
  AND4_X1   g170(.A1(new_n317), .A2(new_n323), .A3(new_n369), .A4(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT38), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n319), .A2(new_n373), .A3(new_n321), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(KEYINPUT87), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n253), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n311), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n318), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT30), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n378), .B1(new_n379), .B2(new_n313), .ZN(new_n380));
  XOR2_X1   g179(.A(KEYINPUT79), .B(KEYINPUT30), .Z(new_n381));
  NAND3_X1  g180(.A1(new_n314), .A2(new_n316), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT80), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n314), .A2(KEYINPUT80), .A3(new_n316), .A4(new_n381), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n380), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n354), .A2(new_n348), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n387), .A2(G225gat), .A3(G233gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n342), .A2(new_n343), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(KEYINPUT39), .A3(new_n389), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n390), .B(new_n359), .C1(KEYINPUT39), .C2(new_n388), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT40), .ZN(new_n392));
  OR2_X1    g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n391), .A2(new_n392), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(new_n394), .A3(new_n361), .ZN(new_n395));
  OR2_X1    g194(.A1(new_n386), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n376), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT36), .ZN(new_n398));
  XNOR2_X1  g197(.A(G15gat), .B(G43gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(G71gat), .B(G99gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n399), .B(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n305), .A2(new_n337), .ZN(new_n402));
  INV_X1    g201(.A(G227gat), .ZN(new_n403));
  INV_X1    g202(.A(G233gat), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n347), .B(new_n274), .C1(new_n297), .C2(new_n304), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n402), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n401), .B1(new_n407), .B2(KEYINPUT32), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT73), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT33), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n407), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n409), .B1(new_n407), .B2(new_n410), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n408), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OR2_X1    g212(.A1(new_n401), .A2(new_n410), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n407), .A2(KEYINPUT32), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT74), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n407), .A2(KEYINPUT74), .A3(KEYINPUT32), .A4(new_n414), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n413), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n405), .B1(new_n402), .B2(new_n406), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT34), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n421), .A2(new_n422), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n413), .A2(new_n419), .A3(new_n425), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT75), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT76), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT75), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n413), .A2(new_n419), .A3(new_n431), .A4(new_n425), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n429), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n430), .B1(new_n429), .B2(new_n432), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n398), .B(new_n427), .C1(new_n433), .C2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n429), .A2(new_n432), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n427), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT36), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n367), .A2(new_n362), .A3(new_n361), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n370), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n386), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n253), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n397), .A2(new_n439), .A3(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n427), .B1(new_n433), .B2(new_n434), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT35), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n248), .A2(new_n447), .A3(new_n252), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n448), .B1(new_n369), .B2(new_n371), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n446), .A2(new_n386), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n253), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n451), .A2(new_n436), .A3(new_n427), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT35), .B1(new_n442), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n444), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT94), .ZN(new_n456));
  XNOR2_X1  g255(.A(G113gat), .B(G141gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n457), .B(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G169gat), .B(G197gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n459), .B(new_n460), .ZN(new_n461));
  XOR2_X1   g260(.A(new_n461), .B(KEYINPUT12), .Z(new_n462));
  NAND2_X1  g261(.A1(G229gat), .A2(G233gat), .ZN(new_n463));
  XOR2_X1   g262(.A(new_n463), .B(KEYINPUT13), .Z(new_n464));
  XNOR2_X1  g263(.A(G15gat), .B(G22gat), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT16), .ZN(new_n466));
  AOI21_X1  g265(.A(G1gat), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n202), .A2(G15gat), .ZN(new_n468));
  INV_X1    g267(.A(G15gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(G22gat), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n470), .A3(KEYINPUT92), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(G8gat), .ZN(new_n472));
  INV_X1    g271(.A(G8gat), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n465), .A2(KEYINPUT92), .A3(new_n473), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n467), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(G1gat), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n468), .A2(new_n470), .A3(new_n466), .ZN(new_n477));
  AOI22_X1  g276(.A1(new_n472), .A2(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(G43gat), .B(G50gat), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NOR3_X1   g281(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n483));
  OAI22_X1  g282(.A1(new_n480), .A2(KEYINPUT15), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n238), .A2(G43gat), .ZN(new_n485));
  INV_X1    g284(.A(G43gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(G50gat), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(new_n487), .A3(KEYINPUT15), .ZN(new_n488));
  NAND2_X1  g287(.A1(G29gat), .A2(G36gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n484), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n481), .A2(KEYINPUT90), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT90), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n493), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n495));
  INV_X1    g294(.A(G36gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n492), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n488), .B1(new_n498), .B2(new_n489), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT91), .B1(new_n491), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n487), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT15), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n497), .A2(new_n481), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n503), .A2(new_n488), .A3(new_n489), .A4(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT91), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n481), .A2(KEYINPUT90), .B1(new_n495), .B2(new_n496), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n507), .A2(new_n494), .B1(G29gat), .B2(G36gat), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n505), .B(new_n506), .C1(new_n508), .C2(new_n488), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n479), .A2(new_n500), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n479), .B1(new_n500), .B2(new_n509), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n464), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT17), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n500), .A2(new_n509), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n489), .ZN(new_n516));
  INV_X1    g315(.A(new_n488), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n501), .A2(new_n502), .B1(new_n497), .B2(new_n481), .ZN(new_n518));
  AOI22_X1  g317(.A1(new_n480), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n472), .A2(new_n474), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n477), .A2(new_n476), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n467), .A2(new_n472), .A3(new_n474), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n520), .A2(KEYINPUT17), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n515), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n526), .A2(KEYINPUT18), .A3(new_n510), .A4(new_n463), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n510), .A2(new_n463), .ZN(new_n528));
  AOI21_X1  g327(.A(KEYINPUT18), .B1(new_n528), .B2(new_n526), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT93), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n513), .B(new_n527), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n526), .A2(new_n510), .A3(new_n463), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT18), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(KEYINPUT93), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n456), .B(new_n462), .C1(new_n531), .C2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n462), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n527), .A2(new_n513), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n529), .A2(new_n530), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n537), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n527), .A2(new_n513), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n543), .A2(new_n537), .A3(new_n534), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT94), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n536), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n455), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G99gat), .A2(G106gat), .ZN(new_n549));
  INV_X1    g348(.A(G85gat), .ZN(new_n550));
  INV_X1    g349(.A(G92gat), .ZN(new_n551));
  AOI22_X1  g350(.A1(KEYINPUT8), .A2(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT97), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT7), .ZN(new_n554));
  NAND2_X1  g353(.A1(G85gat), .A2(G92gat), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n553), .B(new_n554), .C1(new_n555), .C2(KEYINPUT98), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n553), .B1(new_n555), .B2(KEYINPUT98), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n558), .B(KEYINPUT7), .C1(new_n553), .C2(new_n555), .ZN(new_n559));
  INV_X1    g358(.A(new_n549), .ZN(new_n560));
  NOR2_X1   g359(.A1(G99gat), .A2(G106gat), .ZN(new_n561));
  OAI21_X1  g360(.A(KEYINPUT99), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n561), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT99), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n564), .A3(new_n549), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n557), .A2(new_n559), .A3(new_n562), .A4(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(G85gat), .A2(G92gat), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT98), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT97), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT7), .B1(new_n555), .B2(new_n553), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n556), .B(new_n552), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n565), .A2(new_n562), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AND4_X1   g372(.A1(new_n500), .A2(new_n509), .A3(new_n566), .A4(new_n573), .ZN(new_n574));
  AND2_X1   g373(.A1(G232gat), .A2(G233gat), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n574), .B1(KEYINPUT41), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n520), .A2(KEYINPUT17), .B1(new_n566), .B2(new_n573), .ZN(new_n577));
  AND3_X1   g376(.A1(new_n515), .A2(KEYINPUT100), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT100), .B1(new_n515), .B2(new_n577), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n576), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G190gat), .B(G218gat), .Z(new_n581));
  OR2_X1    g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n575), .A2(KEYINPUT41), .ZN(new_n583));
  XNOR2_X1  g382(.A(G134gat), .B(G162gat), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n583), .B(new_n584), .Z(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n580), .A2(new_n581), .ZN(new_n587));
  AND4_X1   g386(.A1(KEYINPUT101), .A2(new_n582), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n585), .B(KEYINPUT101), .Z(new_n589));
  AOI21_X1  g388(.A(new_n589), .B1(new_n582), .B2(new_n587), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G71gat), .A2(G78gat), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT95), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(G71gat), .A2(G78gat), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT95), .B1(G71gat), .B2(G78gat), .ZN(new_n597));
  NOR3_X1   g396(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(G57gat), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n599), .A2(G64gat), .ZN(new_n600));
  INV_X1    g399(.A(G64gat), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n601), .A2(G57gat), .ZN(new_n602));
  OAI22_X1  g401(.A1(new_n600), .A2(new_n602), .B1(new_n594), .B2(KEYINPUT9), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT96), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n605), .B1(new_n599), .B2(G64gat), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n601), .A2(KEYINPUT96), .A3(G57gat), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n606), .B(new_n607), .C1(G57gat), .C2(new_n601), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n596), .A2(KEYINPUT9), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(new_n593), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n604), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT21), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(G127gat), .ZN(new_n617));
  AOI22_X1  g416(.A1(new_n603), .A2(new_n598), .B1(new_n608), .B2(new_n610), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n479), .B1(KEYINPUT21), .B2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n617), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(G155gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(G183gat), .B(G211gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n620), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G120gat), .B(G148gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(G176gat), .B(G204gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G230gat), .A2(G233gat), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n571), .A2(new_n572), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n571), .A2(new_n572), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n612), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT10), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n566), .A2(new_n618), .A3(new_n573), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n638), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(KEYINPUT10), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n633), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n632), .B1(new_n636), .B2(new_n638), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n631), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT104), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n642), .A2(new_n643), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n645), .B1(new_n646), .B2(new_n630), .ZN(new_n647));
  NOR4_X1   g446(.A1(new_n642), .A2(new_n643), .A3(KEYINPUT104), .A4(new_n631), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n644), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n592), .A2(new_n625), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n548), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n441), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G1gat), .ZN(G1324gat));
  AOI22_X1  g454(.A1(new_n376), .A2(new_n396), .B1(new_n442), .B2(new_n253), .ZN(new_n656));
  AOI22_X1  g455(.A1(new_n656), .A2(new_n439), .B1(new_n453), .B2(new_n450), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n657), .A2(new_n386), .A3(new_n546), .ZN(new_n658));
  INV_X1    g457(.A(new_n651), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT16), .B(G8gat), .Z(new_n660));
  AND3_X1   g459(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n661), .A2(KEYINPUT105), .A3(KEYINPUT42), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT42), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n658), .A2(new_n659), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n663), .B1(new_n664), .B2(G8gat), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n665), .A2(new_n661), .ZN(new_n666));
  AOI21_X1  g465(.A(KEYINPUT105), .B1(new_n661), .B2(KEYINPUT42), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n662), .B1(new_n666), .B2(new_n667), .ZN(G1325gat));
  NAND3_X1  g467(.A1(new_n652), .A2(new_n469), .A3(new_n446), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n548), .A2(new_n439), .A3(new_n651), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n669), .B1(new_n670), .B2(new_n469), .ZN(G1326gat));
  NAND2_X1  g470(.A1(new_n652), .A2(new_n253), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT43), .B(G22gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(G1327gat));
  NAND2_X1  g473(.A1(new_n455), .A2(new_n591), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n625), .A2(new_n649), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n677), .A2(new_n546), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NOR4_X1   g478(.A1(new_n675), .A2(G29gat), .A3(new_n441), .A4(new_n679), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n680), .B(KEYINPUT45), .Z(new_n681));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(new_n657), .B2(new_n592), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n592), .B1(new_n444), .B2(new_n454), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT44), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n678), .ZN(new_n687));
  OAI21_X1  g486(.A(G29gat), .B1(new_n687), .B2(new_n441), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n681), .A2(new_n688), .ZN(G1328gat));
  NOR2_X1   g488(.A1(new_n677), .A2(new_n592), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n658), .A2(new_n496), .A3(new_n690), .ZN(new_n691));
  XOR2_X1   g490(.A(new_n691), .B(KEYINPUT46), .Z(new_n692));
  OAI21_X1  g491(.A(G36gat), .B1(new_n687), .B2(new_n386), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(G1329gat));
  NAND3_X1  g493(.A1(new_n446), .A2(new_n486), .A3(new_n690), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n548), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n435), .A2(new_n438), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n683), .A2(new_n685), .A3(new_n697), .A4(new_n678), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n696), .B1(new_n698), .B2(G43gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g499(.A1(new_n683), .A2(new_n685), .A3(new_n253), .A4(new_n678), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT106), .B1(new_n701), .B2(G50gat), .ZN(new_n702));
  AND4_X1   g501(.A1(new_n238), .A2(new_n684), .A3(new_n253), .A4(new_n678), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n703), .B1(new_n701), .B2(G50gat), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT48), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n702), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  AOI221_X4 g505(.A(new_n703), .B1(KEYINPUT106), .B2(KEYINPUT48), .C1(new_n701), .C2(G50gat), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(G1331gat));
  INV_X1    g507(.A(new_n625), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(new_n547), .A3(new_n591), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n455), .A2(new_n710), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n711), .A2(new_n649), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n653), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g513(.A1(new_n386), .A2(new_n650), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n716), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n717));
  XOR2_X1   g516(.A(KEYINPUT49), .B(G64gat), .Z(new_n718));
  OAI21_X1  g517(.A(new_n717), .B1(new_n716), .B2(new_n718), .ZN(G1333gat));
  NAND4_X1  g518(.A1(new_n455), .A2(new_n446), .A3(new_n649), .A4(new_n710), .ZN(new_n720));
  OR2_X1    g519(.A1(new_n720), .A2(KEYINPUT107), .ZN(new_n721));
  AOI21_X1  g520(.A(G71gat), .B1(new_n720), .B2(KEYINPUT107), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n697), .A2(G71gat), .ZN(new_n723));
  AOI22_X1  g522(.A1(new_n721), .A2(new_n722), .B1(new_n712), .B2(new_n723), .ZN(new_n724));
  XOR2_X1   g523(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1334gat));
  NAND2_X1  g525(.A1(new_n712), .A2(new_n253), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g527(.A1(new_n709), .A2(new_n546), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT109), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n649), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n731), .B(KEYINPUT110), .Z(new_n732));
  NAND2_X1  g531(.A1(new_n686), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G85gat), .B1(new_n733), .B2(new_n441), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n684), .A2(KEYINPUT51), .A3(new_n730), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT51), .B1(new_n684), .B2(new_n730), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n653), .A2(new_n550), .A3(new_n649), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n734), .B1(new_n738), .B2(new_n739), .ZN(G1336gat));
  OAI21_X1  g539(.A(new_n715), .B1(new_n736), .B2(new_n737), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n551), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n386), .A2(new_n551), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n683), .A2(new_n685), .A3(new_n732), .A4(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT52), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(KEYINPUT111), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n745), .A2(KEYINPUT111), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n742), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n750), .B1(new_n742), .B2(new_n748), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n751), .A2(new_n752), .ZN(G1337gat));
  OAI21_X1  g552(.A(G99gat), .B1(new_n733), .B2(new_n439), .ZN(new_n754));
  OR3_X1    g553(.A1(new_n445), .A2(G99gat), .A3(new_n650), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n754), .B1(new_n738), .B2(new_n755), .ZN(G1338gat));
  NAND4_X1  g555(.A1(new_n683), .A2(new_n685), .A3(new_n253), .A4(new_n732), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(G106gat), .ZN(new_n758));
  OR3_X1    g557(.A1(new_n451), .A2(G106gat), .A3(new_n650), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n758), .B1(new_n738), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g560(.A1(new_n529), .A2(new_n462), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n511), .A2(new_n512), .A3(new_n464), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n463), .B1(new_n526), .B2(new_n510), .ZN(new_n764));
  OR2_X1    g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI22_X1  g564(.A1(new_n762), .A2(new_n543), .B1(new_n765), .B2(new_n461), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n649), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n639), .A2(new_n641), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n632), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n639), .A2(new_n641), .A3(new_n633), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n769), .A2(KEYINPUT54), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n630), .B1(new_n642), .B2(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n771), .A2(new_n773), .A3(KEYINPUT55), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT113), .ZN(new_n775));
  INV_X1    g574(.A(new_n643), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n769), .A2(new_n776), .A3(new_n630), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT104), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n646), .A2(new_n645), .A3(new_n630), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n771), .A2(new_n773), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n771), .A2(new_n773), .A3(new_n784), .A4(KEYINPUT55), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n775), .A2(new_n780), .A3(new_n783), .A4(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n767), .B1(new_n546), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI211_X1 g588(.A(KEYINPUT115), .B(new_n767), .C1(new_n546), .C2(new_n786), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(new_n592), .A3(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n461), .B1(new_n763), .B2(new_n764), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n544), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT114), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  AND3_X1   g594(.A1(new_n775), .A2(new_n780), .A3(new_n785), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n795), .A2(new_n591), .A3(new_n783), .A4(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n625), .B1(new_n791), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n651), .A2(new_n547), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n386), .ZN(new_n801));
  NOR4_X1   g600(.A1(new_n800), .A2(new_n452), .A3(new_n801), .A4(new_n441), .ZN(new_n802));
  AOI21_X1  g601(.A(G113gat), .B1(new_n802), .B2(new_n547), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n800), .A2(new_n253), .ZN(new_n804));
  AOI211_X1 g603(.A(new_n380), .B(new_n441), .C1(new_n384), .C2(new_n385), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n804), .A2(new_n446), .A3(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n546), .A2(new_n327), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n803), .B1(new_n807), .B2(new_n808), .ZN(G1340gat));
  AOI21_X1  g608(.A(G120gat), .B1(new_n802), .B2(new_n649), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n650), .A2(new_n325), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n810), .B1(new_n807), .B2(new_n811), .ZN(G1341gat));
  OAI21_X1  g611(.A(G127gat), .B1(new_n806), .B2(new_n709), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n802), .A2(new_n330), .A3(new_n625), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(G1342gat));
  XOR2_X1   g614(.A(KEYINPUT72), .B(G134gat), .Z(new_n816));
  NAND4_X1  g615(.A1(new_n386), .A2(new_n653), .A3(new_n591), .A4(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n800), .A2(new_n452), .A3(new_n817), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT56), .ZN(new_n819));
  OAI21_X1  g618(.A(G134gat), .B1(new_n806), .B2(new_n592), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(G1343gat));
  INV_X1    g620(.A(KEYINPUT58), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n435), .A2(new_n438), .A3(new_n805), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n253), .B1(new_n798), .B2(new_n799), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n825), .A2(new_n211), .A3(new_n547), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n253), .A2(KEYINPUT57), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n659), .A2(new_n546), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n542), .A2(new_n545), .ZN(new_n829));
  XOR2_X1   g628(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n830));
  NAND2_X1  g629(.A1(new_n781), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n829), .A2(new_n796), .A3(new_n536), .A4(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT116), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n649), .A2(new_n766), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n833), .B1(new_n649), .B2(new_n766), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n591), .B1(new_n832), .B2(new_n836), .ZN(new_n837));
  NOR4_X1   g636(.A1(new_n794), .A2(new_n588), .A3(new_n590), .A4(new_n786), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n709), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n827), .B1(new_n828), .B2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n824), .B2(new_n841), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n842), .A2(new_n546), .A3(new_n823), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n822), .B(new_n826), .C1(new_n843), .C2(new_n211), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT119), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT118), .B1(new_n842), .B2(new_n823), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847));
  INV_X1    g646(.A(new_n823), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n591), .B1(new_n787), .B2(new_n788), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n838), .B1(new_n790), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n828), .B1(new_n850), .B2(new_n625), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT57), .B1(new_n851), .B2(new_n253), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n847), .B(new_n848), .C1(new_n852), .C2(new_n840), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n846), .A2(new_n547), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(G141gat), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n826), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n845), .B1(new_n856), .B2(KEYINPUT58), .ZN(new_n857));
  INV_X1    g656(.A(new_n826), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n858), .B1(new_n854), .B2(G141gat), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n859), .A2(KEYINPUT119), .A3(new_n822), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n844), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g662(.A(KEYINPUT120), .B(new_n844), .C1(new_n857), .C2(new_n860), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(G1344gat));
  NOR2_X1   g664(.A1(new_n212), .A2(KEYINPUT59), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n846), .A2(new_n853), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n866), .B1(new_n867), .B2(new_n650), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n451), .B1(new_n828), .B2(new_n839), .ZN(new_n869));
  OAI22_X1  g668(.A1(new_n800), .A2(new_n827), .B1(new_n869), .B2(KEYINPUT57), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n870), .A2(new_n649), .A3(new_n848), .ZN(new_n871));
  OAI21_X1  g670(.A(KEYINPUT59), .B1(new_n871), .B2(new_n212), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n825), .A2(new_n212), .A3(new_n649), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1345gat));
  OAI21_X1  g674(.A(G155gat), .B1(new_n867), .B2(new_n709), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n825), .A2(new_n207), .A3(new_n625), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1346gat));
  NOR3_X1   g677(.A1(new_n867), .A2(new_n208), .A3(new_n592), .ZN(new_n879));
  AOI21_X1  g678(.A(G162gat), .B1(new_n825), .B2(new_n591), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n879), .A2(new_n880), .ZN(G1347gat));
  NAND4_X1  g680(.A1(new_n804), .A2(new_n441), .A3(new_n446), .A4(new_n801), .ZN(new_n882));
  OAI21_X1  g681(.A(G169gat), .B1(new_n882), .B2(new_n546), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT122), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n851), .A2(new_n441), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT121), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n452), .A2(new_n386), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n259), .A3(new_n547), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n884), .A2(new_n889), .ZN(G1348gat));
  NAND3_X1  g689(.A1(new_n888), .A2(new_n260), .A3(new_n649), .ZN(new_n891));
  OAI21_X1  g690(.A(G176gat), .B1(new_n882), .B2(new_n650), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(G1349gat));
  NAND3_X1  g692(.A1(new_n888), .A2(new_n255), .A3(new_n625), .ZN(new_n894));
  OAI21_X1  g693(.A(G183gat), .B1(new_n882), .B2(new_n709), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT60), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(KEYINPUT123), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n896), .B(new_n898), .ZN(G1350gat));
  OAI21_X1  g698(.A(G190gat), .B1(new_n882), .B2(new_n592), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT61), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n888), .A2(new_n256), .A3(new_n591), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1351gat));
  NOR3_X1   g702(.A1(new_n697), .A2(new_n386), .A3(new_n451), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT124), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n546), .A2(G197gat), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n905), .A2(new_n886), .A3(new_n906), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n907), .A2(KEYINPUT125), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n697), .A2(new_n653), .A3(new_n386), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n909), .A2(new_n870), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(G197gat), .B1(new_n911), .B2(new_n546), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n907), .A2(new_n912), .A3(KEYINPUT125), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n908), .A2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n914), .B(new_n915), .ZN(G1352gat));
  NAND2_X1  g715(.A1(new_n905), .A2(new_n886), .ZN(new_n917));
  OR3_X1    g716(.A1(new_n917), .A2(G204gat), .A3(new_n650), .ZN(new_n918));
  OR2_X1    g717(.A1(new_n918), .A2(KEYINPUT62), .ZN(new_n919));
  OAI21_X1  g718(.A(G204gat), .B1(new_n911), .B2(new_n650), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(KEYINPUT62), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(G1353gat));
  INV_X1    g721(.A(G211gat), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT63), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(KEYINPUT127), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n925), .B1(new_n911), .B2(new_n709), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n924), .A2(KEYINPUT127), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n625), .A2(new_n923), .ZN(new_n930));
  OAI22_X1  g729(.A1(new_n928), .A2(new_n929), .B1(new_n917), .B2(new_n930), .ZN(G1354gat));
  OAI21_X1  g730(.A(G218gat), .B1(new_n911), .B2(new_n592), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n592), .A2(G218gat), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n917), .B2(new_n933), .ZN(G1355gat));
endmodule


