//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n444, new_n445, new_n447, new_n451, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n562, new_n564, new_n565, new_n567,
    new_n568, new_n569, new_n570, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n607, new_n609, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1153, new_n1154,
    new_n1155, new_n1156;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  INV_X1    g017(.A(G2072), .ZN(new_n443));
  INV_X1    g018(.A(G2078), .ZN(new_n444));
  NOR2_X1   g019(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g020(.A1(new_n445), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g023(.A(G452), .Z(G391));
  AND2_X1   g024(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g027(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR4_X1   g032(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n457), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  NAND2_X1  g036(.A1(new_n457), .A2(G2106), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n459), .A2(G567), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n466), .B1(KEYINPUT3), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT67), .B(KEYINPUT3), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n469), .B2(new_n467), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT67), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(new_n466), .A3(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(G2105), .B1(new_n470), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G137), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n471), .A2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(G125), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n479), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n467), .A2(G2105), .ZN(new_n485));
  AOI22_X1  g060(.A1(new_n484), .A2(G2105), .B1(G101), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n478), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G160));
  NAND2_X1  g063(.A1(new_n477), .A2(G136), .ZN(new_n489));
  INV_X1    g064(.A(G2105), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(new_n470), .B2(new_n476), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G124), .ZN(new_n492));
  OR2_X1    g067(.A1(G100), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G112), .C2(new_n490), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n489), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n490), .A2(G138), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n482), .A2(KEYINPUT4), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n498), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n480), .A2(KEYINPUT68), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n501), .B1(new_n475), .B2(G2104), .ZN(new_n502));
  AOI211_X1 g077(.A(KEYINPUT68), .B(new_n467), .C1(new_n472), .C2(new_n474), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n500), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n499), .B1(new_n504), .B2(KEYINPUT4), .ZN(new_n505));
  OAI211_X1 g080(.A(G126), .B(G2105), .C1(new_n502), .C2(new_n503), .ZN(new_n506));
  OAI21_X1  g081(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n507));
  INV_X1    g082(.A(G114), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(G2105), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n497), .B1(new_n505), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n499), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n498), .B1(new_n470), .B2(new_n476), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT4), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n509), .B1(new_n491), .B2(G126), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT69), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n512), .A2(new_n518), .ZN(G164));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n520), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n522), .A2(KEYINPUT70), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(KEYINPUT70), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT5), .B(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n523), .A2(new_n524), .B1(G88), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT71), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n528), .A2(new_n529), .ZN(new_n532));
  INV_X1    g107(.A(G651), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n525), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n531), .A2(new_n532), .B1(new_n533), .B2(new_n534), .ZN(G303));
  INV_X1    g110(.A(G303), .ZN(G166));
  NAND2_X1  g111(.A1(new_n527), .A2(G89), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n540));
  INV_X1    g115(.A(new_n521), .ZN(new_n541));
  INV_X1    g116(.A(G51), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI211_X1 g118(.A(new_n537), .B(new_n539), .C1(new_n543), .C2(KEYINPUT72), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n543), .A2(KEYINPUT72), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n544), .A2(new_n545), .ZN(G286));
  INV_X1    g121(.A(G286), .ZN(G168));
  NAND2_X1  g122(.A1(new_n521), .A2(G52), .ZN(new_n548));
  INV_X1    g123(.A(G90), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n549), .B2(new_n526), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(new_n533), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n550), .A2(new_n552), .ZN(G171));
  AOI22_X1  g128(.A1(new_n525), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n554), .A2(new_n533), .ZN(new_n555));
  INV_X1    g130(.A(G43), .ZN(new_n556));
  INV_X1    g131(.A(G81), .ZN(new_n557));
  OAI221_X1 g132(.A(new_n555), .B1(new_n556), .B2(new_n541), .C1(new_n557), .C2(new_n526), .ZN(new_n558));
  INV_X1    g133(.A(G860), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT73), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT74), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(G188));
  NAND2_X1  g141(.A1(new_n521), .A2(G53), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n527), .A2(G91), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n525), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n570));
  OAI211_X1 g145(.A(new_n568), .B(new_n569), .C1(new_n533), .C2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  OR2_X1    g147(.A1(new_n525), .A2(G74), .ZN(new_n573));
  AOI22_X1  g148(.A1(G651), .A2(new_n573), .B1(new_n521), .B2(G49), .ZN(new_n574));
  INV_X1    g149(.A(G87), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n575), .B2(new_n526), .ZN(new_n576));
  XOR2_X1   g151(.A(new_n576), .B(KEYINPUT75), .Z(G288));
  AOI22_X1  g152(.A1(new_n525), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n578), .A2(new_n533), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n521), .A2(G48), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  AOI211_X1 g156(.A(new_n579), .B(new_n581), .C1(G86), .C2(new_n527), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G305));
  NAND2_X1  g158(.A1(new_n521), .A2(G47), .ZN(new_n584));
  INV_X1    g159(.A(G85), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n585), .B2(new_n526), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n533), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n586), .A2(new_n588), .ZN(G290));
  INV_X1    g164(.A(G868), .ZN(new_n590));
  NOR2_X1   g165(.A1(G301), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n527), .A2(G92), .ZN(new_n592));
  XOR2_X1   g167(.A(new_n592), .B(KEYINPUT10), .Z(new_n593));
  NAND2_X1  g168(.A1(new_n525), .A2(G66), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n533), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n596), .B1(G54), .B2(new_n521), .ZN(new_n597));
  AND3_X1   g172(.A1(new_n593), .A2(KEYINPUT76), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(KEYINPUT76), .B1(new_n593), .B2(new_n597), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n591), .B1(new_n601), .B2(new_n590), .ZN(G284));
  AOI21_X1  g177(.A(new_n591), .B1(new_n601), .B2(new_n590), .ZN(G321));
  NAND2_X1  g178(.A1(G299), .A2(new_n590), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G168), .B2(new_n590), .ZN(G297));
  OAI21_X1  g180(.A(new_n604), .B1(G168), .B2(new_n590), .ZN(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n601), .B1(new_n607), .B2(G860), .ZN(G148));
  NAND2_X1  g183(.A1(new_n601), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(new_n558), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(G868), .B2(new_n611), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n491), .A2(G123), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n490), .A2(G111), .ZN(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(G135), .B2(new_n477), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT77), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2096), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n490), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT12), .Z(new_n622));
  XOR2_X1   g197(.A(KEYINPUT13), .B(G2100), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n620), .A2(new_n624), .ZN(G156));
  INV_X1    g200(.A(KEYINPUT14), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2427), .B(G2438), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2430), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT15), .B(G2435), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n626), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(new_n629), .B2(new_n628), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(G1341), .B(G1348), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n631), .B(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2443), .B(G2446), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(G14), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n640), .B1(new_n639), .B2(new_n637), .ZN(G401));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT78), .ZN(new_n643));
  XOR2_X1   g218(.A(G2072), .B(G2078), .Z(new_n644));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  NOR3_X1   g221(.A1(new_n643), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT18), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n643), .A2(new_n644), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n644), .B(KEYINPUT17), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n649), .B(new_n646), .C1(new_n643), .C2(new_n650), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(new_n643), .A3(new_n645), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n648), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2096), .B(G2100), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT79), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n653), .B(new_n655), .ZN(G227));
  XOR2_X1   g231(.A(G1971), .B(G1976), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1956), .B(G2474), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1961), .B(G1966), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n658), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n658), .A2(new_n661), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT20), .Z(new_n665));
  NAND2_X1  g240(.A1(new_n658), .A2(new_n662), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(KEYINPUT80), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(KEYINPUT80), .ZN(new_n668));
  AOI211_X1 g243(.A(new_n663), .B(new_n665), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1991), .B(G1996), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1981), .B(G1986), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G229));
  INV_X1    g250(.A(G16), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(G22), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT84), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(G166), .B2(new_n676), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n679), .A2(G1971), .ZN(new_n680));
  NOR2_X1   g255(.A1(G6), .A2(G16), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n582), .B2(G16), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT32), .ZN(new_n683));
  INV_X1    g258(.A(G1981), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n679), .A2(G1971), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n676), .A2(G23), .ZN(new_n687));
  INV_X1    g262(.A(new_n576), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n688), .B2(new_n676), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT33), .B(G1976), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND4_X1  g266(.A1(new_n680), .A2(new_n685), .A3(new_n686), .A4(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT83), .B(KEYINPUT34), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  INV_X1    g271(.A(G29), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G25), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT81), .Z(new_n699));
  OR2_X1    g274(.A1(new_n490), .A2(G107), .ZN(new_n700));
  OAI21_X1  g275(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  AOI22_X1  g277(.A1(new_n491), .A2(G119), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n477), .A2(G131), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n699), .B1(new_n705), .B2(G29), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT82), .Z(new_n707));
  XOR2_X1   g282(.A(KEYINPUT35), .B(G1991), .Z(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n707), .A2(new_n709), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n676), .A2(G24), .ZN(new_n712));
  INV_X1    g287(.A(G290), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(new_n676), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G1986), .ZN(new_n715));
  NOR3_X1   g290(.A1(new_n710), .A2(new_n711), .A3(new_n715), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n695), .A2(new_n696), .A3(new_n716), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT85), .B(KEYINPUT36), .Z(new_n718));
  AND2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n717), .A2(new_n718), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n676), .A2(G21), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G168), .B2(new_n676), .ZN(new_n722));
  INV_X1    g297(.A(G1966), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n601), .A2(G16), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G4), .B2(G16), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT86), .B(G1348), .Z(new_n727));
  OAI21_X1  g302(.A(new_n724), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n676), .A2(G20), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT23), .Z(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G299), .B2(G16), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1956), .ZN(new_n732));
  INV_X1    g307(.A(G34), .ZN(new_n733));
  AOI21_X1  g308(.A(G29), .B1(new_n733), .B2(KEYINPUT24), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(KEYINPUT24), .B2(new_n733), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n487), .B2(new_n697), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G2084), .ZN(new_n737));
  NOR2_X1   g312(.A1(G16), .A2(G19), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n611), .B2(G16), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(G1341), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT30), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n741), .A2(G28), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n697), .B1(new_n741), .B2(G28), .ZN(new_n743));
  AND2_X1   g318(.A1(KEYINPUT31), .A2(G11), .ZN(new_n744));
  NOR2_X1   g319(.A1(KEYINPUT31), .A2(G11), .ZN(new_n745));
  OAI22_X1  g320(.A1(new_n742), .A2(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n740), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(G5), .A2(G16), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT88), .Z(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G301), .B2(new_n676), .ZN(new_n750));
  INV_X1    g325(.A(G1961), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n739), .A2(G1341), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n732), .A2(new_n737), .A3(new_n747), .A4(new_n752), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n728), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n697), .A2(G32), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n477), .A2(G141), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n491), .A2(G129), .ZN(new_n757));
  NAND3_X1  g332(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT26), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n760), .A2(new_n761), .B1(G105), .B2(new_n485), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n756), .A2(new_n757), .A3(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n755), .B1(new_n764), .B2(new_n697), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT27), .B(G1996), .Z(new_n766));
  NOR2_X1   g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n726), .B2(new_n727), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n697), .A2(G35), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G162), .B2(new_n697), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT29), .Z(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G2090), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n619), .A2(G29), .B1(new_n765), .B2(new_n766), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n768), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G27), .A2(G29), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G164), .B2(G29), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G2078), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n750), .A2(new_n751), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT89), .Z(new_n780));
  NAND2_X1  g355(.A1(new_n697), .A2(G26), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT28), .Z(new_n782));
  NAND2_X1  g357(.A1(new_n477), .A2(G140), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n491), .A2(G128), .ZN(new_n784));
  OR2_X1    g359(.A1(G104), .A2(G2105), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n785), .B(G2104), .C1(G116), .C2(new_n490), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n783), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n782), .B1(new_n787), .B2(G29), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G2067), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n477), .A2(G139), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT87), .B(KEYINPUT25), .Z(new_n791));
  NAND3_X1  g366(.A1(new_n490), .A2(G103), .A3(G2104), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  NAND2_X1  g369(.A1(G115), .A2(G2104), .ZN(new_n795));
  INV_X1    g370(.A(G127), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n795), .B1(new_n482), .B2(new_n796), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n793), .A2(new_n794), .B1(G2105), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n790), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(G29), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G29), .B2(G33), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(new_n443), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n443), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n780), .A2(new_n789), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  NOR4_X1   g380(.A1(new_n754), .A2(new_n775), .A3(new_n778), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n772), .A2(G2090), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT90), .Z(new_n808));
  NAND2_X1  g383(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n719), .A2(new_n720), .A3(new_n809), .ZN(G311));
  INV_X1    g385(.A(G311), .ZN(G150));
  NOR2_X1   g386(.A1(new_n600), .A2(new_n607), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT38), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n527), .A2(G93), .B1(new_n521), .B2(G55), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n525), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(new_n533), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n558), .B(new_n817), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n813), .B(new_n818), .Z(new_n819));
  OR2_X1    g394(.A1(new_n819), .A2(KEYINPUT39), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(KEYINPUT39), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n820), .A2(new_n559), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n817), .A2(new_n559), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT37), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(G145));
  INV_X1    g400(.A(KEYINPUT91), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n516), .A2(new_n826), .ZN(new_n827));
  OAI211_X1 g402(.A(KEYINPUT91), .B(new_n513), .C1(new_n514), .C2(new_n515), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n511), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(new_n787), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(new_n799), .ZN(new_n831));
  INV_X1    g406(.A(new_n787), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n829), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(new_n800), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(new_n763), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n831), .A2(new_n834), .A3(new_n764), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n477), .A2(G142), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n491), .A2(G130), .ZN(new_n839));
  OR2_X1    g414(.A1(G106), .A2(G2105), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n840), .B(G2104), .C1(G118), .C2(new_n490), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  AND3_X1   g418(.A1(new_n703), .A2(KEYINPUT92), .A3(new_n704), .ZN(new_n844));
  AOI21_X1  g419(.A(KEYINPUT92), .B1(new_n703), .B2(new_n704), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n622), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n622), .B1(new_n844), .B2(new_n845), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n843), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n848), .A2(new_n843), .A3(new_n849), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n851), .A2(KEYINPUT93), .A3(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT93), .ZN(new_n854));
  INV_X1    g429(.A(new_n852), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n855), .B2(new_n850), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n836), .A2(new_n837), .A3(new_n853), .A4(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT95), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n858), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n836), .A2(new_n837), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n856), .A2(new_n853), .ZN(new_n862));
  AOI21_X1  g437(.A(KEYINPUT94), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AND3_X1   g438(.A1(new_n861), .A2(KEYINPUT94), .A3(new_n862), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n859), .B(new_n860), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n619), .B(G160), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n495), .ZN(new_n867));
  AOI21_X1  g442(.A(KEYINPUT96), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n865), .A2(KEYINPUT96), .A3(new_n867), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n864), .A2(new_n863), .ZN(new_n872));
  NOR3_X1   g447(.A1(new_n861), .A2(new_n855), .A3(new_n850), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n873), .A2(new_n867), .ZN(new_n874));
  AOI21_X1  g449(.A(G37), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(KEYINPUT40), .B1(new_n871), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n870), .ZN(new_n877));
  OAI211_X1 g452(.A(KEYINPUT40), .B(new_n875), .C1(new_n877), .C2(new_n868), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n876), .A2(new_n879), .ZN(G395));
  NAND2_X1  g455(.A1(G166), .A2(new_n582), .ZN(new_n881));
  NAND2_X1  g456(.A1(G303), .A2(G305), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n688), .B(G290), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT98), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n881), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n883), .A2(new_n884), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n886), .A2(new_n884), .A3(new_n883), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT42), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n888), .A2(KEYINPUT42), .A3(new_n889), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n609), .B(new_n818), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n593), .A2(new_n597), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n896), .B(G299), .Z(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT41), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  XOR2_X1   g475(.A(KEYINPUT97), .B(KEYINPUT41), .Z(new_n901));
  OAI21_X1  g476(.A(new_n900), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n894), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n898), .A2(new_n903), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n892), .B(new_n893), .C1(new_n904), .C2(KEYINPUT99), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(KEYINPUT99), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n904), .A2(new_n892), .A3(KEYINPUT99), .A4(new_n893), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n590), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n817), .A2(G868), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(G295));
  OR3_X1    g488(.A1(new_n909), .A2(KEYINPUT100), .A3(new_n911), .ZN(new_n914));
  OAI21_X1  g489(.A(KEYINPUT100), .B1(new_n909), .B2(new_n911), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(G331));
  XNOR2_X1  g491(.A(new_n818), .B(G171), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(G286), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n897), .A2(new_n901), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n919), .B(KEYINPUT103), .C1(new_n899), .C2(new_n897), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n918), .B(new_n920), .C1(KEYINPUT103), .C2(new_n919), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n917), .B(G168), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n897), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n921), .A2(KEYINPUT104), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n890), .A2(new_n925), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n923), .A2(KEYINPUT104), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n888), .A2(KEYINPUT102), .A3(new_n889), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n924), .A2(new_n926), .A3(new_n927), .A4(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(G37), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n918), .A2(new_n902), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n923), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n930), .B1(new_n932), .B2(new_n890), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n929), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT43), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT43), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n926), .A2(new_n928), .A3(new_n932), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n934), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT106), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  OAI211_X1 g517(.A(KEYINPUT44), .B(new_n936), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n926), .A2(new_n928), .A3(new_n932), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT43), .B1(new_n944), .B2(new_n933), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n929), .A2(new_n934), .A3(new_n937), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  XOR2_X1   g522(.A(KEYINPUT101), .B(KEYINPUT44), .Z(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT105), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n951));
  AOI211_X1 g526(.A(new_n951), .B(new_n948), .C1(new_n945), .C2(new_n946), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n943), .B1(new_n950), .B2(new_n952), .ZN(G397));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(new_n829), .B2(G1384), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(G160), .A2(G40), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G1996), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(KEYINPUT46), .A3(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n962), .B(KEYINPUT125), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT46), .B1(new_n960), .B2(new_n961), .ZN(new_n964));
  INV_X1    g539(.A(G2067), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n787), .B(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n959), .B1(new_n764), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n963), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n969), .B(KEYINPUT47), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n705), .A2(new_n709), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n971), .B(KEYINPUT124), .Z(new_n972));
  XNOR2_X1  g547(.A(new_n763), .B(new_n961), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n973), .A2(new_n966), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n832), .A2(new_n965), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n959), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n959), .A2(G1986), .A3(G290), .ZN(new_n978));
  OR2_X1    g553(.A1(new_n978), .A2(KEYINPUT48), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n705), .B(new_n708), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n974), .A2(new_n980), .ZN(new_n981));
  AOI22_X1  g556(.A1(new_n978), .A2(KEYINPUT48), .B1(new_n960), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n977), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n970), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n984), .B(KEYINPUT126), .ZN(new_n985));
  INV_X1    g560(.A(G8), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n827), .A2(new_n828), .ZN(new_n987));
  AOI21_X1  g562(.A(G1384), .B1(new_n987), .B2(new_n517), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n986), .B1(new_n988), .B2(new_n958), .ZN(new_n989));
  OAI21_X1  g564(.A(G1981), .B1(new_n579), .B2(KEYINPUT110), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n990), .B(KEYINPUT49), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(new_n582), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n992), .A2(G1976), .A3(G288), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n582), .A2(new_n684), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT111), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n989), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(G166), .B2(new_n986), .ZN(new_n998));
  NAND3_X1  g573(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G1384), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n512), .A2(new_n1001), .A3(new_n518), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n954), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT91), .B1(new_n1004), .B2(new_n513), .ZN(new_n1005));
  INV_X1    g580(.A(new_n828), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n517), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1007), .A2(KEYINPUT45), .A3(new_n1001), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1003), .A2(new_n1008), .A3(new_n958), .ZN(new_n1009));
  INV_X1    g584(.A(G1971), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT107), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1009), .A2(KEYINPUT107), .A3(new_n1010), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NOR4_X1   g590(.A1(new_n829), .A2(KEYINPUT108), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT108), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1017), .B1(new_n988), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1002), .A2(KEYINPUT50), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1016), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT109), .B(G2090), .Z(new_n1022));
  NOR3_X1   g597(.A1(new_n1021), .A2(new_n957), .A3(new_n1022), .ZN(new_n1023));
  OAI211_X1 g598(.A(G8), .B(new_n1000), .C1(new_n1015), .C2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n688), .A2(G1976), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n989), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT52), .ZN(new_n1027));
  INV_X1    g602(.A(G1976), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT52), .B1(G288), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1029), .A2(new_n989), .A3(new_n1025), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n992), .A2(new_n989), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1027), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n996), .B1(new_n1024), .B2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n512), .A2(KEYINPUT45), .A3(new_n1001), .A4(new_n518), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n955), .A2(new_n958), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n723), .ZN(new_n1036));
  OR2_X1    g611(.A1(new_n957), .A2(G2084), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1036), .B1(new_n1021), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1038), .A2(G8), .A3(G168), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n988), .A2(new_n1018), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n958), .B1(new_n1002), .B2(KEYINPUT50), .ZN(new_n1042));
  OR2_X1    g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1011), .B1(new_n1043), .B2(new_n1022), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G8), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1000), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1032), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1024), .A2(new_n1040), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT112), .B(KEYINPUT63), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(G8), .B1(new_n1015), .B2(new_n1023), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n1046), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT63), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1039), .A2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1053), .A2(new_n1024), .A3(new_n1048), .A4(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1033), .B1(new_n1051), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1024), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n751), .B1(new_n1021), .B2(new_n957), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1003), .A2(new_n1008), .A3(new_n444), .A4(new_n958), .ZN(new_n1060));
  XOR2_X1   g635(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT119), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1060), .A2(KEYINPUT119), .A3(new_n1061), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1059), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n955), .A2(new_n444), .A3(new_n958), .A4(new_n1034), .ZN(new_n1065));
  OR2_X1    g640(.A1(new_n1065), .A2(KEYINPUT117), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(KEYINPUT117), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1066), .A2(KEYINPUT53), .A3(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(G171), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1058), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1007), .A2(new_n1018), .A3(new_n1001), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1020), .A2(new_n1071), .A3(KEYINPUT108), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n988), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1037), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1035), .A2(new_n723), .ZN(new_n1075));
  OAI21_X1  g650(.A(G8), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n1077));
  NAND2_X1  g652(.A1(G286), .A2(G8), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1078), .B(KEYINPUT116), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT51), .B1(new_n1081), .B2(new_n1079), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1079), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1083), .B1(new_n1038), .B2(G8), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1080), .B(KEYINPUT62), .C1(new_n1082), .C2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1080), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT62), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1077), .B1(new_n1038), .B2(new_n1083), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1093), .A2(KEYINPUT122), .A3(KEYINPUT62), .A4(new_n1080), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1070), .A2(new_n1087), .A3(new_n1090), .A4(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT114), .ZN(new_n1096));
  XOR2_X1   g671(.A(G299), .B(KEYINPUT57), .Z(new_n1097));
  XOR2_X1   g672(.A(KEYINPUT113), .B(G1956), .Z(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT56), .B(G2072), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1003), .A2(new_n1008), .A3(new_n958), .A4(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1097), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n988), .A2(new_n965), .A3(new_n958), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n957), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1103), .B1(new_n1104), .B2(G1348), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1102), .B1(new_n1105), .B2(new_n601), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1099), .A2(new_n1097), .A3(new_n1101), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1096), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G1348), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1110), .B1(new_n1021), .B2(new_n957), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n600), .B1(new_n1111), .B2(new_n1103), .ZN(new_n1112));
  OAI211_X1 g687(.A(KEYINPUT114), .B(new_n1107), .C1(new_n1112), .C2(new_n1102), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1109), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT60), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n600), .B1(new_n1105), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1105), .A2(new_n1115), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1111), .A2(KEYINPUT60), .A3(new_n601), .A4(new_n1103), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT115), .B1(new_n1108), .B2(new_n1102), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT61), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OAI211_X1 g697(.A(KEYINPUT115), .B(KEYINPUT61), .C1(new_n1108), .C2(new_n1102), .ZN(new_n1123));
  OR2_X1    g698(.A1(new_n1009), .A2(G1996), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n988), .A2(new_n958), .ZN(new_n1125));
  XOR2_X1   g700(.A(KEYINPUT58), .B(G1341), .Z(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n558), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n1129));
  OR2_X1    g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1122), .A2(new_n1123), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1114), .B1(new_n1119), .B2(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1059), .B(KEYINPUT120), .ZN(new_n1134));
  XOR2_X1   g709(.A(G171), .B(KEYINPUT54), .Z(new_n1135));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n1136));
  OAI211_X1 g711(.A(KEYINPUT53), .B(new_n444), .C1(new_n957), .C2(new_n1136), .ZN(new_n1137));
  AOI211_X1 g712(.A(new_n1137), .B(new_n956), .C1(new_n1136), .C2(new_n957), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1135), .B1(new_n1138), .B2(new_n1008), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1134), .B(new_n1139), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1058), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1088), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1135), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1057), .B(new_n1095), .C1(new_n1133), .C2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT123), .ZN(new_n1146));
  XNOR2_X1  g721(.A(G290), .B(G1986), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n960), .B1(new_n981), .B2(new_n1147), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1145), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1146), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n985), .B1(new_n1149), .B2(new_n1150), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g726(.A1(G401), .A2(new_n464), .A3(G227), .ZN(new_n1153));
  XNOR2_X1  g727(.A(new_n1153), .B(KEYINPUT127), .ZN(new_n1154));
  AOI211_X1 g728(.A(G229), .B(new_n1154), .C1(new_n946), .C2(new_n945), .ZN(new_n1155));
  NAND2_X1  g729(.A1(new_n871), .A2(new_n875), .ZN(new_n1156));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n1156), .ZN(G225));
  INV_X1    g731(.A(G225), .ZN(G308));
endmodule


