//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 1 0 1 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 1 1 0 1 1 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n206));
  INV_X1    g0006(.A(G116), .ZN(new_n207));
  INV_X1    g0007(.A(G270), .ZN(new_n208));
  OAI21_X1  g0008(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n209), .B(new_n215), .C1(G58), .C2(G232), .ZN(new_n216));
  INV_X1    g0016(.A(G1), .ZN(new_n217));
  INV_X1    g0017(.A(G20), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT65), .ZN(new_n223));
  INV_X1    g0023(.A(G13), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT0), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n218), .A2(KEYINPUT64), .ZN(new_n229));
  INV_X1    g0029(.A(KEYINPUT64), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G20), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  OAI21_X1  g0033(.A(G50), .B1(G58), .B2(G68), .ZN(new_n234));
  NOR3_X1   g0034(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(new_n221), .B2(KEYINPUT1), .ZN(new_n236));
  NAND3_X1  g0036(.A1(new_n223), .A2(new_n228), .A3(new_n236), .ZN(new_n237));
  INV_X1    g0037(.A(new_n237), .ZN(G361));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT2), .ZN(new_n241));
  INV_X1    g0041(.A(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G264), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n208), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(G107), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(new_n207), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n250), .B(new_n253), .Z(G351));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n233), .ZN(new_n256));
  AND2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT7), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n232), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT3), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n264), .A2(new_n218), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT7), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n261), .A2(new_n267), .A3(G68), .ZN(new_n268));
  INV_X1    g0068(.A(G58), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(new_n211), .ZN(new_n270));
  OAI21_X1  g0070(.A(G20), .B1(new_n270), .B2(new_n201), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G20), .A2(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G159), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n268), .A2(KEYINPUT16), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n271), .A2(new_n273), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n232), .A2(new_n259), .A3(KEYINPUT7), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n266), .A2(new_n260), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n276), .B1(new_n279), .B2(G68), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n256), .B(new_n275), .C1(new_n280), .C2(KEYINPUT16), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n255), .A2(new_n233), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n217), .A2(G13), .A3(G20), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n217), .A2(KEYINPUT68), .A3(G20), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT68), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n285), .B1(new_n218), .B2(G1), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n282), .A2(new_n283), .A3(new_n284), .A4(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n269), .A2(KEYINPUT8), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT8), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G58), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT66), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n269), .A2(KEYINPUT66), .A3(KEYINPUT8), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n287), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n283), .B1(new_n292), .B2(new_n293), .ZN(new_n296));
  OAI21_X1  g0096(.A(KEYINPUT73), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n296), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT73), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n298), .B(new_n299), .C1(new_n294), .C2(new_n287), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g0101(.A(G226), .B(G1698), .C1(new_n257), .C2(new_n258), .ZN(new_n302));
  INV_X1    g0102(.A(G1698), .ZN(new_n303));
  OAI211_X1 g0103(.A(G223), .B(new_n303), .C1(new_n257), .C2(new_n258), .ZN(new_n304));
  NAND2_X1  g0104(.A1(G33), .A2(G87), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G41), .ZN(new_n307));
  OAI211_X1 g0107(.A(G1), .B(G13), .C1(new_n263), .C2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n217), .B1(G41), .B2(G45), .ZN(new_n311));
  INV_X1    g0111(.A(G274), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n308), .A2(new_n311), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G232), .ZN(new_n316));
  AND4_X1   g0116(.A1(G179), .A2(new_n310), .A3(new_n314), .A4(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G169), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n313), .B1(new_n306), .B2(new_n309), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n318), .B1(new_n319), .B2(new_n316), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT74), .B1(new_n317), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n310), .A2(new_n314), .A3(new_n316), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G169), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT74), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n319), .A2(G179), .A3(new_n316), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  AOI221_X4 g0126(.A(KEYINPUT18), .B1(new_n281), .B2(new_n301), .C1(new_n321), .C2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT18), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n321), .A2(new_n326), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n281), .A2(new_n301), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n322), .A2(G200), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n319), .A2(G190), .A3(new_n316), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n281), .A2(new_n301), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n335), .A2(KEYINPUT17), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(KEYINPUT17), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AND2_X1   g0138(.A1(new_n332), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(G33), .A2(G97), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT3), .B(G33), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n303), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(G232), .ZN(new_n343));
  OAI221_X1 g0143(.A(new_n340), .B1(new_n342), .B2(new_n242), .C1(new_n303), .C2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n313), .B1(new_n344), .B2(new_n309), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT13), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n315), .A2(G238), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n346), .B1(new_n345), .B2(new_n347), .ZN(new_n350));
  OAI21_X1  g0150(.A(G169), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT14), .ZN(new_n352));
  INV_X1    g0152(.A(new_n350), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n353), .A2(G179), .A3(new_n348), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT72), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT14), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n357), .B(G169), .C1(new_n349), .C2(new_n350), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n353), .A2(KEYINPUT72), .A3(G179), .A4(new_n348), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n352), .A2(new_n356), .A3(new_n358), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n272), .A2(G50), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT67), .ZN(new_n362));
  XNOR2_X1  g0162(.A(KEYINPUT64), .B(G20), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n362), .B1(new_n363), .B2(new_n263), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n230), .A2(G20), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n218), .A2(KEYINPUT64), .ZN(new_n366));
  OAI211_X1 g0166(.A(KEYINPUT67), .B(G33), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G77), .ZN(new_n369));
  OAI221_X1 g0169(.A(new_n361), .B1(new_n218), .B2(G68), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n370), .A2(new_n256), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n371), .A2(KEYINPUT11), .ZN(new_n372));
  INV_X1    g0172(.A(new_n283), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n211), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n374), .B(KEYINPUT12), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n371), .A2(KEYINPUT11), .ZN(new_n376));
  INV_X1    g0176(.A(new_n287), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G68), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n372), .A2(new_n375), .A3(new_n376), .A4(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n360), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G190), .ZN(new_n381));
  NOR3_X1   g0181(.A1(new_n349), .A2(new_n350), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G200), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n383), .B1(new_n353), .B2(new_n348), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n379), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n363), .A2(new_n256), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n369), .B1(new_n287), .B2(new_n387), .ZN(new_n388));
  XOR2_X1   g0188(.A(KEYINPUT15), .B(G87), .Z(new_n389));
  NAND3_X1  g0189(.A1(new_n364), .A2(new_n367), .A3(new_n389), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n288), .A2(new_n290), .ZN(new_n391));
  INV_X1    g0191(.A(new_n272), .ZN(new_n392));
  OR2_X1    g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n388), .B1(new_n394), .B2(new_n256), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT70), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n283), .A2(G77), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n395), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n396), .B1(new_n395), .B2(new_n398), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n259), .A2(G107), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n341), .A2(G1698), .ZN(new_n403));
  OAI221_X1 g0203(.A(new_n402), .B1(new_n403), .B2(new_n212), .C1(G1698), .C2(new_n343), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n309), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n315), .A2(G244), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n314), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G200), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n401), .B(new_n408), .C1(new_n381), .C2(new_n407), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n339), .A2(new_n380), .A3(new_n386), .A4(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n272), .A2(G150), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n203), .A2(G20), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n411), .B(new_n412), .C1(new_n368), .C2(new_n294), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n413), .A2(new_n256), .B1(new_n202), .B2(new_n373), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n377), .A2(G50), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(KEYINPUT71), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(KEYINPUT71), .B1(new_n414), .B2(new_n415), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT9), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n341), .A2(G223), .A3(G1698), .ZN(new_n420));
  INV_X1    g0220(.A(G222), .ZN(new_n421));
  OAI221_X1 g0221(.A(new_n420), .B1(new_n369), .B2(new_n341), .C1(new_n342), .C2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n309), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n315), .A2(G226), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(new_n424), .A3(new_n314), .ZN(new_n425));
  OR2_X1    g0225(.A1(new_n425), .A2(new_n381), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n413), .A2(new_n256), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n373), .A2(new_n202), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(new_n428), .A3(new_n415), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT71), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT9), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n431), .A2(new_n432), .A3(new_n416), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n425), .A2(G200), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n419), .A2(new_n426), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT10), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n431), .A2(new_n416), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n437), .A2(KEYINPUT9), .B1(G200), .B2(new_n425), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT10), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n438), .A2(new_n439), .A3(new_n426), .A4(new_n433), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n436), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G179), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n423), .A2(new_n442), .A3(new_n424), .A4(new_n314), .ZN(new_n443));
  XNOR2_X1  g0243(.A(new_n443), .B(KEYINPUT69), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n425), .A2(new_n318), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(new_n429), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  OR2_X1    g0247(.A1(new_n407), .A2(G179), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n407), .A2(new_n318), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n448), .B(new_n449), .C1(new_n399), .C2(new_n400), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n410), .A2(new_n447), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT75), .ZN(new_n453));
  XNOR2_X1  g0253(.A(new_n452), .B(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n341), .A2(G250), .A3(new_n303), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G294), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n456), .B(new_n457), .C1(new_n403), .C2(new_n214), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n309), .ZN(new_n459));
  INV_X1    g0259(.A(G45), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(G1), .ZN(new_n461));
  AND2_X1   g0261(.A1(KEYINPUT5), .A2(G41), .ZN(new_n462));
  NOR2_X1   g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OR2_X1    g0264(.A1(new_n464), .A2(new_n312), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n464), .A2(new_n308), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G264), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n459), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT84), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n468), .A2(new_n469), .A3(new_n442), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n459), .A2(new_n465), .A3(new_n467), .ZN(new_n471));
  OAI21_X1  g0271(.A(KEYINPUT84), .B1(new_n471), .B2(new_n318), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(G179), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n283), .A2(G107), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT25), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI211_X1 g0277(.A(new_n256), .B(new_n373), .C1(new_n217), .C2(G33), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(G107), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(KEYINPUT23), .B1(new_n218), .B2(G107), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G116), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n482), .B1(G20), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(KEYINPUT23), .A2(G107), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n484), .B1(new_n363), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT82), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT24), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT22), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n229), .A2(new_n231), .B1(new_n264), .B2(new_n265), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n489), .B1(new_n490), .B2(G87), .ZN(new_n491));
  AND4_X1   g0291(.A1(new_n489), .A2(new_n232), .A3(new_n341), .A4(G87), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n486), .B(new_n488), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n487), .A2(KEYINPUT24), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n232), .A2(new_n341), .A3(G87), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT22), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n490), .A2(new_n489), .A3(G87), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n494), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n499), .A2(new_n486), .A3(new_n488), .A4(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n495), .A2(new_n256), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT83), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n495), .A2(KEYINPUT83), .A3(new_n256), .A4(new_n501), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n481), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n475), .A2(new_n476), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n474), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n504), .A2(new_n505), .ZN(new_n510));
  INV_X1    g0310(.A(new_n481), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n471), .A2(G190), .ZN(new_n512));
  AND4_X1   g0312(.A1(new_n508), .A2(new_n510), .A3(new_n511), .A4(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n468), .A2(G200), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n509), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n389), .A2(new_n283), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n364), .A2(G97), .A3(new_n367), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT19), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n518), .A2(KEYINPUT77), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(KEYINPUT77), .B1(new_n518), .B2(new_n519), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n490), .A2(G68), .ZN(new_n522));
  NOR2_X1   g0322(.A1(G97), .A2(G107), .ZN(new_n523));
  INV_X1    g0323(.A(G87), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n340), .A2(new_n519), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n525), .B1(new_n363), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  NOR3_X1   g0328(.A1(new_n520), .A2(new_n521), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n517), .B1(new_n529), .B2(new_n282), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(KEYINPUT78), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n518), .A2(new_n519), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT77), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n528), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n518), .A2(KEYINPUT77), .A3(new_n519), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n256), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT78), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n538), .A2(new_n539), .A3(new_n517), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n531), .A2(new_n540), .B1(G87), .B2(new_n478), .ZN(new_n541));
  INV_X1    g0341(.A(G244), .ZN(new_n542));
  OAI221_X1 g0342(.A(new_n483), .B1(new_n403), .B2(new_n542), .C1(new_n212), .C2(new_n342), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n309), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n308), .B(G250), .C1(G1), .C2(new_n460), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n461), .A2(G274), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n383), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(G190), .B2(new_n547), .ZN(new_n549));
  INV_X1    g0349(.A(new_n389), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n479), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n539), .B1(new_n538), .B2(new_n517), .ZN(new_n553));
  AOI211_X1 g0353(.A(KEYINPUT78), .B(new_n516), .C1(new_n537), .C2(new_n256), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n547), .A2(G179), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n556), .B1(new_n318), .B2(new_n547), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n541), .A2(new_n549), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n466), .A2(G270), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n465), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT79), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n341), .A2(G264), .A3(G1698), .ZN(new_n562));
  INV_X1    g0362(.A(G303), .ZN(new_n563));
  OAI221_X1 g0363(.A(new_n562), .B1(new_n563), .B2(new_n341), .C1(new_n342), .C2(new_n214), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n309), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT79), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n559), .A2(new_n566), .A3(new_n465), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n561), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  OR2_X1    g0368(.A1(new_n568), .A2(new_n442), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n568), .A2(KEYINPUT21), .A3(G169), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n373), .A2(new_n207), .ZN(new_n572));
  XNOR2_X1  g0372(.A(new_n572), .B(KEYINPUT80), .ZN(new_n573));
  NAND2_X1  g0373(.A1(G33), .A2(G283), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n232), .B(new_n574), .C1(G33), .C2(new_n213), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n575), .B(new_n256), .C1(new_n218), .C2(G116), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT20), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n576), .A2(new_n577), .ZN(new_n579));
  OAI221_X1 g0379(.A(new_n573), .B1(new_n207), .B2(new_n479), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n571), .A2(new_n580), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n568), .A2(G169), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n580), .ZN(new_n583));
  XOR2_X1   g0383(.A(KEYINPUT81), .B(KEYINPUT21), .Z(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n580), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n568), .A2(G200), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n586), .B(new_n587), .C1(new_n381), .C2(new_n568), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n581), .A2(new_n585), .A3(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(G244), .B(new_n303), .C1(new_n257), .C2(new_n258), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT4), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n341), .A2(KEYINPUT4), .A3(G244), .A4(new_n303), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n341), .A2(G250), .A3(G1698), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n574), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n309), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n466), .A2(G257), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n596), .A2(new_n465), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT76), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n596), .A2(KEYINPUT76), .A3(new_n465), .A4(new_n597), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n600), .A2(G200), .A3(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n283), .A2(G97), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n279), .A2(G107), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n392), .A2(new_n369), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT6), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n213), .A2(new_n480), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n607), .B1(new_n608), .B2(new_n523), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n480), .A2(KEYINPUT6), .A3(G97), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n604), .B(new_n606), .C1(new_n232), .C2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n603), .B1(new_n612), .B2(new_n256), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n478), .A2(G97), .ZN(new_n614));
  INV_X1    g0414(.A(new_n598), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G190), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n602), .A2(new_n613), .A3(new_n614), .A4(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n613), .A2(new_n614), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n598), .A2(new_n318), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n615), .A2(new_n442), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n515), .A2(new_n558), .A3(new_n589), .A4(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n455), .A2(new_n623), .ZN(G372));
  INV_X1    g0424(.A(new_n446), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n386), .A2(new_n338), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n451), .B1(new_n360), .B2(new_n379), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n323), .A2(new_n325), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT18), .B1(new_n330), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n330), .A2(new_n628), .A3(KEYINPUT18), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  OAI22_X1  g0431(.A1(new_n626), .A2(new_n627), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n625), .B1(new_n632), .B2(new_n441), .ZN(new_n633));
  AOI211_X1 g0433(.A(new_n507), .B(new_n481), .C1(new_n504), .C2(new_n505), .ZN(new_n634));
  OAI21_X1  g0434(.A(KEYINPUT85), .B1(new_n634), .B2(new_n474), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n571), .A2(new_n580), .B1(new_n583), .B2(new_n584), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n510), .A2(new_n508), .A3(new_n511), .ZN(new_n637));
  INV_X1    g0437(.A(new_n474), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT85), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n635), .A2(new_n636), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n555), .A2(new_n557), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n478), .A2(G87), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n643), .B(new_n549), .C1(new_n553), .C2(new_n554), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n506), .A2(new_n508), .A3(new_n514), .A4(new_n512), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n642), .A2(new_n622), .A3(new_n644), .A4(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT86), .B1(new_n641), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n642), .ZN(new_n648));
  INV_X1    g0448(.A(new_n621), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n551), .B1(new_n531), .B2(new_n540), .ZN(new_n650));
  INV_X1    g0450(.A(new_n557), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n644), .B(new_n649), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT26), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n642), .A2(KEYINPUT26), .A3(new_n644), .A4(new_n649), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n648), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n642), .A2(new_n644), .A3(new_n622), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n635), .A2(new_n636), .A3(new_n640), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT86), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n657), .A2(new_n658), .A3(new_n659), .A4(new_n645), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n647), .A2(new_n656), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n633), .B1(new_n455), .B2(new_n662), .ZN(G369));
  NAND2_X1  g0463(.A1(new_n581), .A2(new_n585), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n363), .A2(new_n224), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n217), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G213), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(G343), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n586), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n664), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n581), .A2(new_n585), .A3(new_n588), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n674), .B1(new_n675), .B2(new_n673), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(G330), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n515), .B1(new_n634), .B2(new_n672), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n637), .A2(new_n638), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n679), .B1(new_n680), .B2(new_n672), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n635), .A2(new_n640), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n672), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n664), .A2(new_n672), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n515), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n682), .A2(new_n684), .A3(new_n687), .ZN(G399));
  NOR2_X1   g0488(.A1(new_n225), .A2(G41), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n525), .A2(G116), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(G1), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n234), .B2(new_n690), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n661), .A2(new_n672), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT29), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT88), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n657), .B(new_n645), .C1(new_n664), .C2(new_n509), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n671), .B1(new_n700), .B2(new_n656), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT29), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n695), .A2(KEYINPUT88), .A3(new_n696), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n699), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n568), .A2(new_n442), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n547), .A2(new_n468), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n705), .A2(new_n706), .A3(new_n596), .A4(new_n597), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n615), .A2(new_n471), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(new_n442), .A3(new_n568), .A4(new_n547), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n707), .A2(new_n708), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n709), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n671), .ZN(new_n714));
  OAI211_X1 g0514(.A(KEYINPUT31), .B(new_n714), .C1(new_n623), .C2(new_n671), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(KEYINPUT31), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n715), .A2(G330), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(KEYINPUT87), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT87), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n715), .A2(new_n720), .A3(G330), .A4(new_n717), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n704), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n694), .B1(new_n723), .B2(G1), .ZN(G364));
  AOI21_X1  g0524(.A(new_n217), .B1(new_n665), .B2(G45), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n690), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT89), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n678), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(G330), .B2(new_n676), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n250), .A2(G45), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n225), .A2(new_n341), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n730), .B(new_n731), .C1(G45), .C2(new_n234), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n226), .A2(new_n341), .ZN(new_n733));
  XNOR2_X1  g0533(.A(G355), .B(KEYINPUT90), .ZN(new_n734));
  OAI221_X1 g0534(.A(new_n732), .B1(G116), .B2(new_n226), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n233), .B1(G20), .B2(new_n318), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n736), .A2(KEYINPUT91), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(KEYINPUT91), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G13), .A2(G33), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G20), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n735), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n727), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n232), .A2(new_n442), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(G190), .A3(new_n383), .ZN(new_n747));
  INV_X1    g0547(.A(G322), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR4_X1   g0549(.A1(new_n232), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n341), .B1(new_n750), .B2(G329), .ZN(new_n751));
  INV_X1    g0551(.A(G294), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n381), .A2(G179), .A3(G200), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n232), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n751), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n746), .A2(new_n381), .A3(new_n383), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT92), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n749), .B(new_n755), .C1(new_n760), .C2(G311), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n383), .A2(G179), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n363), .A2(new_n381), .A3(new_n762), .ZN(new_n763));
  XOR2_X1   g0563(.A(new_n763), .B(KEYINPUT93), .Z(new_n764));
  INV_X1    g0564(.A(G283), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n746), .A2(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G190), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  XOR2_X1   g0568(.A(KEYINPUT33), .B(G317), .Z(new_n769));
  OAI22_X1  g0569(.A1(new_n764), .A2(new_n765), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n766), .A2(new_n381), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n770), .B1(G326), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n762), .A2(G20), .A3(G190), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n761), .B(new_n772), .C1(new_n563), .C2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n524), .ZN(new_n775));
  INV_X1    g0575(.A(new_n750), .ZN(new_n776));
  INV_X1    g0576(.A(G159), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT32), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n778), .A2(new_n779), .B1(new_n269), .B2(new_n747), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n775), .B(new_n780), .C1(G77), .C2(new_n760), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n764), .A2(new_n480), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(G68), .B2(new_n767), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n754), .A2(new_n213), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n259), .B(new_n784), .C1(new_n778), .C2(new_n779), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n781), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n771), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n202), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n774), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n745), .B1(new_n789), .B2(new_n739), .ZN(new_n790));
  INV_X1    g0590(.A(new_n742), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n744), .B(new_n790), .C1(new_n676), .C2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n729), .A2(new_n792), .ZN(G396));
  OAI21_X1  g0593(.A(new_n671), .B1(new_n399), .B2(new_n400), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n451), .A2(KEYINPUT96), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT96), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n450), .A2(new_n796), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n409), .B(new_n794), .C1(new_n795), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n451), .A2(new_n671), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n695), .A2(new_n801), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n795), .A2(new_n797), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n803), .A2(new_n409), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n661), .A2(new_n672), .A3(new_n804), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n722), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n727), .B1(new_n808), .B2(KEYINPUT97), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n806), .A2(new_n807), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n809), .B(new_n810), .C1(KEYINPUT97), .C2(new_n808), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n739), .A2(new_n740), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n745), .B1(new_n369), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT94), .ZN(new_n814));
  INV_X1    g0614(.A(G137), .ZN(new_n815));
  INV_X1    g0615(.A(G150), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n815), .A2(new_n787), .B1(new_n768), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(G159), .B2(new_n760), .ZN(new_n818));
  INV_X1    g0618(.A(G143), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n818), .B1(new_n819), .B2(new_n747), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT34), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n341), .B1(new_n754), .B2(new_n269), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n764), .A2(new_n211), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n822), .B(new_n823), .C1(G132), .C2(new_n750), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n821), .B(new_n824), .C1(new_n202), .C2(new_n773), .ZN(new_n825));
  INV_X1    g0625(.A(G311), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n776), .A2(new_n826), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n784), .B(new_n827), .C1(new_n760), .C2(G116), .ZN(new_n828));
  INV_X1    g0628(.A(new_n764), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(G87), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G283), .A2(new_n767), .B1(new_n771), .B2(G303), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n259), .B1(new_n773), .B2(new_n480), .ZN(new_n832));
  INV_X1    g0632(.A(new_n747), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(new_n833), .B2(G294), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n828), .A2(new_n830), .A3(new_n831), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n825), .A2(new_n835), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT95), .Z(new_n837));
  INV_X1    g0637(.A(new_n739), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n814), .B1(new_n741), .B2(new_n800), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n811), .A2(new_n839), .ZN(G384));
  INV_X1    g0640(.A(G330), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT31), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n642), .A2(new_n644), .A3(new_n622), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n680), .A2(new_n645), .ZN(new_n844));
  NOR3_X1   g0644(.A1(new_n843), .A2(new_n844), .A3(new_n675), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n842), .B1(new_n845), .B2(new_n672), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n716), .B1(new_n846), .B2(new_n714), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n454), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n379), .A2(new_n671), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n380), .A2(new_n386), .A3(new_n849), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n379), .B(new_n671), .C1(new_n360), .C2(new_n385), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n850), .A2(new_n851), .B1(new_n798), .B2(new_n799), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n715), .A2(new_n717), .A3(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT38), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n275), .A2(new_n256), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT16), .B1(new_n268), .B2(new_n274), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n298), .B1(new_n294), .B2(new_n287), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n669), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n332), .B2(new_n338), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n321), .A2(new_n326), .B1(new_n281), .B2(new_n301), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT37), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n335), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n669), .B1(new_n281), .B2(new_n301), .ZN(new_n864));
  NOR3_X1   g0664(.A1(new_n861), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n857), .B1(new_n628), .B2(new_n858), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n862), .B1(new_n866), .B2(new_n335), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n854), .B1(new_n860), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n329), .A2(new_n330), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT18), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n861), .A2(new_n328), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n338), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n859), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OR2_X1    g0675(.A1(new_n865), .A2(new_n867), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n875), .A2(new_n876), .A3(KEYINPUT38), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT99), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n869), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT40), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n875), .A2(new_n876), .A3(KEYINPUT99), .A4(KEYINPUT38), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n330), .A2(new_n628), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n328), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n336), .A2(new_n337), .B1(new_n884), .B2(new_n630), .ZN(new_n885));
  INV_X1    g0685(.A(new_n864), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT102), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n281), .A2(new_n301), .A3(new_n334), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n888), .A2(new_n333), .B1(new_n330), .B2(new_n628), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n862), .B1(new_n889), .B2(new_n886), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT101), .B1(new_n890), .B2(new_n865), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n883), .A2(new_n335), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT37), .B1(new_n892), .B2(new_n864), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT101), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n870), .A2(new_n886), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n893), .B(new_n894), .C1(new_n863), .C2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n337), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n335), .A2(KEYINPUT17), .ZN(new_n898));
  OAI22_X1  g0698(.A1(new_n897), .A2(new_n898), .B1(new_n631), .B2(new_n629), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT102), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n899), .A2(new_n900), .A3(new_n864), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n887), .A2(new_n891), .A3(new_n896), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n854), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n877), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n904), .A2(new_n715), .A3(new_n717), .A4(new_n852), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n853), .A2(new_n882), .B1(new_n905), .B2(KEYINPUT40), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n841), .B1(new_n848), .B2(new_n906), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n907), .B(KEYINPUT104), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n848), .B2(new_n906), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n803), .A2(new_n671), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n805), .A2(new_n911), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n850), .A2(new_n851), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n879), .A2(new_n881), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n912), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n884), .A2(new_n630), .A3(new_n669), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n380), .A2(new_n671), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n879), .A2(KEYINPUT39), .A3(new_n881), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT100), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT39), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n903), .A2(new_n924), .A3(new_n877), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n921), .B1(new_n920), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n916), .B(new_n917), .C1(new_n919), .C2(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n909), .B(new_n928), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n699), .A2(new_n454), .A3(new_n702), .A4(new_n703), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n633), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT103), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n929), .B(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n217), .B2(new_n665), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT35), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n233), .B(new_n232), .C1(new_n611), .C2(new_n935), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n936), .B(G116), .C1(new_n935), .C2(new_n611), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT36), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT98), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n211), .B2(G50), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n202), .A2(KEYINPUT98), .A3(G68), .ZN(new_n941));
  OAI21_X1  g0741(.A(G77), .B1(new_n269), .B2(new_n211), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n940), .B(new_n941), .C1(new_n942), .C2(new_n234), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n943), .A2(G1), .A3(new_n224), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n934), .A2(new_n938), .A3(new_n944), .ZN(G367));
  NAND2_X1  g0745(.A1(new_n618), .A2(new_n671), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n622), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n649), .A2(new_n671), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n687), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT42), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n621), .B1(new_n947), .B2(new_n680), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT106), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n672), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n541), .A2(new_n672), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n648), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n558), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n958), .B1(new_n959), .B2(new_n957), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(KEYINPUT105), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT105), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n958), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n956), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n956), .A2(new_n965), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT107), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NOR3_X1   g0770(.A1(new_n956), .A2(KEYINPUT107), .A3(new_n965), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n967), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n682), .A2(new_n950), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n972), .B(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n687), .A2(new_n684), .A3(new_n949), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT45), .Z(new_n976));
  AOI21_X1  g0776(.A(new_n949), .B1(new_n687), .B2(new_n684), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT44), .ZN(new_n978));
  AND3_X1   g0778(.A1(new_n976), .A2(new_n682), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n682), .B1(new_n976), .B2(new_n978), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n687), .B1(new_n681), .B2(new_n686), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(new_n677), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n723), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n689), .B(KEYINPUT41), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n725), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n974), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n961), .A2(new_n742), .A3(new_n963), .ZN(new_n990));
  INV_X1    g0790(.A(new_n731), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n743), .B1(new_n226), .B2(new_n550), .C1(new_n246), .C2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n773), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(G116), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT46), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n213), .B2(new_n763), .C1(new_n480), .C2(new_n754), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n752), .A2(new_n768), .B1(new_n787), .B2(new_n826), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n259), .B1(new_n747), .B2(new_n563), .ZN(new_n998));
  NOR3_X1   g0798(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n760), .ZN(new_n1000));
  INV_X1    g0800(.A(G317), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n999), .B1(new_n765), .B2(new_n1000), .C1(new_n1001), .C2(new_n776), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n819), .A2(new_n787), .B1(new_n768), .B2(new_n777), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n747), .A2(new_n816), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n211), .A2(new_n754), .B1(new_n763), .B2(new_n369), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n341), .B1(new_n776), .B2(new_n815), .ZN(new_n1006));
  NOR4_X1   g0806(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1007), .B1(new_n202), .B2(new_n1000), .C1(new_n269), .C2(new_n773), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1002), .A2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n1010));
  XNOR2_X1  g0810(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n745), .B1(new_n1011), .B2(new_n739), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n990), .A2(new_n992), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n989), .A2(new_n1013), .ZN(G387));
  INV_X1    g0814(.A(new_n984), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n723), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n723), .A2(new_n1015), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1016), .A2(new_n689), .A3(new_n1017), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(G311), .A2(new_n767), .B1(new_n771), .B2(G322), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n1001), .B2(new_n747), .C1(new_n1000), .C2(new_n563), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1021), .A2(KEYINPUT48), .B1(G294), .B2(new_n993), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n765), .B2(new_n754), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT111), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1021), .A2(KEYINPUT48), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AND2_X1   g0826(.A1(new_n1026), .A2(KEYINPUT49), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n763), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n341), .B1(new_n1028), .B2(G116), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n1026), .B2(KEYINPUT49), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n750), .A2(G326), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n1027), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n764), .A2(new_n213), .B1(new_n768), .B2(new_n294), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n389), .B1(new_n232), .B2(new_n753), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n369), .B2(new_n773), .C1(new_n776), .C2(new_n816), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(G68), .B2(new_n760), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n259), .B1(new_n833), .B2(G50), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n1033), .B(new_n1038), .C1(G159), .C2(new_n771), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n739), .B1(new_n1032), .B2(new_n1039), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n681), .A2(new_n791), .ZN(new_n1041));
  AND3_X1   g0841(.A1(new_n1040), .A2(new_n727), .A3(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n391), .A2(G50), .ZN(new_n1043));
  XOR2_X1   g0843(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n1044));
  OR2_X1    g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n691), .B(KEYINPUT109), .ZN(new_n1046));
  AOI21_X1  g0846(.A(G45), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(G68), .A2(G77), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n731), .B(new_n1049), .C1(new_n243), .C2(new_n460), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(G107), .B2(new_n226), .C1(new_n691), .C2(new_n733), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n743), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n1042), .A2(new_n1052), .B1(new_n988), .B2(new_n1015), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1018), .A2(new_n1053), .ZN(G393));
  NAND3_X1  g0854(.A1(new_n976), .A2(new_n682), .A3(new_n978), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1055), .A2(KEYINPUT112), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n981), .B2(KEYINPUT112), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1017), .A2(new_n1057), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1058), .B(new_n689), .C1(new_n1017), .C2(new_n982), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1057), .A2(new_n725), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n754), .A2(new_n369), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1000), .A2(new_n391), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n259), .B1(new_n993), .B2(G68), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n830), .B(new_n1063), .C1(new_n819), .C2(new_n776), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT113), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1061), .B(new_n1062), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n767), .A2(G50), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n787), .A2(new_n816), .B1(new_n777), .B2(new_n747), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT51), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .A4(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G317), .A2(new_n771), .B1(new_n833), .B2(G311), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT114), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n1073), .A2(KEYINPUT52), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(KEYINPUT52), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1000), .A2(new_n752), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n768), .A2(new_n563), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n259), .B1(new_n207), .B2(new_n754), .C1(new_n776), .C2(new_n748), .ZN(new_n1078));
  NOR4_X1   g0878(.A1(new_n1076), .A2(new_n782), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1074), .A2(new_n1075), .A3(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n773), .A2(new_n765), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1071), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n745), .B1(new_n1082), .B2(new_n739), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n950), .A2(new_n742), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n743), .B1(new_n213), .B2(new_n226), .C1(new_n253), .C2(new_n991), .ZN(new_n1085));
  AND3_X1   g0885(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1060), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1059), .A2(new_n1087), .ZN(G390));
  AOI21_X1  g0888(.A(new_n910), .B1(new_n701), .B2(new_n804), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n919), .B(new_n904), .C1(new_n1089), .C2(new_n913), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n918), .B1(new_n912), .B2(new_n914), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n920), .A2(new_n925), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(KEYINPUT100), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n922), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1090), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n719), .A2(new_n721), .A3(new_n852), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT115), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n719), .A2(KEYINPUT115), .A3(new_n721), .A4(new_n852), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1095), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n913), .B1(new_n805), .B2(new_n911), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n927), .B1(new_n1102), .B2(new_n918), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n718), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1103), .A2(new_n1090), .B1(new_n1104), .B2(new_n852), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n454), .A2(G330), .A3(new_n847), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n930), .A2(new_n633), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(KEYINPUT116), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT116), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n930), .A2(new_n1110), .A3(new_n633), .A4(new_n1107), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n914), .B1(new_n1104), .B2(new_n800), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n719), .A2(new_n721), .A3(new_n800), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n913), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1104), .A2(new_n852), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1114), .A2(new_n1089), .B1(new_n1118), .B2(new_n912), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1106), .B1(new_n1112), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1113), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1100), .A2(new_n1089), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1118), .A2(new_n912), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1095), .A2(new_n1117), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1103), .A2(new_n1090), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1124), .A2(new_n1127), .A3(new_n1111), .A4(new_n1109), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1120), .A2(new_n689), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n927), .A2(new_n740), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n812), .A2(new_n294), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n760), .A2(G97), .B1(G107), .B2(new_n767), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT118), .ZN(new_n1133));
  OR2_X1    g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1061), .B(new_n823), .C1(G283), .C2(new_n771), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n259), .B1(new_n776), .B2(new_n752), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n775), .B(new_n1137), .C1(new_n833), .C2(G116), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n750), .A2(G125), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n777), .B2(new_n754), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n833), .B2(G132), .ZN(new_n1142));
  XOR2_X1   g0942(.A(KEYINPUT54), .B(G143), .Z(new_n1143));
  NAND2_X1  g0943(.A1(new_n760), .A2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n773), .A2(new_n816), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT53), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G128), .A2(new_n771), .B1(new_n767), .B2(G137), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1142), .A2(new_n1144), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n341), .B1(new_n763), .B2(new_n202), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT117), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1139), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT119), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n745), .B1(new_n1152), .B2(new_n739), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1130), .A2(new_n1131), .A3(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n1106), .B2(new_n725), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1129), .A2(new_n1156), .ZN(G378));
  AOI22_X1  g0957(.A1(new_n760), .A2(G137), .B1(G132), .B2(new_n767), .ZN(new_n1158));
  XOR2_X1   g0958(.A(new_n1158), .B(KEYINPUT120), .Z(new_n1159));
  NAND2_X1  g0959(.A1(new_n993), .A2(new_n1143), .ZN(new_n1160));
  INV_X1    g0960(.A(G128), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n747), .A2(new_n1161), .B1(new_n816), .B2(new_n754), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(G125), .B2(new_n771), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1159), .A2(new_n1160), .A3(new_n1163), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n1164), .B(KEYINPUT59), .Z(new_n1165));
  AOI21_X1  g0965(.A(G41), .B1(new_n750), .B2(G124), .ZN(new_n1166));
  AOI21_X1  g0966(.A(G33), .B1(new_n1028), .B2(G159), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n763), .A2(new_n269), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G283), .B2(new_n750), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n211), .B2(new_n754), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n768), .A2(new_n213), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n307), .B(new_n259), .C1(new_n773), .C2(new_n369), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n747), .A2(new_n480), .ZN(new_n1174));
  NOR4_X1   g0974(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1175), .B1(new_n207), .B2(new_n787), .C1(new_n550), .C2(new_n1000), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT58), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n202), .B1(new_n257), .B2(G41), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1168), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT121), .Z(new_n1180));
  AOI21_X1  g0980(.A(new_n745), .B1(new_n1180), .B2(new_n739), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n812), .A2(new_n202), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n437), .A2(new_n669), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n447), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT55), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1183), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n441), .A2(new_n446), .A3(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1184), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1186), .B1(new_n441), .B2(new_n446), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n625), .B(new_n1183), .C1(new_n436), .C2(new_n440), .ZN(new_n1190));
  OAI21_X1  g0990(.A(KEYINPUT55), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1188), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT56), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1188), .A2(new_n1191), .A3(KEYINPUT56), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1181), .B(new_n1182), .C1(new_n741), .C2(new_n1196), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n1197), .A2(KEYINPUT122), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(KEYINPUT122), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1188), .A2(new_n1191), .A3(KEYINPUT56), .ZN(new_n1200));
  AOI21_X1  g1000(.A(KEYINPUT56), .B1(new_n1188), .B2(new_n1191), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NOR3_X1   g1002(.A1(new_n906), .A2(new_n1202), .A3(new_n841), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n905), .A2(KEYINPUT40), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n847), .A2(new_n852), .A3(new_n882), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1196), .B1(new_n1206), .B2(G330), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n928), .B1(new_n1203), .B2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1202), .B1(new_n906), .B2(new_n841), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1094), .A2(new_n918), .B1(new_n1102), .B2(new_n915), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1206), .A2(G330), .A3(new_n1196), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1209), .A2(new_n1210), .A3(new_n917), .A4(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1208), .A2(new_n1212), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1198), .A2(new_n1199), .B1(new_n988), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1112), .B1(new_n1127), .B2(new_n1124), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1208), .A2(new_n1212), .A3(KEYINPUT123), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT123), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n928), .B(new_n1217), .C1(new_n1203), .C2(new_n1207), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1216), .A2(KEYINPUT57), .A3(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n689), .B1(new_n1215), .B2(new_n1219), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1111), .B(new_n1109), .C1(new_n1106), .C2(new_n1119), .ZN(new_n1221));
  AOI21_X1  g1021(.A(KEYINPUT57), .B1(new_n1221), .B2(new_n1213), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1214), .B1(new_n1220), .B2(new_n1222), .ZN(G375));
  NAND2_X1  g1023(.A1(new_n1112), .A2(new_n1119), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1124), .A2(new_n1111), .A3(new_n1109), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1224), .A2(new_n1225), .A3(new_n986), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n913), .A2(new_n740), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1034), .B1(new_n563), .B2(new_n776), .C1(new_n1000), .C2(new_n480), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n764), .A2(new_n369), .B1(new_n768), .B2(new_n207), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n259), .B1(new_n213), .B2(new_n773), .C1(new_n747), .C2(new_n765), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n752), .B2(new_n787), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n771), .A2(G132), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1169), .B(new_n1233), .C1(new_n767), .C2(new_n1143), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n993), .A2(G159), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n1235), .B1(new_n202), .B2(new_n754), .C1(new_n776), .C2(new_n1161), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(G137), .B2(new_n833), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n760), .A2(G150), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1234), .A2(new_n341), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n838), .B1(new_n1232), .B2(new_n1239), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n745), .B(new_n1240), .C1(new_n211), .C2(new_n812), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT124), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1124), .A2(new_n988), .B1(new_n1227), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1226), .A2(new_n1243), .ZN(G381));
  NAND4_X1  g1044(.A1(new_n1018), .A2(new_n792), .A3(new_n729), .A4(new_n1053), .ZN(new_n1245));
  OR3_X1    g1045(.A1(G387), .A2(G384), .A3(new_n1245), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1216), .A2(KEYINPUT57), .A3(new_n1218), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n690), .B1(new_n1247), .B2(new_n1221), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT57), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1213), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1249), .B1(new_n1215), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1112), .A2(new_n1119), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n690), .B1(new_n1253), .B2(new_n1127), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1155), .B1(new_n1254), .B2(new_n1120), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1252), .A2(new_n1255), .A3(new_n1214), .ZN(new_n1256));
  OR4_X1    g1056(.A1(G390), .A2(new_n1246), .A3(new_n1256), .A4(G381), .ZN(G407));
  OAI211_X1 g1057(.A(G407), .B(G213), .C1(G343), .C2(new_n1256), .ZN(G409));
  AOI21_X1  g1058(.A(new_n1124), .B1(new_n1111), .B2(new_n1109), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n689), .B1(new_n1259), .B2(KEYINPUT60), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1112), .A2(KEYINPUT60), .A3(new_n1119), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1225), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1243), .B1(new_n1260), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(G384), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT60), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1224), .A2(new_n1266), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1267), .A2(new_n689), .A3(new_n1225), .A4(new_n1261), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1268), .A2(G384), .A3(new_n1243), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1265), .A2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1255), .B1(new_n1252), .B2(new_n1214), .ZN(new_n1271));
  INV_X1    g1071(.A(G213), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1272), .A2(G343), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1129), .A2(new_n1156), .A3(new_n1197), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1221), .A2(new_n986), .A3(new_n1213), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1216), .A2(new_n988), .A3(new_n1218), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1274), .B1(new_n1275), .B2(new_n1278), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1270), .A2(new_n1271), .A3(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT62), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1268), .A2(G384), .A3(new_n1243), .ZN(new_n1283));
  AOI21_X1  g1083(.A(G384), .B1(new_n1268), .B2(new_n1243), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(G375), .A2(G378), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1129), .A2(new_n1156), .A3(new_n1197), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1277), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1112), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1250), .B1(new_n1128), .B2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1288), .B1(new_n1290), .B2(new_n986), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1273), .B1(new_n1287), .B2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1285), .A2(new_n1286), .A3(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(KEYINPUT62), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT61), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1292), .A2(new_n1286), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1273), .A2(G2897), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1265), .A2(new_n1269), .A3(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1297), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1299), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1296), .A2(new_n1298), .A3(new_n1300), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1282), .A2(new_n1294), .A3(new_n1295), .A4(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT126), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(G393), .A2(G396), .ZN(new_n1304));
  AND2_X1   g1104(.A1(new_n1304), .A2(new_n1245), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n989), .A2(G390), .A3(new_n1013), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n973), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(new_n972), .B(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n988), .B1(new_n985), .B2(new_n986), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1013), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1087), .B(new_n1059), .C1(new_n1310), .C2(new_n1311), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1305), .A2(new_n1306), .A3(new_n1312), .ZN(new_n1313));
  AOI22_X1  g1113(.A1(new_n1312), .A2(new_n1306), .B1(new_n1245), .B2(new_n1304), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1303), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1312), .A2(new_n1306), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1305), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1305), .A2(new_n1312), .A3(new_n1306), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1318), .A2(KEYINPUT126), .A3(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1315), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1302), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1300), .A2(new_n1298), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1271), .A2(new_n1279), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1293), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(KEYINPUT63), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1318), .A2(new_n1295), .A3(new_n1319), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT63), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1327), .B1(new_n1293), .B2(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(KEYINPUT125), .B1(new_n1326), .B2(new_n1329), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1328), .B1(new_n1301), .B2(new_n1293), .ZN(new_n1331));
  NOR3_X1   g1131(.A1(new_n1313), .A2(new_n1314), .A3(KEYINPUT61), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1332), .B1(new_n1280), .B2(KEYINPUT63), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT125), .ZN(new_n1334));
  NOR3_X1   g1134(.A1(new_n1331), .A2(new_n1333), .A3(new_n1334), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1322), .B1(new_n1330), .B2(new_n1335), .ZN(G405));
  NAND3_X1  g1136(.A1(new_n1285), .A2(new_n1256), .A3(new_n1286), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1256), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1270), .B1(new_n1338), .B2(new_n1271), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1321), .A2(new_n1337), .A3(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(KEYINPUT127), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1339), .A2(new_n1337), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1342), .A2(new_n1320), .A3(new_n1315), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT127), .ZN(new_n1344));
  NAND4_X1  g1144(.A1(new_n1321), .A2(new_n1344), .A3(new_n1337), .A4(new_n1339), .ZN(new_n1345));
  AND3_X1   g1145(.A1(new_n1341), .A2(new_n1343), .A3(new_n1345), .ZN(G402));
endmodule


