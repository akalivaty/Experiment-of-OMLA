

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U552 ( .A1(G1384), .A2(n683), .ZN(n684) );
  NOR2_X2 U553 ( .A1(G2104), .A2(n529), .ZN(n516) );
  INV_X1 U554 ( .A(KEYINPUT26), .ZN(n686) );
  INV_X1 U555 ( .A(KEYINPUT64), .ZN(n692) );
  NOR2_X1 U556 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U557 ( .A1(G651), .A2(n649), .ZN(n644) );
  BUF_X1 U558 ( .A(n691), .Z(n937) );
  NOR2_X1 U559 ( .A1(G543), .A2(G651), .ZN(n637) );
  NAND2_X1 U560 ( .A1(n637), .A2(G89), .ZN(n517) );
  XNOR2_X1 U561 ( .A(n517), .B(KEYINPUT4), .ZN(n519) );
  XOR2_X1 U562 ( .A(G543), .B(KEYINPUT0), .Z(n649) );
  XNOR2_X1 U563 ( .A(KEYINPUT65), .B(G651), .ZN(n521) );
  NOR2_X1 U564 ( .A1(n649), .A2(n521), .ZN(n634) );
  NAND2_X1 U565 ( .A1(G76), .A2(n634), .ZN(n518) );
  NAND2_X1 U566 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U567 ( .A(n520), .B(KEYINPUT5), .ZN(n527) );
  NAND2_X1 U568 ( .A1(G51), .A2(n644), .ZN(n524) );
  NOR2_X1 U569 ( .A1(n521), .A2(G543), .ZN(n522) );
  XOR2_X1 U570 ( .A(KEYINPUT1), .B(n522), .Z(n648) );
  NAND2_X1 U571 ( .A1(G63), .A2(n648), .ZN(n523) );
  NAND2_X1 U572 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U573 ( .A(KEYINPUT6), .B(n525), .Z(n526) );
  NAND2_X1 U574 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U575 ( .A(n528), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U576 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U577 ( .A(G2105), .ZN(n529) );
  NAND2_X1 U578 ( .A1(n516), .A2(G125), .ZN(n532) );
  AND2_X1 U579 ( .A1(n529), .A2(G2104), .ZN(n569) );
  NAND2_X1 U580 ( .A1(G101), .A2(n569), .ZN(n530) );
  XOR2_X1 U581 ( .A(n530), .B(KEYINPUT23), .Z(n531) );
  NAND2_X1 U582 ( .A1(n532), .A2(n531), .ZN(n537) );
  NOR2_X1 U583 ( .A1(G2104), .A2(G2105), .ZN(n533) );
  XOR2_X2 U584 ( .A(KEYINPUT17), .B(n533), .Z(n864) );
  NAND2_X1 U585 ( .A1(G137), .A2(n864), .ZN(n535) );
  AND2_X1 U586 ( .A1(G2104), .A2(G2105), .ZN(n861) );
  NAND2_X1 U587 ( .A1(G113), .A2(n861), .ZN(n534) );
  NAND2_X1 U588 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X1 U589 ( .A1(n537), .A2(n536), .ZN(G160) );
  NAND2_X1 U590 ( .A1(G47), .A2(n644), .ZN(n539) );
  NAND2_X1 U591 ( .A1(G85), .A2(n637), .ZN(n538) );
  NAND2_X1 U592 ( .A1(n539), .A2(n538), .ZN(n543) );
  NAND2_X1 U593 ( .A1(G72), .A2(n634), .ZN(n541) );
  NAND2_X1 U594 ( .A1(G60), .A2(n648), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n541), .A2(n540), .ZN(n542) );
  OR2_X1 U596 ( .A1(n543), .A2(n542), .ZN(G290) );
  XOR2_X1 U597 ( .A(G2435), .B(G2454), .Z(n545) );
  XNOR2_X1 U598 ( .A(KEYINPUT105), .B(G2438), .ZN(n544) );
  XNOR2_X1 U599 ( .A(n545), .B(n544), .ZN(n552) );
  XOR2_X1 U600 ( .A(G2446), .B(G2430), .Z(n547) );
  XNOR2_X1 U601 ( .A(G2451), .B(G2443), .ZN(n546) );
  XNOR2_X1 U602 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U603 ( .A(n548), .B(G2427), .Z(n550) );
  XNOR2_X1 U604 ( .A(G1348), .B(G1341), .ZN(n549) );
  XNOR2_X1 U605 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U606 ( .A(n552), .B(n551), .ZN(n553) );
  AND2_X1 U607 ( .A1(n553), .A2(G14), .ZN(G401) );
  NAND2_X1 U608 ( .A1(G138), .A2(n864), .ZN(n558) );
  AND2_X1 U609 ( .A1(G102), .A2(n569), .ZN(n557) );
  NAND2_X1 U610 ( .A1(G126), .A2(n516), .ZN(n555) );
  NAND2_X1 U611 ( .A1(G114), .A2(n861), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U613 ( .A1(n557), .A2(n556), .ZN(n683) );
  AND2_X1 U614 ( .A1(n558), .A2(n683), .ZN(G164) );
  XNOR2_X1 U615 ( .A(KEYINPUT67), .B(KEYINPUT9), .ZN(n562) );
  NAND2_X1 U616 ( .A1(n637), .A2(G90), .ZN(n560) );
  NAND2_X1 U617 ( .A1(G77), .A2(n634), .ZN(n559) );
  NAND2_X1 U618 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U619 ( .A(n562), .B(n561), .ZN(n567) );
  NAND2_X1 U620 ( .A1(n644), .A2(G52), .ZN(n563) );
  XNOR2_X1 U621 ( .A(n563), .B(KEYINPUT66), .ZN(n565) );
  NAND2_X1 U622 ( .A1(G64), .A2(n648), .ZN(n564) );
  NAND2_X1 U623 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U624 ( .A1(n567), .A2(n566), .ZN(G171) );
  AND2_X1 U625 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U626 ( .A1(G123), .A2(n516), .ZN(n568) );
  XNOR2_X1 U627 ( .A(n568), .B(KEYINPUT18), .ZN(n577) );
  INV_X1 U628 ( .A(n569), .ZN(n570) );
  INV_X1 U629 ( .A(n570), .ZN(n866) );
  NAND2_X1 U630 ( .A1(G99), .A2(n866), .ZN(n572) );
  NAND2_X1 U631 ( .A1(G111), .A2(n861), .ZN(n571) );
  NAND2_X1 U632 ( .A1(n572), .A2(n571), .ZN(n575) );
  NAND2_X1 U633 ( .A1(G135), .A2(n864), .ZN(n573) );
  XNOR2_X1 U634 ( .A(KEYINPUT75), .B(n573), .ZN(n574) );
  NOR2_X1 U635 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U636 ( .A1(n577), .A2(n576), .ZN(n1005) );
  XNOR2_X1 U637 ( .A(G2096), .B(n1005), .ZN(n578) );
  OR2_X1 U638 ( .A1(G2100), .A2(n578), .ZN(G156) );
  NAND2_X1 U639 ( .A1(G50), .A2(n644), .ZN(n580) );
  NAND2_X1 U640 ( .A1(G62), .A2(n648), .ZN(n579) );
  NAND2_X1 U641 ( .A1(n580), .A2(n579), .ZN(n585) );
  NAND2_X1 U642 ( .A1(n637), .A2(G88), .ZN(n582) );
  NAND2_X1 U643 ( .A1(G75), .A2(n634), .ZN(n581) );
  NAND2_X1 U644 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U645 ( .A(KEYINPUT79), .B(n583), .Z(n584) );
  NOR2_X1 U646 ( .A1(n585), .A2(n584), .ZN(G166) );
  NAND2_X1 U647 ( .A1(G7), .A2(G661), .ZN(n586) );
  XNOR2_X1 U648 ( .A(n586), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U649 ( .A(G223), .ZN(n837) );
  NAND2_X1 U650 ( .A1(n837), .A2(G567), .ZN(n587) );
  XOR2_X1 U651 ( .A(KEYINPUT11), .B(n587), .Z(G234) );
  NAND2_X1 U652 ( .A1(n648), .A2(G56), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(KEYINPUT71), .ZN(n589) );
  XNOR2_X1 U654 ( .A(KEYINPUT14), .B(n589), .ZN(n596) );
  NAND2_X1 U655 ( .A1(n637), .A2(G81), .ZN(n590) );
  XOR2_X1 U656 ( .A(KEYINPUT12), .B(n590), .Z(n593) );
  NAND2_X1 U657 ( .A1(G68), .A2(n634), .ZN(n591) );
  XOR2_X1 U658 ( .A(KEYINPUT72), .B(n591), .Z(n592) );
  XNOR2_X1 U659 ( .A(KEYINPUT13), .B(n594), .ZN(n595) );
  NOR2_X1 U660 ( .A1(n596), .A2(n595), .ZN(n598) );
  NAND2_X1 U661 ( .A1(n644), .A2(G43), .ZN(n597) );
  NAND2_X1 U662 ( .A1(n598), .A2(n597), .ZN(n691) );
  INV_X1 U663 ( .A(G860), .ZN(n626) );
  OR2_X1 U664 ( .A1(n937), .A2(n626), .ZN(G153) );
  INV_X1 U665 ( .A(G171), .ZN(G301) );
  NAND2_X1 U666 ( .A1(G868), .A2(G301), .ZN(n607) );
  NAND2_X1 U667 ( .A1(G79), .A2(n634), .ZN(n600) );
  NAND2_X1 U668 ( .A1(G66), .A2(n648), .ZN(n599) );
  NAND2_X1 U669 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U670 ( .A1(G54), .A2(n644), .ZN(n602) );
  NAND2_X1 U671 ( .A1(G92), .A2(n637), .ZN(n601) );
  NAND2_X1 U672 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U673 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U674 ( .A(n605), .B(KEYINPUT15), .ZN(n919) );
  INV_X1 U675 ( .A(n919), .ZN(n706) );
  OR2_X1 U676 ( .A1(n706), .A2(G868), .ZN(n606) );
  NAND2_X1 U677 ( .A1(n607), .A2(n606), .ZN(G284) );
  NAND2_X1 U678 ( .A1(n637), .A2(G91), .ZN(n609) );
  NAND2_X1 U679 ( .A1(G78), .A2(n634), .ZN(n608) );
  NAND2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U681 ( .A(KEYINPUT68), .B(n610), .ZN(n614) );
  NAND2_X1 U682 ( .A1(G53), .A2(n644), .ZN(n612) );
  NAND2_X1 U683 ( .A1(G65), .A2(n648), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U685 ( .A1(n614), .A2(n613), .ZN(n926) );
  XNOR2_X1 U686 ( .A(n926), .B(KEYINPUT69), .ZN(G299) );
  XNOR2_X1 U687 ( .A(KEYINPUT73), .B(G868), .ZN(n615) );
  NOR2_X1 U688 ( .A1(G286), .A2(n615), .ZN(n617) );
  NOR2_X1 U689 ( .A1(G868), .A2(G299), .ZN(n616) );
  NOR2_X1 U690 ( .A1(n617), .A2(n616), .ZN(G297) );
  NAND2_X1 U691 ( .A1(n626), .A2(G559), .ZN(n618) );
  NAND2_X1 U692 ( .A1(n618), .A2(n706), .ZN(n619) );
  XNOR2_X1 U693 ( .A(n619), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U694 ( .A1(n706), .A2(G868), .ZN(n620) );
  NOR2_X1 U695 ( .A1(G559), .A2(n620), .ZN(n621) );
  XNOR2_X1 U696 ( .A(n621), .B(KEYINPUT74), .ZN(n623) );
  NOR2_X1 U697 ( .A1(n937), .A2(G868), .ZN(n622) );
  NOR2_X1 U698 ( .A1(n623), .A2(n622), .ZN(G282) );
  NAND2_X1 U699 ( .A1(G559), .A2(n706), .ZN(n624) );
  XOR2_X1 U700 ( .A(KEYINPUT76), .B(n624), .Z(n625) );
  XNOR2_X1 U701 ( .A(n937), .B(n625), .ZN(n660) );
  NAND2_X1 U702 ( .A1(n626), .A2(n660), .ZN(n633) );
  NAND2_X1 U703 ( .A1(G55), .A2(n644), .ZN(n628) );
  NAND2_X1 U704 ( .A1(G67), .A2(n648), .ZN(n627) );
  NAND2_X1 U705 ( .A1(n628), .A2(n627), .ZN(n632) );
  NAND2_X1 U706 ( .A1(n637), .A2(G93), .ZN(n630) );
  NAND2_X1 U707 ( .A1(G80), .A2(n634), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U709 ( .A1(n632), .A2(n631), .ZN(n662) );
  XOR2_X1 U710 ( .A(n633), .B(n662), .Z(G145) );
  XOR2_X1 U711 ( .A(KEYINPUT78), .B(KEYINPUT2), .Z(n636) );
  NAND2_X1 U712 ( .A1(G73), .A2(n634), .ZN(n635) );
  XNOR2_X1 U713 ( .A(n636), .B(n635), .ZN(n641) );
  NAND2_X1 U714 ( .A1(G48), .A2(n644), .ZN(n639) );
  NAND2_X1 U715 ( .A1(G86), .A2(n637), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U717 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U718 ( .A1(G61), .A2(n648), .ZN(n642) );
  NAND2_X1 U719 ( .A1(n643), .A2(n642), .ZN(G305) );
  NAND2_X1 U720 ( .A1(G49), .A2(n644), .ZN(n646) );
  NAND2_X1 U721 ( .A1(G74), .A2(G651), .ZN(n645) );
  NAND2_X1 U722 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U723 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U724 ( .A1(G87), .A2(n649), .ZN(n650) );
  XOR2_X1 U725 ( .A(KEYINPUT77), .B(n650), .Z(n651) );
  NAND2_X1 U726 ( .A1(n652), .A2(n651), .ZN(G288) );
  XNOR2_X1 U727 ( .A(n662), .B(G290), .ZN(n657) );
  XNOR2_X1 U728 ( .A(KEYINPUT19), .B(KEYINPUT81), .ZN(n654) );
  XNOR2_X1 U729 ( .A(G305), .B(KEYINPUT80), .ZN(n653) );
  XNOR2_X1 U730 ( .A(n654), .B(n653), .ZN(n655) );
  XOR2_X1 U731 ( .A(n655), .B(G288), .Z(n656) );
  XNOR2_X1 U732 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U733 ( .A(G166), .B(n658), .ZN(n659) );
  XNOR2_X1 U734 ( .A(n659), .B(G299), .ZN(n884) );
  XNOR2_X1 U735 ( .A(n660), .B(n884), .ZN(n661) );
  NAND2_X1 U736 ( .A1(n661), .A2(G868), .ZN(n664) );
  OR2_X1 U737 ( .A1(n662), .A2(G868), .ZN(n663) );
  NAND2_X1 U738 ( .A1(n664), .A2(n663), .ZN(G295) );
  NAND2_X1 U739 ( .A1(G2078), .A2(G2084), .ZN(n665) );
  XOR2_X1 U740 ( .A(KEYINPUT20), .B(n665), .Z(n666) );
  NAND2_X1 U741 ( .A1(G2090), .A2(n666), .ZN(n668) );
  XNOR2_X1 U742 ( .A(KEYINPUT21), .B(KEYINPUT82), .ZN(n667) );
  XNOR2_X1 U743 ( .A(n668), .B(n667), .ZN(n669) );
  NAND2_X1 U744 ( .A1(G2072), .A2(n669), .ZN(G158) );
  XOR2_X1 U745 ( .A(KEYINPUT70), .B(G57), .Z(G237) );
  XNOR2_X1 U746 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U747 ( .A1(G108), .A2(G120), .ZN(n670) );
  NOR2_X1 U748 ( .A1(G237), .A2(n670), .ZN(n671) );
  NAND2_X1 U749 ( .A1(G69), .A2(n671), .ZN(n841) );
  NAND2_X1 U750 ( .A1(n841), .A2(G567), .ZN(n678) );
  XOR2_X1 U751 ( .A(KEYINPUT83), .B(KEYINPUT22), .Z(n673) );
  NAND2_X1 U752 ( .A1(G132), .A2(G82), .ZN(n672) );
  XNOR2_X1 U753 ( .A(n673), .B(n672), .ZN(n674) );
  NOR2_X1 U754 ( .A1(G218), .A2(n674), .ZN(n675) );
  NAND2_X1 U755 ( .A1(G96), .A2(n675), .ZN(n676) );
  XNOR2_X1 U756 ( .A(KEYINPUT84), .B(n676), .ZN(n842) );
  NAND2_X1 U757 ( .A1(n842), .A2(G2106), .ZN(n677) );
  NAND2_X1 U758 ( .A1(n678), .A2(n677), .ZN(n917) );
  NAND2_X1 U759 ( .A1(G661), .A2(G483), .ZN(n679) );
  XOR2_X1 U760 ( .A(KEYINPUT85), .B(n679), .Z(n680) );
  NOR2_X1 U761 ( .A1(n917), .A2(n680), .ZN(n840) );
  NAND2_X1 U762 ( .A1(n840), .A2(G36), .ZN(G176) );
  INV_X1 U763 ( .A(G166), .ZN(G303) );
  INV_X1 U764 ( .A(G1384), .ZN(n681) );
  AND2_X1 U765 ( .A1(G138), .A2(n681), .ZN(n682) );
  NAND2_X1 U766 ( .A1(n864), .A2(n682), .ZN(n685) );
  NAND2_X1 U767 ( .A1(n685), .A2(n684), .ZN(n783) );
  AND2_X1 U768 ( .A1(G160), .A2(G40), .ZN(n782) );
  NAND2_X2 U769 ( .A1(n783), .A2(n782), .ZN(n734) );
  INV_X1 U770 ( .A(G1996), .ZN(n973) );
  NOR2_X1 U771 ( .A1(n734), .A2(n973), .ZN(n687) );
  XNOR2_X1 U772 ( .A(n687), .B(n686), .ZN(n689) );
  NAND2_X1 U773 ( .A1(n734), .A2(G1341), .ZN(n688) );
  NAND2_X1 U774 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U775 ( .A1(n691), .A2(n690), .ZN(n693) );
  XNOR2_X1 U776 ( .A(n693), .B(n692), .ZN(n708) );
  NOR2_X1 U777 ( .A1(n708), .A2(n919), .ZN(n694) );
  XNOR2_X1 U778 ( .A(n694), .B(KEYINPUT96), .ZN(n695) );
  INV_X1 U779 ( .A(n695), .ZN(n703) );
  XNOR2_X1 U780 ( .A(KEYINPUT95), .B(n734), .ZN(n718) );
  NAND2_X1 U781 ( .A1(G2067), .A2(n718), .ZN(n697) );
  NAND2_X1 U782 ( .A1(G1348), .A2(n734), .ZN(n696) );
  NAND2_X1 U783 ( .A1(n697), .A2(n696), .ZN(n701) );
  NAND2_X1 U784 ( .A1(n718), .A2(G2072), .ZN(n698) );
  XNOR2_X1 U785 ( .A(n698), .B(KEYINPUT27), .ZN(n700) );
  INV_X1 U786 ( .A(G1956), .ZN(n908) );
  NOR2_X1 U787 ( .A1(n908), .A2(n718), .ZN(n699) );
  NOR2_X1 U788 ( .A1(n700), .A2(n699), .ZN(n709) );
  NAND2_X1 U789 ( .A1(n709), .A2(n926), .ZN(n704) );
  AND2_X1 U790 ( .A1(n701), .A2(n704), .ZN(n702) );
  NAND2_X1 U791 ( .A1(n703), .A2(n702), .ZN(n714) );
  INV_X1 U792 ( .A(n704), .ZN(n705) );
  NOR2_X1 U793 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U794 ( .A1(n708), .A2(n707), .ZN(n712) );
  NOR2_X1 U795 ( .A1(n926), .A2(n709), .ZN(n710) );
  XOR2_X1 U796 ( .A(n710), .B(KEYINPUT28), .Z(n711) );
  AND2_X1 U797 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U798 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U799 ( .A(n715), .B(KEYINPUT29), .ZN(n722) );
  INV_X1 U800 ( .A(n734), .ZN(n716) );
  NOR2_X1 U801 ( .A1(n716), .A2(G1961), .ZN(n717) );
  XOR2_X1 U802 ( .A(KEYINPUT94), .B(n717), .Z(n720) );
  XNOR2_X1 U803 ( .A(G2078), .B(KEYINPUT25), .ZN(n972) );
  NAND2_X1 U804 ( .A1(n718), .A2(n972), .ZN(n719) );
  NAND2_X1 U805 ( .A1(n720), .A2(n719), .ZN(n728) );
  AND2_X1 U806 ( .A1(G171), .A2(n728), .ZN(n721) );
  NOR2_X1 U807 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U808 ( .A(n723), .B(KEYINPUT97), .ZN(n733) );
  NAND2_X1 U809 ( .A1(G8), .A2(n734), .ZN(n768) );
  NOR2_X1 U810 ( .A1(G1966), .A2(n768), .ZN(n748) );
  NOR2_X1 U811 ( .A1(n734), .A2(G2084), .ZN(n724) );
  XNOR2_X1 U812 ( .A(n724), .B(KEYINPUT93), .ZN(n744) );
  NAND2_X1 U813 ( .A1(G8), .A2(n744), .ZN(n725) );
  NOR2_X1 U814 ( .A1(n748), .A2(n725), .ZN(n726) );
  XOR2_X1 U815 ( .A(KEYINPUT30), .B(n726), .Z(n727) );
  NOR2_X1 U816 ( .A1(G168), .A2(n727), .ZN(n730) );
  NOR2_X1 U817 ( .A1(G171), .A2(n728), .ZN(n729) );
  NOR2_X1 U818 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U819 ( .A(KEYINPUT31), .B(n731), .Z(n732) );
  NAND2_X1 U820 ( .A1(n733), .A2(n732), .ZN(n746) );
  NAND2_X1 U821 ( .A1(n746), .A2(G286), .ZN(n739) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n768), .ZN(n736) );
  NOR2_X1 U823 ( .A1(G2090), .A2(n734), .ZN(n735) );
  NOR2_X1 U824 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U825 ( .A1(n737), .A2(G303), .ZN(n738) );
  NAND2_X1 U826 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U827 ( .A(n740), .B(KEYINPUT98), .ZN(n741) );
  NAND2_X1 U828 ( .A1(n741), .A2(G8), .ZN(n743) );
  XOR2_X1 U829 ( .A(KEYINPUT32), .B(KEYINPUT99), .Z(n742) );
  XNOR2_X1 U830 ( .A(n743), .B(n742), .ZN(n752) );
  INV_X1 U831 ( .A(n744), .ZN(n745) );
  NAND2_X1 U832 ( .A1(G8), .A2(n745), .ZN(n750) );
  INV_X1 U833 ( .A(n746), .ZN(n747) );
  NOR2_X1 U834 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U835 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U836 ( .A1(n752), .A2(n751), .ZN(n764) );
  NOR2_X1 U837 ( .A1(G2090), .A2(G303), .ZN(n753) );
  NAND2_X1 U838 ( .A1(G8), .A2(n753), .ZN(n754) );
  NAND2_X1 U839 ( .A1(n764), .A2(n754), .ZN(n755) );
  XNOR2_X1 U840 ( .A(n755), .B(KEYINPUT102), .ZN(n756) );
  NAND2_X1 U841 ( .A1(n756), .A2(n768), .ZN(n758) );
  INV_X1 U842 ( .A(KEYINPUT103), .ZN(n757) );
  XNOR2_X1 U843 ( .A(n758), .B(n757), .ZN(n781) );
  NOR2_X1 U844 ( .A1(G288), .A2(G1976), .ZN(n759) );
  XNOR2_X1 U845 ( .A(n759), .B(KEYINPUT100), .ZN(n763) );
  NAND2_X1 U846 ( .A1(KEYINPUT33), .A2(n763), .ZN(n760) );
  NOR2_X1 U847 ( .A1(n768), .A2(n760), .ZN(n761) );
  XNOR2_X1 U848 ( .A(G1981), .B(G305), .ZN(n924) );
  NOR2_X1 U849 ( .A1(n761), .A2(n924), .ZN(n767) );
  NOR2_X1 U850 ( .A1(G1971), .A2(G303), .ZN(n762) );
  NOR2_X1 U851 ( .A1(n763), .A2(n762), .ZN(n932) );
  NAND2_X1 U852 ( .A1(n932), .A2(n764), .ZN(n765) );
  NAND2_X1 U853 ( .A1(n767), .A2(n765), .ZN(n770) );
  NAND2_X1 U854 ( .A1(G288), .A2(G1976), .ZN(n766) );
  XNOR2_X1 U855 ( .A(n766), .B(KEYINPUT101), .ZN(n930) );
  NAND2_X1 U856 ( .A1(KEYINPUT33), .A2(n767), .ZN(n773) );
  AND2_X1 U857 ( .A1(n773), .A2(n768), .ZN(n771) );
  OR2_X1 U858 ( .A1(n930), .A2(n771), .ZN(n769) );
  NOR2_X1 U859 ( .A1(n770), .A2(n769), .ZN(n779) );
  INV_X1 U860 ( .A(n771), .ZN(n777) );
  NOR2_X1 U861 ( .A1(G1981), .A2(G305), .ZN(n772) );
  XNOR2_X1 U862 ( .A(KEYINPUT24), .B(n772), .ZN(n775) );
  INV_X1 U863 ( .A(n773), .ZN(n774) );
  OR2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n776) );
  AND2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U866 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U867 ( .A1(n781), .A2(n780), .ZN(n821) );
  XNOR2_X1 U868 ( .A(G1986), .B(G290), .ZN(n929) );
  INV_X1 U869 ( .A(n782), .ZN(n784) );
  NOR2_X1 U870 ( .A1(n784), .A2(n783), .ZN(n832) );
  NAND2_X1 U871 ( .A1(n929), .A2(n832), .ZN(n819) );
  NAND2_X1 U872 ( .A1(G104), .A2(n866), .ZN(n786) );
  NAND2_X1 U873 ( .A1(G140), .A2(n864), .ZN(n785) );
  NAND2_X1 U874 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U875 ( .A(KEYINPUT34), .B(n787), .ZN(n792) );
  NAND2_X1 U876 ( .A1(G128), .A2(n516), .ZN(n789) );
  NAND2_X1 U877 ( .A1(G116), .A2(n861), .ZN(n788) );
  NAND2_X1 U878 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U879 ( .A(n790), .B(KEYINPUT35), .Z(n791) );
  NOR2_X1 U880 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U881 ( .A(KEYINPUT36), .B(n793), .Z(n794) );
  XOR2_X1 U882 ( .A(KEYINPUT86), .B(n794), .Z(n851) );
  XNOR2_X1 U883 ( .A(KEYINPUT37), .B(G2067), .ZN(n830) );
  NOR2_X1 U884 ( .A1(n851), .A2(n830), .ZN(n1002) );
  NAND2_X1 U885 ( .A1(n1002), .A2(n832), .ZN(n795) );
  XOR2_X1 U886 ( .A(KEYINPUT87), .B(n795), .Z(n828) );
  NAND2_X1 U887 ( .A1(G95), .A2(n866), .ZN(n796) );
  XNOR2_X1 U888 ( .A(n796), .B(KEYINPUT91), .ZN(n803) );
  NAND2_X1 U889 ( .A1(n861), .A2(G107), .ZN(n797) );
  XNOR2_X1 U890 ( .A(KEYINPUT89), .B(n797), .ZN(n800) );
  NAND2_X1 U891 ( .A1(n516), .A2(G119), .ZN(n798) );
  XOR2_X1 U892 ( .A(KEYINPUT88), .B(n798), .Z(n799) );
  NOR2_X1 U893 ( .A1(n800), .A2(n799), .ZN(n801) );
  XOR2_X1 U894 ( .A(KEYINPUT90), .B(n801), .Z(n802) );
  NOR2_X1 U895 ( .A1(n803), .A2(n802), .ZN(n805) );
  NAND2_X1 U896 ( .A1(n864), .A2(G131), .ZN(n804) );
  NAND2_X1 U897 ( .A1(n805), .A2(n804), .ZN(n850) );
  AND2_X1 U898 ( .A1(n850), .A2(G1991), .ZN(n815) );
  NAND2_X1 U899 ( .A1(G105), .A2(n866), .ZN(n806) );
  XNOR2_X1 U900 ( .A(n806), .B(KEYINPUT38), .ZN(n813) );
  NAND2_X1 U901 ( .A1(G141), .A2(n864), .ZN(n808) );
  NAND2_X1 U902 ( .A1(G129), .A2(n516), .ZN(n807) );
  NAND2_X1 U903 ( .A1(n808), .A2(n807), .ZN(n811) );
  NAND2_X1 U904 ( .A1(n861), .A2(G117), .ZN(n809) );
  XOR2_X1 U905 ( .A(KEYINPUT92), .B(n809), .Z(n810) );
  NOR2_X1 U906 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n875) );
  AND2_X1 U908 ( .A1(n875), .A2(G1996), .ZN(n814) );
  NOR2_X1 U909 ( .A1(n815), .A2(n814), .ZN(n1004) );
  INV_X1 U910 ( .A(n832), .ZN(n816) );
  NOR2_X1 U911 ( .A1(n1004), .A2(n816), .ZN(n825) );
  INV_X1 U912 ( .A(n825), .ZN(n817) );
  AND2_X1 U913 ( .A1(n828), .A2(n817), .ZN(n818) );
  AND2_X1 U914 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U915 ( .A1(n821), .A2(n820), .ZN(n835) );
  NOR2_X1 U916 ( .A1(n875), .A2(G1996), .ZN(n822) );
  XNOR2_X1 U917 ( .A(n822), .B(KEYINPUT104), .ZN(n999) );
  NOR2_X1 U918 ( .A1(G1986), .A2(G290), .ZN(n823) );
  NOR2_X1 U919 ( .A1(G1991), .A2(n850), .ZN(n1008) );
  NOR2_X1 U920 ( .A1(n823), .A2(n1008), .ZN(n824) );
  NOR2_X1 U921 ( .A1(n825), .A2(n824), .ZN(n826) );
  NOR2_X1 U922 ( .A1(n999), .A2(n826), .ZN(n827) );
  XNOR2_X1 U923 ( .A(n827), .B(KEYINPUT39), .ZN(n829) );
  NAND2_X1 U924 ( .A1(n829), .A2(n828), .ZN(n831) );
  NAND2_X1 U925 ( .A1(n851), .A2(n830), .ZN(n1003) );
  NAND2_X1 U926 ( .A1(n831), .A2(n1003), .ZN(n833) );
  NAND2_X1 U927 ( .A1(n833), .A2(n832), .ZN(n834) );
  NAND2_X1 U928 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U929 ( .A(KEYINPUT40), .B(n836), .ZN(G329) );
  NAND2_X1 U930 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U931 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U932 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U934 ( .A1(n840), .A2(n839), .ZN(G188) );
  XOR2_X1 U935 ( .A(G120), .B(KEYINPUT106), .Z(G236) );
  INV_X1 U937 ( .A(G132), .ZN(G219) );
  INV_X1 U938 ( .A(G108), .ZN(G238) );
  INV_X1 U939 ( .A(G96), .ZN(G221) );
  INV_X1 U940 ( .A(G82), .ZN(G220) );
  INV_X1 U941 ( .A(G69), .ZN(G235) );
  NOR2_X1 U942 ( .A1(n842), .A2(n841), .ZN(G325) );
  INV_X1 U943 ( .A(G325), .ZN(G261) );
  NAND2_X1 U944 ( .A1(G124), .A2(n516), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n843), .B(KEYINPUT44), .ZN(n845) );
  NAND2_X1 U946 ( .A1(n866), .A2(G100), .ZN(n844) );
  NAND2_X1 U947 ( .A1(n845), .A2(n844), .ZN(n849) );
  NAND2_X1 U948 ( .A1(G136), .A2(n864), .ZN(n847) );
  NAND2_X1 U949 ( .A1(G112), .A2(n861), .ZN(n846) );
  NAND2_X1 U950 ( .A1(n847), .A2(n846), .ZN(n848) );
  NOR2_X1 U951 ( .A1(n849), .A2(n848), .ZN(G162) );
  XOR2_X1 U952 ( .A(n851), .B(n850), .Z(n860) );
  NAND2_X1 U953 ( .A1(G103), .A2(n866), .ZN(n853) );
  NAND2_X1 U954 ( .A1(G139), .A2(n864), .ZN(n852) );
  NAND2_X1 U955 ( .A1(n853), .A2(n852), .ZN(n859) );
  NAND2_X1 U956 ( .A1(n861), .A2(G115), .ZN(n854) );
  XNOR2_X1 U957 ( .A(n854), .B(KEYINPUT112), .ZN(n856) );
  NAND2_X1 U958 ( .A1(G127), .A2(n516), .ZN(n855) );
  NAND2_X1 U959 ( .A1(n856), .A2(n855), .ZN(n857) );
  XOR2_X1 U960 ( .A(KEYINPUT47), .B(n857), .Z(n858) );
  NOR2_X1 U961 ( .A1(n859), .A2(n858), .ZN(n1014) );
  XNOR2_X1 U962 ( .A(n860), .B(n1014), .ZN(n882) );
  NAND2_X1 U963 ( .A1(G130), .A2(n516), .ZN(n863) );
  NAND2_X1 U964 ( .A1(G118), .A2(n861), .ZN(n862) );
  NAND2_X1 U965 ( .A1(n863), .A2(n862), .ZN(n871) );
  NAND2_X1 U966 ( .A1(n864), .A2(G142), .ZN(n865) );
  XNOR2_X1 U967 ( .A(n865), .B(KEYINPUT110), .ZN(n868) );
  NAND2_X1 U968 ( .A1(G106), .A2(n866), .ZN(n867) );
  NAND2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U970 ( .A(KEYINPUT45), .B(n869), .Z(n870) );
  NOR2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n879) );
  XOR2_X1 U972 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n873) );
  XNOR2_X1 U973 ( .A(G164), .B(KEYINPUT111), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n873), .B(n872), .ZN(n874) );
  XOR2_X1 U975 ( .A(n874), .B(G162), .Z(n877) );
  XOR2_X1 U976 ( .A(G160), .B(n875), .Z(n876) );
  XNOR2_X1 U977 ( .A(n877), .B(n876), .ZN(n878) );
  XNOR2_X1 U978 ( .A(n879), .B(n878), .ZN(n880) );
  XNOR2_X1 U979 ( .A(n880), .B(n1005), .ZN(n881) );
  XNOR2_X1 U980 ( .A(n882), .B(n881), .ZN(n883) );
  NOR2_X1 U981 ( .A1(G37), .A2(n883), .ZN(G395) );
  XNOR2_X1 U982 ( .A(G286), .B(n937), .ZN(n885) );
  XNOR2_X1 U983 ( .A(n885), .B(n884), .ZN(n887) );
  XOR2_X1 U984 ( .A(n919), .B(G171), .Z(n886) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n888) );
  NOR2_X1 U986 ( .A1(G37), .A2(n888), .ZN(G397) );
  XOR2_X1 U987 ( .A(G2678), .B(KEYINPUT107), .Z(n890) );
  XNOR2_X1 U988 ( .A(KEYINPUT43), .B(KEYINPUT108), .ZN(n889) );
  XNOR2_X1 U989 ( .A(n890), .B(n889), .ZN(n894) );
  XOR2_X1 U990 ( .A(KEYINPUT42), .B(G2090), .Z(n892) );
  XNOR2_X1 U991 ( .A(G2067), .B(G2072), .ZN(n891) );
  XNOR2_X1 U992 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U993 ( .A(n894), .B(n893), .Z(n896) );
  XNOR2_X1 U994 ( .A(G2096), .B(G2100), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n898) );
  XOR2_X1 U996 ( .A(G2078), .B(G2084), .Z(n897) );
  XNOR2_X1 U997 ( .A(n898), .B(n897), .ZN(G227) );
  XOR2_X1 U998 ( .A(G1981), .B(G1961), .Z(n900) );
  XNOR2_X1 U999 ( .A(G1986), .B(G1966), .ZN(n899) );
  XNOR2_X1 U1000 ( .A(n900), .B(n899), .ZN(n904) );
  XOR2_X1 U1001 ( .A(G1971), .B(G1976), .Z(n902) );
  XNOR2_X1 U1002 ( .A(G1996), .B(G1991), .ZN(n901) );
  XNOR2_X1 U1003 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1004 ( .A(n904), .B(n903), .Z(n906) );
  XNOR2_X1 U1005 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n905) );
  XNOR2_X1 U1006 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1007 ( .A(G2474), .B(n907), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(n909), .B(n908), .ZN(G229) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n910) );
  XNOR2_X1 U1010 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1011 ( .A1(G397), .A2(n911), .ZN(n914) );
  NOR2_X1 U1012 ( .A1(n917), .A2(G401), .ZN(n912) );
  XOR2_X1 U1013 ( .A(KEYINPUT113), .B(n912), .Z(n913) );
  NAND2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(n915) );
  NOR2_X1 U1015 ( .A1(G395), .A2(n915), .ZN(n916) );
  XNOR2_X1 U1016 ( .A(KEYINPUT114), .B(n916), .ZN(G308) );
  INV_X1 U1017 ( .A(G308), .ZN(G225) );
  INV_X1 U1018 ( .A(n917), .ZN(G319) );
  INV_X1 U1019 ( .A(G16), .ZN(n968) );
  XOR2_X1 U1020 ( .A(KEYINPUT56), .B(KEYINPUT122), .Z(n918) );
  XNOR2_X1 U1021 ( .A(n968), .B(n918), .ZN(n943) );
  XNOR2_X1 U1022 ( .A(G171), .B(G1961), .ZN(n921) );
  XOR2_X1 U1023 ( .A(G1348), .B(n919), .Z(n920) );
  NAND2_X1 U1024 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1025 ( .A(n922), .B(KEYINPUT123), .ZN(n941) );
  XOR2_X1 U1026 ( .A(G168), .B(G1966), .Z(n923) );
  NOR2_X1 U1027 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1028 ( .A(KEYINPUT57), .B(n925), .Z(n936) );
  XNOR2_X1 U1029 ( .A(G1956), .B(n926), .ZN(n928) );
  NAND2_X1 U1030 ( .A1(G1971), .A2(G303), .ZN(n927) );
  NAND2_X1 U1031 ( .A1(n928), .A2(n927), .ZN(n934) );
  NOR2_X1 U1032 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1033 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n939) );
  XNOR2_X1 U1036 ( .A(G1341), .B(n937), .ZN(n938) );
  NOR2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1038 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n970) );
  XNOR2_X1 U1040 ( .A(KEYINPUT125), .B(G1981), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(n944), .B(G6), .ZN(n951) );
  XOR2_X1 U1042 ( .A(G4), .B(KEYINPUT126), .Z(n946) );
  XNOR2_X1 U1043 ( .A(G1348), .B(KEYINPUT59), .ZN(n945) );
  XNOR2_X1 U1044 ( .A(n946), .B(n945), .ZN(n949) );
  XNOR2_X1 U1045 ( .A(KEYINPUT124), .B(G1341), .ZN(n947) );
  XNOR2_X1 U1046 ( .A(G19), .B(n947), .ZN(n948) );
  NOR2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n953) );
  XNOR2_X1 U1049 ( .A(G20), .B(G1956), .ZN(n952) );
  NOR2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(KEYINPUT60), .B(n954), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(G1966), .B(G21), .ZN(n956) );
  XNOR2_X1 U1053 ( .A(G1961), .B(G5), .ZN(n955) );
  NOR2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n965) );
  XNOR2_X1 U1056 ( .A(G1976), .B(G23), .ZN(n960) );
  XNOR2_X1 U1057 ( .A(G1971), .B(G22), .ZN(n959) );
  NOR2_X1 U1058 ( .A1(n960), .A2(n959), .ZN(n962) );
  XOR2_X1 U1059 ( .A(G1986), .B(G24), .Z(n961) );
  NAND2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1061 ( .A(KEYINPUT58), .B(n963), .ZN(n964) );
  NOR2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1063 ( .A(KEYINPUT61), .B(n966), .ZN(n967) );
  NAND2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1066 ( .A(KEYINPUT127), .B(n971), .ZN(n997) );
  XOR2_X1 U1067 ( .A(G2090), .B(G35), .Z(n989) );
  XNOR2_X1 U1068 ( .A(G1991), .B(G25), .ZN(n984) );
  XNOR2_X1 U1069 ( .A(n972), .B(G27), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(KEYINPUT118), .B(G32), .ZN(n974) );
  XNOR2_X1 U1071 ( .A(n974), .B(n973), .ZN(n975) );
  NAND2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(G2067), .B(G26), .ZN(n978) );
  XNOR2_X1 U1074 ( .A(G2072), .B(G33), .ZN(n977) );
  NOR2_X1 U1075 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1076 ( .A(n979), .B(KEYINPUT117), .ZN(n980) );
  NOR2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1078 ( .A(KEYINPUT119), .B(n982), .ZN(n983) );
  NOR2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1080 ( .A1(n985), .A2(G28), .ZN(n986) );
  XNOR2_X1 U1081 ( .A(n986), .B(KEYINPUT53), .ZN(n987) );
  XNOR2_X1 U1082 ( .A(n987), .B(KEYINPUT120), .ZN(n988) );
  NAND2_X1 U1083 ( .A1(n989), .A2(n988), .ZN(n992) );
  XNOR2_X1 U1084 ( .A(G34), .B(G2084), .ZN(n990) );
  XNOR2_X1 U1085 ( .A(KEYINPUT54), .B(n990), .ZN(n991) );
  NOR2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1087 ( .A(KEYINPUT55), .B(n993), .Z(n994) );
  NOR2_X1 U1088 ( .A1(G29), .A2(n994), .ZN(n995) );
  XNOR2_X1 U1089 ( .A(KEYINPUT121), .B(n995), .ZN(n996) );
  NAND2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n1026) );
  XOR2_X1 U1091 ( .A(G2090), .B(G162), .Z(n998) );
  NOR2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1093 ( .A(n1000), .B(KEYINPUT51), .ZN(n1001) );
  NOR2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1013) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1011) );
  XNOR2_X1 U1096 ( .A(G160), .B(G2084), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(KEYINPUT115), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1019) );
  XOR2_X1 U1102 ( .A(G2072), .B(n1014), .Z(n1016) );
  XOR2_X1 U1103 ( .A(G164), .B(G2078), .Z(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1105 ( .A(KEYINPUT50), .B(n1017), .Z(n1018) );
  NOR2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(KEYINPUT52), .B(n1020), .ZN(n1022) );
  INV_X1 U1108 ( .A(KEYINPUT55), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1023), .A2(G29), .ZN(n1024) );
  XOR2_X1 U1111 ( .A(KEYINPUT116), .B(n1024), .Z(n1025) );
  NOR2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1113 ( .A1(n1027), .A2(G11), .ZN(n1028) );
  XOR2_X1 U1114 ( .A(KEYINPUT62), .B(n1028), .Z(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

