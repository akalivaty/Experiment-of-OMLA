//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 1 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 0 0 0 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1220, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n207), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT1), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(KEYINPUT64), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT64), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G20), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n202), .A2(new_n203), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(G50), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n207), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT0), .ZN(new_n228));
  AOI22_X1  g0028(.A1(new_n222), .A2(new_n225), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n229), .B1(new_n228), .B2(new_n227), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n215), .A2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  NAND2_X1  g0039(.A1(new_n201), .A2(G68), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n203), .A2(G50), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n244), .B(KEYINPUT65), .Z(new_n245));
  INV_X1    g0045(.A(G107), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G97), .ZN(new_n247));
  INV_X1    g0047(.A(G97), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G107), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n245), .B(new_n252), .ZN(G351));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  AND2_X1   g0054(.A1(new_n254), .A2(new_n221), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n216), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  AOI22_X1  g0058(.A1(new_n258), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n220), .A2(G33), .A3(G77), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n255), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  XOR2_X1   g0061(.A(new_n261), .B(KEYINPUT11), .Z(new_n262));
  NOR2_X1   g0062(.A1(new_n216), .A2(G1), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT71), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(new_n264), .A3(G13), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(G13), .A3(G20), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT71), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n255), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n266), .A2(G20), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT12), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G68), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT12), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(G68), .ZN(new_n277));
  AOI22_X1  g0077(.A1(new_n269), .A2(new_n277), .B1(new_n276), .B2(new_n267), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n262), .A2(new_n275), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT13), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT67), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT66), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n283), .B(new_n266), .C1(G41), .C2(G45), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G1), .A3(G13), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(new_n286), .A3(G274), .ZN(new_n287));
  OR2_X1    g0087(.A1(G41), .A2(G45), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n283), .B1(new_n288), .B2(new_n266), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n282), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G274), .ZN(new_n291));
  INV_X1    g0091(.A(new_n221), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n291), .B1(new_n292), .B2(new_n285), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT66), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n293), .A2(new_n295), .A3(KEYINPUT67), .A4(new_n284), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT3), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G33), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n298), .A2(new_n300), .A3(G232), .A4(G1698), .ZN(new_n301));
  INV_X1    g0101(.A(G1698), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n298), .A2(new_n300), .A3(G226), .A4(new_n302), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n301), .B(new_n303), .C1(new_n256), .C2(new_n248), .ZN(new_n304));
  INV_X1    g0104(.A(new_n286), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n286), .A2(new_n294), .ZN(new_n307));
  INV_X1    g0107(.A(G238), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  AND4_X1   g0110(.A1(new_n281), .A2(new_n297), .A3(new_n306), .A4(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n309), .B1(new_n290), .B2(new_n296), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n281), .B1(new_n312), .B2(new_n306), .ZN(new_n313));
  OAI21_X1  g0113(.A(G169), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT74), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(KEYINPUT14), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n297), .A2(new_n306), .A3(new_n310), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT13), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n312), .A2(new_n281), .A3(new_n306), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n316), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n321), .A2(G169), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n317), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n319), .A2(G179), .A3(new_n320), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n315), .A2(KEYINPUT14), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n280), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n321), .A2(G200), .ZN(new_n331));
  INV_X1    g0131(.A(G190), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n280), .B(new_n331), .C1(new_n332), .C2(new_n321), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n272), .A2(G50), .ZN(new_n335));
  XNOR2_X1  g0135(.A(new_n335), .B(KEYINPUT68), .ZN(new_n336));
  INV_X1    g0136(.A(new_n267), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n270), .A2(new_n337), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n336), .A2(new_n338), .B1(new_n201), .B2(new_n337), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  XOR2_X1   g0140(.A(KEYINPUT8), .B(G58), .Z(new_n341));
  NAND3_X1  g0141(.A1(new_n341), .A2(G33), .A3(new_n220), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n258), .A2(G150), .B1(new_n204), .B2(G20), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n344), .A2(new_n255), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g0146(.A(KEYINPUT3), .B(G33), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n347), .A2(G222), .A3(new_n302), .ZN(new_n348));
  INV_X1    g0148(.A(G77), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(G1698), .ZN(new_n350));
  INV_X1    g0150(.A(G223), .ZN(new_n351));
  OAI221_X1 g0151(.A(new_n348), .B1(new_n349), .B2(new_n347), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n305), .ZN(new_n353));
  INV_X1    g0153(.A(new_n307), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n290), .A2(new_n296), .B1(G226), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(G169), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  OR3_X1    g0156(.A1(new_n346), .A2(new_n356), .A3(KEYINPUT69), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT69), .B1(new_n346), .B2(new_n356), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n353), .A2(new_n355), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n357), .B(new_n358), .C1(G179), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(G200), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(new_n332), .B2(new_n359), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT9), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n340), .B2(new_n345), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n339), .B(KEYINPUT9), .C1(new_n255), .C2(new_n344), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(KEYINPUT72), .B1(KEYINPUT73), .B2(KEYINPUT10), .ZN(new_n367));
  OR3_X1    g0167(.A1(new_n362), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(KEYINPUT72), .B1(new_n364), .B2(new_n365), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT73), .ZN(new_n370));
  NOR3_X1   g0170(.A1(new_n369), .A2(new_n362), .A3(new_n370), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n360), .B(new_n368), .C1(new_n371), .C2(KEYINPUT10), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n290), .A2(new_n296), .B1(G232), .B2(new_n354), .ZN(new_n373));
  INV_X1    g0173(.A(G179), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n347), .A2(G226), .A3(G1698), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n347), .A2(G223), .A3(new_n302), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G33), .A2(G87), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n305), .ZN(new_n379));
  AND3_X1   g0179(.A1(new_n373), .A2(new_n374), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(G169), .B1(new_n373), .B2(new_n379), .ZN(new_n381));
  OAI21_X1  g0181(.A(KEYINPUT77), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n354), .A2(G232), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n379), .A2(new_n297), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G169), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT77), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n373), .A2(new_n374), .A3(new_n379), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n341), .ZN(new_n390));
  NOR3_X1   g0190(.A1(new_n390), .A2(new_n270), .A3(new_n263), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n391), .B1(new_n337), .B2(new_n390), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G58), .A2(G68), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n223), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(G20), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n258), .A2(G159), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(KEYINPUT75), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT75), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n216), .B1(new_n223), .B2(new_n393), .ZN(new_n399));
  INV_X1    g0199(.A(G159), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n257), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n398), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n397), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT7), .B1(new_n347), .B2(G20), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n298), .A2(new_n300), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n220), .A2(new_n405), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n404), .B(G68), .C1(new_n406), .C2(KEYINPUT7), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n403), .A2(new_n407), .A3(KEYINPUT16), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n270), .ZN(new_n409));
  XOR2_X1   g0209(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n410));
  INV_X1    g0210(.A(KEYINPUT7), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n405), .A2(new_n411), .A3(new_n216), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n217), .A2(new_n219), .B1(new_n298), .B2(new_n300), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n412), .B(G68), .C1(new_n413), .C2(new_n411), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n399), .A2(new_n401), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n410), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n392), .B1(new_n409), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n382), .A2(new_n389), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT18), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n382), .A2(new_n389), .A3(new_n417), .A4(KEYINPUT18), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n384), .A2(G200), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n373), .A2(G190), .A3(new_n379), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT17), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n414), .A2(new_n415), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n270), .B(new_n408), .C1(new_n427), .C2(new_n410), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n425), .A2(new_n426), .A3(new_n428), .A4(new_n392), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n428), .A2(new_n392), .A3(new_n424), .A4(new_n423), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT17), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n422), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n347), .A2(G232), .A3(new_n302), .ZN(new_n434));
  OAI221_X1 g0234(.A(new_n434), .B1(new_n246), .B2(new_n347), .C1(new_n350), .C2(new_n308), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n305), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n290), .A2(new_n296), .B1(G244), .B2(new_n354), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT70), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n436), .A2(KEYINPUT70), .A3(new_n437), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G190), .ZN(new_n443));
  INV_X1    g0243(.A(new_n220), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n444), .A2(G77), .B1(new_n341), .B2(new_n258), .ZN(new_n445));
  XOR2_X1   g0245(.A(KEYINPUT15), .B(G87), .Z(new_n446));
  NAND3_X1  g0246(.A1(new_n446), .A2(G33), .A3(new_n220), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n255), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n448), .B1(new_n349), .B2(new_n269), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n271), .A2(G77), .A3(new_n272), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(G200), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n443), .B(new_n452), .C1(new_n453), .C2(new_n442), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n442), .A2(new_n374), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n440), .A2(new_n385), .A3(new_n441), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(new_n451), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  NOR4_X1   g0258(.A1(new_n334), .A2(new_n372), .A3(new_n433), .A4(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(KEYINPUT80), .A2(G41), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT5), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT5), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n462), .B1(KEYINPUT80), .B2(G41), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G45), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(G1), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G274), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n461), .A2(new_n463), .A3(new_n466), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n469), .A2(new_n286), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n468), .B1(new_n470), .B2(G257), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n298), .A2(new_n300), .A3(G250), .A4(G1698), .ZN(new_n472));
  NAND2_X1  g0272(.A1(G33), .A2(G283), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n298), .A2(new_n300), .A3(G244), .A4(new_n302), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT4), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT4), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n347), .A2(new_n477), .A3(G244), .A4(new_n302), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n474), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n305), .B1(new_n479), .B2(KEYINPUT79), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n476), .A2(new_n478), .ZN(new_n481));
  INV_X1    g0281(.A(new_n474), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n481), .A2(KEYINPUT79), .A3(new_n482), .ZN(new_n483));
  OAI211_X1 g0283(.A(KEYINPUT81), .B(new_n471), .C1(new_n480), .C2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n481), .A2(new_n482), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT79), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n479), .A2(KEYINPUT79), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(new_n305), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(KEYINPUT81), .B1(new_n490), .B2(new_n471), .ZN(new_n491));
  OAI21_X1  g0291(.A(G190), .B1(new_n485), .B2(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n255), .B(new_n267), .C1(G1), .C2(new_n256), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G97), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n337), .A2(new_n248), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n257), .A2(new_n349), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT6), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n247), .A2(new_n249), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n246), .A2(KEYINPUT6), .A3(G97), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(KEYINPUT78), .B(new_n499), .C1(new_n503), .C2(new_n220), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n412), .B(G107), .C1(new_n413), .C2(new_n411), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT78), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n220), .B1(new_n501), .B2(new_n502), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n506), .B1(new_n507), .B2(new_n498), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n504), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n497), .B1(new_n509), .B2(new_n270), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n471), .B1(new_n480), .B2(new_n483), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n511), .B1(G200), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT81), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n515), .A2(new_n385), .A3(new_n484), .ZN(new_n516));
  INV_X1    g0316(.A(new_n471), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n286), .B1(new_n486), .B2(new_n487), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n517), .B1(new_n518), .B2(new_n489), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n510), .B1(new_n519), .B2(new_n374), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n492), .A2(new_n513), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT88), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n298), .A2(new_n300), .A3(G257), .A4(G1698), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT87), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n347), .A2(KEYINPUT87), .A3(G257), .A4(G1698), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G294), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n347), .A2(G250), .A3(new_n302), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n525), .A2(new_n526), .A3(new_n527), .A4(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n305), .ZN(new_n530));
  INV_X1    g0330(.A(new_n468), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n470), .A2(G264), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n522), .B1(new_n533), .B2(new_n374), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n529), .A2(new_n305), .B1(G264), .B2(new_n470), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n535), .A2(KEYINPUT88), .A3(G179), .A4(new_n531), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n533), .A2(G169), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n220), .A2(new_n347), .A3(G87), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT22), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT22), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n220), .A2(new_n347), .A3(new_n541), .A4(G87), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  OR2_X1    g0343(.A1(KEYINPUT83), .A2(G116), .ZN(new_n544));
  NAND2_X1  g0344(.A1(KEYINPUT83), .A2(G116), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n544), .A2(G33), .A3(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT23), .ZN(new_n547));
  AOI21_X1  g0347(.A(G20), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(KEYINPUT23), .A2(G107), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n246), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n549), .B1(new_n220), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n543), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT24), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n543), .A2(KEYINPUT24), .A3(new_n552), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n555), .A2(new_n270), .A3(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT25), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n267), .B2(G107), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n337), .A2(KEYINPUT25), .A3(new_n246), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n494), .A2(G107), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n538), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n533), .A2(G200), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n535), .A2(G190), .A3(new_n531), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n557), .A2(new_n564), .A3(new_n561), .A4(new_n565), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT86), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n298), .A2(new_n300), .A3(G264), .A4(G1698), .ZN(new_n569));
  INV_X1    g0369(.A(G303), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n569), .B1(new_n570), .B2(new_n347), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n347), .A2(G257), .A3(new_n302), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n305), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n469), .A2(G270), .A3(new_n286), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n531), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G169), .ZN(new_n576));
  INV_X1    g0376(.A(G116), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n577), .B1(new_n266), .B2(G33), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n265), .A2(new_n255), .A3(new_n268), .A4(new_n578), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n265), .A2(new_n268), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n544), .A2(new_n545), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n579), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT20), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n270), .B1(new_n582), .B2(new_n216), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n473), .B1(new_n248), .B2(G33), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n444), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n584), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n255), .B1(G20), .B2(new_n581), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n589), .B(KEYINPUT20), .C1(new_n444), .C2(new_n586), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n583), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n568), .B1(new_n576), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT21), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT21), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n568), .B(new_n594), .C1(new_n576), .C2(new_n591), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n575), .A2(G200), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n596), .B(new_n591), .C1(new_n332), .C2(new_n575), .ZN(new_n597));
  INV_X1    g0397(.A(new_n591), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n575), .A2(new_n374), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n593), .A2(new_n595), .A3(new_n597), .A4(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n580), .A2(new_n446), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT19), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(KEYINPUT84), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT84), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT19), .ZN(new_n606));
  AND2_X1   g0406(.A1(G33), .A2(G97), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n604), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n220), .ZN(new_n609));
  INV_X1    g0409(.A(G87), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n610), .A2(KEYINPUT85), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n610), .A2(KEYINPUT85), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n248), .B(new_n246), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n220), .A2(G33), .A3(G97), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n604), .A2(new_n606), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n220), .A2(new_n347), .A3(G68), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n614), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n602), .B1(new_n619), .B2(new_n270), .ZN(new_n620));
  INV_X1    g0420(.A(new_n446), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n620), .B1(new_n621), .B2(new_n493), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n286), .B(G250), .C1(G1), .C2(new_n465), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n467), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n298), .A2(new_n300), .A3(G244), .A4(G1698), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n546), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n298), .A2(new_n300), .A3(G238), .A4(new_n302), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT82), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n347), .A2(KEYINPUT82), .A3(G238), .A4(new_n302), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n627), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n625), .B1(new_n632), .B2(new_n286), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n385), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n630), .A2(new_n631), .ZN(new_n635));
  INV_X1    g0435(.A(new_n627), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n286), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n637), .A2(new_n624), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n374), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n622), .A2(new_n634), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n638), .A2(G190), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n493), .A2(new_n610), .ZN(new_n642));
  AOI211_X1 g0442(.A(new_n642), .B(new_n602), .C1(new_n619), .C2(new_n270), .ZN(new_n643));
  OAI21_X1  g0443(.A(G200), .B1(new_n637), .B2(new_n624), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n641), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n640), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n601), .A2(new_n646), .ZN(new_n647));
  AND4_X1   g0447(.A1(new_n459), .A2(new_n521), .A3(new_n567), .A4(new_n647), .ZN(G372));
  INV_X1    g0448(.A(new_n457), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n329), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n432), .A2(new_n333), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n422), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n371), .A2(KEYINPUT10), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(new_n653), .A3(new_n368), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n654), .A2(new_n360), .ZN(new_n655));
  INV_X1    g0455(.A(new_n642), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n644), .A2(KEYINPUT89), .A3(new_n656), .A4(new_n620), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n641), .ZN(new_n658));
  AOI21_X1  g0458(.A(KEYINPUT89), .B1(new_n643), .B2(new_n644), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n566), .B(new_n640), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n592), .A2(KEYINPUT21), .B1(new_n598), .B2(new_n599), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n563), .A2(new_n595), .A3(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n521), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n516), .A2(new_n520), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n658), .A2(new_n659), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n665), .A2(new_n666), .A3(new_n640), .A4(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n516), .A2(new_n520), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT26), .B1(new_n669), .B2(new_n646), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n664), .A2(new_n640), .A3(new_n668), .A4(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n459), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n655), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g0473(.A(new_n673), .B(KEYINPUT90), .Z(G369));
  NAND2_X1  g0474(.A1(new_n662), .A2(new_n595), .ZN(new_n675));
  INV_X1    g0475(.A(G13), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n444), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n266), .ZN(new_n678));
  OAI21_X1  g0478(.A(G213), .B1(new_n678), .B2(KEYINPUT27), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT91), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n678), .A2(KEYINPUT91), .A3(KEYINPUT27), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n679), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(new_n591), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n675), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n601), .B2(new_n686), .ZN(new_n688));
  XOR2_X1   g0488(.A(new_n688), .B(KEYINPUT92), .Z(new_n689));
  INV_X1    g0489(.A(new_n685), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n562), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n567), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n563), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n690), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n689), .A2(G330), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n675), .A2(new_n685), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n567), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n563), .B2(new_n690), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n696), .A2(new_n701), .ZN(G399));
  NOR2_X1   g0502(.A1(new_n613), .A2(G116), .ZN(new_n703));
  INV_X1    g0503(.A(new_n226), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G41), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n703), .A2(new_n706), .A3(G1), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n224), .B2(new_n706), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT28), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT95), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT29), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n671), .A2(new_n711), .A3(new_n685), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n665), .A2(new_n666), .A3(new_n645), .A4(new_n640), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n640), .B1(new_n658), .B2(new_n659), .ZN(new_n714));
  OAI21_X1  g0514(.A(KEYINPUT26), .B1(new_n669), .B2(new_n714), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n664), .A2(new_n640), .A3(new_n713), .A4(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n711), .B1(new_n716), .B2(new_n685), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n712), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n485), .A2(new_n491), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n530), .A2(new_n532), .ZN(new_n722));
  OAI21_X1  g0522(.A(KEYINPUT93), .B1(new_n722), .B2(new_n633), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT93), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n638), .A2(new_n724), .A3(new_n535), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n723), .A2(new_n725), .A3(new_n599), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n720), .B1(new_n721), .B2(new_n726), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n723), .A2(new_n725), .A3(new_n599), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n728), .B(KEYINPUT30), .C1(new_n491), .C2(new_n485), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n633), .B(KEYINPUT94), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n533), .A2(new_n374), .A3(new_n575), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(new_n512), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n727), .A2(new_n729), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n690), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n647), .A2(new_n521), .A3(new_n567), .A4(new_n685), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n734), .A2(new_n735), .A3(KEYINPUT31), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT31), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n733), .A2(new_n737), .A3(new_n690), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n736), .A2(G330), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n710), .B1(new_n719), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n718), .A2(KEYINPUT95), .A3(new_n739), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n709), .B1(new_n743), .B2(G1), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n744), .B(KEYINPUT96), .Z(G364));
  AOI21_X1  g0545(.A(new_n266), .B1(new_n677), .B2(G45), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n705), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G13), .A2(G33), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n688), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n221), .B1(G20), .B2(new_n385), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n704), .A2(new_n405), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT97), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n759), .A2(G355), .B1(new_n577), .B2(new_n704), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n704), .A2(new_n347), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n762), .B1(new_n465), .B2(new_n225), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(new_n244), .B2(new_n465), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n757), .B1(new_n760), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n220), .A2(G190), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n374), .A2(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G311), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR4_X1   g0570(.A1(new_n216), .A2(new_n332), .A3(new_n453), .A4(G179), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n347), .B1(new_n771), .B2(G303), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n374), .A2(new_n332), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n444), .A2(new_n453), .A3(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G322), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G179), .A2(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G190), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n444), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G294), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n772), .B1(new_n774), .B2(new_n775), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n766), .A2(new_n776), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n770), .B(new_n781), .C1(G329), .C2(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n444), .A2(G200), .A3(new_n773), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT99), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G326), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n766), .A2(G200), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(G179), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n374), .ZN(new_n790));
  XOR2_X1   g0590(.A(KEYINPUT100), .B(G317), .Z(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT33), .ZN(new_n792));
  AOI22_X1  g0592(.A1(G283), .A2(new_n789), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n784), .A2(new_n787), .A3(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(KEYINPUT101), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  INV_X1    g0597(.A(new_n789), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n246), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(G68), .B2(new_n790), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n782), .A2(new_n400), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT32), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n774), .B(KEYINPUT98), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G58), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n778), .A2(G97), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n611), .A2(new_n612), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n405), .B1(new_n771), .B2(new_n806), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n805), .B(new_n807), .C1(new_n201), .C2(new_n785), .ZN(new_n808));
  INV_X1    g0608(.A(new_n768), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n808), .B1(G77), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n800), .A2(new_n802), .A3(new_n804), .A4(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n796), .A2(new_n797), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n765), .B1(new_n812), .B2(new_n755), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n749), .B1(new_n754), .B2(new_n813), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n689), .A2(G330), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n689), .A2(G330), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n814), .B1(new_n817), .B2(new_n749), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT102), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G396));
  NAND2_X1  g0620(.A1(new_n671), .A2(new_n685), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n457), .A2(new_n690), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n454), .B1(new_n452), .B2(new_n685), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n822), .B1(new_n823), .B2(new_n457), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n821), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n740), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n826), .A2(KEYINPUT105), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n826), .A2(KEYINPUT105), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n825), .A2(new_n740), .ZN(new_n829));
  NOR4_X1   g0629(.A1(new_n827), .A2(new_n828), .A3(new_n748), .A4(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n755), .A2(new_n750), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n748), .B1(G77), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n785), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n809), .A2(G159), .B1(new_n834), .B2(G137), .ZN(new_n835));
  INV_X1    g0635(.A(G150), .ZN(new_n836));
  INV_X1    g0636(.A(new_n790), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(G143), .B2(new_n803), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT34), .Z(new_n840));
  NAND2_X1  g0640(.A1(new_n789), .A2(G68), .ZN(new_n841));
  INV_X1    g0641(.A(new_n771), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n347), .B1(new_n842), .B2(new_n201), .C1(new_n779), .C2(new_n202), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(G132), .B2(new_n783), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n840), .A2(new_n841), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n805), .B1(new_n780), .B2(new_n774), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT103), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n405), .B1(new_n842), .B2(new_n246), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n782), .A2(new_n769), .B1(new_n785), .B2(new_n570), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n848), .B(new_n849), .C1(new_n582), .C2(new_n809), .ZN(new_n850));
  INV_X1    g0650(.A(G283), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n850), .B1(new_n610), .B2(new_n798), .C1(new_n851), .C2(new_n837), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n845), .B1(new_n847), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n833), .B1(new_n853), .B2(new_n755), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n824), .B2(new_n751), .ZN(new_n855));
  XOR2_X1   g0655(.A(new_n855), .B(KEYINPUT104), .Z(new_n856));
  NOR2_X1   g0656(.A1(new_n830), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(G384));
  NOR2_X1   g0658(.A1(new_n677), .A2(new_n266), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n459), .A2(G330), .A3(new_n736), .A4(new_n738), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n410), .B1(new_n403), .B2(new_n407), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n392), .B1(new_n409), .B2(new_n861), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n382), .A2(new_n389), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n684), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n430), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT37), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT109), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI211_X1 g0668(.A(KEYINPUT109), .B(KEYINPUT37), .C1(new_n863), .C2(new_n865), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n417), .A2(new_n684), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n870), .A2(new_n430), .ZN(new_n871));
  XOR2_X1   g0671(.A(KEYINPUT110), .B(KEYINPUT37), .Z(new_n872));
  NAND3_X1  g0672(.A1(new_n871), .A2(new_n418), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n868), .A2(new_n869), .A3(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT108), .ZN(new_n875));
  INV_X1    g0675(.A(new_n864), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n433), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n420), .A2(new_n421), .B1(new_n431), .B2(new_n429), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT108), .B1(new_n878), .B2(new_n864), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n874), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT38), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n874), .A2(new_n877), .A3(new_n879), .A4(KEYINPUT38), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n690), .A2(new_n279), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n327), .B1(new_n317), .B2(new_n323), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n333), .B(new_n885), .C1(new_n886), .C2(new_n280), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT106), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n329), .B2(new_n690), .ZN(new_n889));
  NOR4_X1   g0689(.A1(new_n886), .A2(KEYINPUT106), .A3(new_n280), .A4(new_n685), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT107), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(KEYINPUT107), .B(new_n887), .C1(new_n889), .C2(new_n890), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n736), .A2(new_n738), .A3(new_n824), .ZN(new_n896));
  NAND2_X1  g0696(.A1(KEYINPUT112), .A2(KEYINPUT40), .ZN(new_n897));
  AND4_X1   g0697(.A1(new_n884), .A2(new_n895), .A3(new_n896), .A4(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n896), .A2(new_n895), .A3(new_n897), .ZN(new_n899));
  XNOR2_X1  g0699(.A(KEYINPUT111), .B(KEYINPUT38), .ZN(new_n900));
  INV_X1    g0700(.A(new_n873), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n872), .B1(new_n871), .B2(new_n418), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n878), .A2(new_n870), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n900), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n883), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n736), .A2(new_n738), .A3(new_n824), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n893), .B2(new_n894), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT112), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n899), .B(new_n906), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n898), .B1(new_n910), .B2(KEYINPUT40), .ZN(new_n911));
  INV_X1    g0711(.A(G330), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n860), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n459), .A2(new_n736), .A3(new_n738), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n913), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n459), .B1(new_n712), .B2(new_n717), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n655), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n915), .B(new_n917), .Z(new_n918));
  INV_X1    g0718(.A(KEYINPUT39), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(new_n882), .B2(new_n883), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n906), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n919), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n330), .A2(new_n690), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n422), .A2(new_n684), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n671), .A2(new_n685), .A3(new_n824), .ZN(new_n928));
  INV_X1    g0728(.A(new_n822), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n895), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n927), .B1(new_n933), .B2(new_n884), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n926), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n859), .B1(new_n918), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n936), .B2(new_n918), .ZN(new_n938));
  INV_X1    g0738(.A(new_n503), .ZN(new_n939));
  OAI211_X1 g0739(.A(G116), .B(new_n222), .C1(new_n939), .C2(KEYINPUT35), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(KEYINPUT35), .B2(new_n939), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n941), .B(KEYINPUT36), .Z(new_n942));
  NAND2_X1  g0742(.A1(new_n393), .A2(G77), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n240), .B1(new_n224), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(G1), .A3(new_n676), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n938), .A2(new_n942), .A3(new_n945), .ZN(G367));
  NOR2_X1   g0746(.A1(new_n238), .A2(new_n762), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n756), .B1(new_n226), .B2(new_n621), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n748), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI221_X1 g0749(.A(new_n347), .B1(new_n842), .B2(new_n202), .C1(new_n779), .C2(new_n203), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(G50), .B2(new_n809), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n786), .A2(G143), .ZN(new_n952));
  INV_X1    g0752(.A(new_n774), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n783), .A2(G137), .B1(new_n953), .B2(G150), .ZN(new_n954));
  AOI22_X1  g0754(.A1(G77), .A2(new_n789), .B1(new_n790), .B2(G159), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n951), .A2(new_n952), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n798), .A2(new_n248), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n347), .B(new_n957), .C1(G317), .C2(new_n783), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT114), .Z(new_n959));
  NAND3_X1  g0759(.A1(new_n771), .A2(KEYINPUT46), .A3(G116), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n842), .A2(new_n581), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n960), .B1(new_n779), .B2(new_n246), .C1(new_n961), .C2(KEYINPUT46), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(G283), .B2(new_n809), .ZN(new_n963));
  XNOR2_X1  g0763(.A(KEYINPUT113), .B(G311), .ZN(new_n964));
  AOI22_X1  g0764(.A1(G303), .A2(new_n803), .B1(new_n786), .B2(new_n964), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n963), .B(new_n965), .C1(new_n780), .C2(new_n837), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n956), .B1(new_n959), .B2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT47), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n755), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(new_n967), .B2(new_n968), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n949), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n685), .A2(new_n643), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n667), .A2(new_n640), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n640), .B2(new_n974), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n972), .B1(new_n753), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n521), .B1(new_n510), .B2(new_n685), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n665), .A2(new_n690), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n700), .A2(new_n981), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT44), .Z(new_n983));
  NOR2_X1   g0783(.A1(new_n700), .A2(new_n981), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT45), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n696), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n986), .B(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n699), .B1(new_n695), .B2(new_n698), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n816), .B(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n743), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n705), .B(KEYINPUT41), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n747), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n698), .A2(new_n521), .A3(new_n567), .A4(new_n663), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n994), .A2(KEYINPUT42), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n492), .A2(new_n513), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n693), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n690), .B1(new_n997), .B2(new_n669), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(new_n994), .B2(KEYINPUT42), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n995), .A2(new_n999), .B1(KEYINPUT43), .B2(new_n976), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n696), .A2(new_n981), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1002), .B(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n977), .B1(new_n993), .B2(new_n1004), .ZN(G387));
  INV_X1    g0805(.A(new_n743), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1006), .A2(new_n990), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1007), .A2(new_n706), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n990), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1008), .B1(new_n743), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n692), .A2(new_n694), .A3(new_n752), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n703), .B(KEYINPUT115), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n465), .B1(new_n203), .B2(new_n349), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n341), .A2(new_n201), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1013), .B1(new_n1014), .B2(KEYINPUT50), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(KEYINPUT50), .B2(new_n1014), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n761), .B1(new_n1012), .B2(new_n1016), .C1(new_n465), .C2(new_n235), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n703), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n759), .A2(new_n1018), .B1(new_n246), .B2(new_n704), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n757), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n779), .A2(new_n621), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n405), .B1(new_n771), .B2(G77), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1022), .B(new_n1023), .C1(new_n768), .C2(new_n203), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G50), .A2(new_n953), .B1(new_n834), .B2(G159), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n836), .B2(new_n782), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n837), .A2(new_n390), .ZN(new_n1027));
  NOR4_X1   g0827(.A1(new_n1024), .A2(new_n1026), .A3(new_n957), .A4(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT116), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n347), .B1(new_n783), .B2(G326), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n786), .A2(G322), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n803), .A2(G317), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n790), .A2(new_n964), .B1(new_n809), .B2(G303), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT48), .Z(new_n1035));
  OAI22_X1  g0835(.A1(new_n779), .A2(new_n851), .B1(new_n780), .B2(new_n842), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1030), .B1(new_n581), .B2(new_n798), .C1(new_n1037), .C2(KEYINPUT49), .ZN(new_n1038));
  AND2_X1   g0838(.A1(new_n1037), .A2(KEYINPUT49), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1029), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n749), .B(new_n1020), .C1(new_n1040), .C2(new_n755), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n1009), .A2(new_n747), .B1(new_n1011), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1010), .A2(new_n1042), .ZN(G393));
  NOR2_X1   g0843(.A1(new_n252), .A2(new_n762), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n757), .B1(G97), .B2(new_n704), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n749), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n405), .B1(new_n842), .B2(new_n851), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n582), .B2(new_n778), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n780), .B2(new_n768), .C1(new_n775), .C2(new_n782), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n799), .B(new_n1050), .C1(G303), .C2(new_n790), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G311), .A2(new_n953), .B1(new_n834), .B2(G317), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT52), .Z(new_n1053));
  AOI21_X1  g0853(.A(new_n405), .B1(new_n771), .B2(G68), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1054), .B1(new_n768), .B2(new_n390), .C1(new_n349), .C2(new_n779), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n201), .A2(new_n837), .B1(new_n798), .B2(new_n610), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1055), .B(new_n1056), .C1(G143), .C2(new_n783), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n836), .A2(new_n785), .B1(new_n774), .B2(new_n400), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT51), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n1051), .A2(new_n1053), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1047), .B1(new_n970), .B2(new_n1060), .C1(new_n980), .C2(new_n753), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n986), .B(new_n696), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1007), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n705), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1007), .A2(new_n1062), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1061), .B1(new_n746), .B2(new_n988), .C1(new_n1064), .C2(new_n1065), .ZN(G390));
  OAI21_X1  g0866(.A(new_n748), .B1(new_n341), .B2(new_n832), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n785), .A2(new_n851), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n405), .B1(new_n842), .B2(new_n610), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(G77), .C2(new_n778), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n768), .A2(new_n248), .B1(new_n774), .B2(new_n577), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(G294), .B2(new_n783), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n790), .A2(G107), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1070), .A2(new_n841), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  NOR3_X1   g0874(.A1(new_n842), .A2(KEYINPUT53), .A3(new_n836), .ZN(new_n1075));
  OAI21_X1  g0875(.A(KEYINPUT53), .B1(new_n842), .B2(new_n836), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n400), .B2(new_n779), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1075), .B(new_n1077), .C1(G137), .C2(new_n790), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n347), .B1(new_n798), .B2(new_n201), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT120), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  XOR2_X1   g0881(.A(KEYINPUT54), .B(G143), .Z(new_n1082));
  AND2_X1   g0882(.A1(new_n809), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G125), .B2(new_n783), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G128), .A2(new_n834), .B1(new_n953), .B2(G132), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1078), .A2(new_n1081), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1074), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1067), .B1(new_n1088), .B2(new_n755), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n924), .B2(new_n751), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n896), .A2(new_n895), .A3(G330), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n925), .B1(new_n930), .B2(new_n895), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n906), .A2(KEYINPUT39), .ZN(new_n1094));
  NOR3_X1   g0894(.A1(new_n1093), .A2(new_n920), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n925), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n906), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n823), .A2(new_n457), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n716), .A2(new_n685), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n929), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1097), .B1(new_n895), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1092), .B1(new_n1095), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1100), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1096), .B(new_n906), .C1(new_n1103), .C2(new_n932), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1091), .B(new_n1104), .C1(new_n924), .C2(new_n1093), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1090), .B1(new_n1106), .B2(new_n746), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n916), .A2(new_n655), .A3(new_n860), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(KEYINPUT117), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT117), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n916), .A2(new_n1110), .A3(new_n655), .A4(new_n860), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n736), .A2(G330), .A3(new_n738), .A4(new_n824), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1112), .A2(new_n893), .A3(new_n894), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n1091), .A2(new_n1103), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n931), .B1(new_n1091), .B2(new_n1113), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1109), .B(new_n1111), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(KEYINPUT118), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1091), .A2(new_n1103), .A3(new_n1113), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n908), .A2(G330), .B1(new_n932), .B2(new_n1112), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1118), .B1(new_n1119), .B2(new_n931), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT118), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1120), .A2(new_n1121), .A3(new_n1111), .A4(new_n1109), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1117), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1123), .A2(KEYINPUT119), .A3(new_n1106), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1117), .A2(new_n1122), .A3(KEYINPUT119), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1106), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n706), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1107), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(G378));
  OAI21_X1  g0929(.A(new_n684), .B1(new_n345), .B2(new_n340), .ZN(new_n1130));
  XOR2_X1   g0930(.A(new_n372), .B(new_n1130), .Z(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1131), .B(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n911), .B2(new_n912), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1133), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT40), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n896), .A2(new_n895), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n922), .B1(new_n1137), .B2(KEYINPUT112), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1136), .B1(new_n1138), .B2(new_n899), .ZN(new_n1139));
  OAI211_X1 g0939(.A(G330), .B(new_n1135), .C1(new_n1139), .C2(new_n898), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1134), .A2(new_n936), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n936), .B1(new_n1134), .B2(new_n1140), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1106), .B1(new_n1117), .B2(new_n1122), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n1141), .A2(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT57), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n706), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1134), .A2(new_n1140), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n935), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1134), .A2(new_n1140), .A3(new_n936), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1148), .A2(new_n1152), .A3(KEYINPUT57), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1147), .A2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n747), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1135), .A2(new_n751), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n347), .A2(G41), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n201), .B1(G33), .B2(G41), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n790), .A2(G97), .B1(new_n809), .B2(new_n446), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT121), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n774), .A2(new_n246), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1157), .B1(new_n842), .B2(new_n349), .C1(new_n782), .C2(new_n851), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1162), .B(new_n1163), .C1(G58), .C2(new_n789), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n834), .A2(G116), .B1(G68), .B2(new_n778), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT122), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1161), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1159), .B1(new_n1168), .B2(KEYINPUT58), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n809), .A2(G137), .B1(new_n834), .B2(G125), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n953), .A2(G128), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n778), .A2(G150), .B1(new_n771), .B2(new_n1082), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G132), .B2(new_n790), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n789), .A2(G159), .ZN(new_n1177));
  AOI211_X1 g0977(.A(G33), .B(G41), .C1(new_n783), .C2(G124), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1169), .B1(KEYINPUT58), .B2(new_n1168), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n755), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1182), .B(new_n748), .C1(G50), .C2(new_n832), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1156), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1155), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1154), .A2(new_n1187), .ZN(G375));
  NAND2_X1  g0988(.A1(new_n1120), .A2(new_n747), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n749), .B1(new_n203), .B2(new_n831), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n783), .A2(G303), .B1(new_n834), .B2(G294), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n246), .B2(new_n768), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n347), .B(new_n1021), .C1(G97), .C2(new_n771), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n789), .A2(G77), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n953), .A2(G283), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1192), .B(new_n1196), .C1(new_n582), .C2(new_n790), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n1197), .A2(KEYINPUT123), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n347), .B1(new_n842), .B2(new_n400), .C1(new_n779), .C2(new_n201), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G128), .B2(new_n783), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n803), .A2(G137), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n809), .A2(G150), .B1(new_n834), .B2(G132), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G58), .A2(new_n789), .B1(new_n790), .B2(new_n1082), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1198), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(KEYINPUT123), .B2(new_n1197), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1190), .B1(new_n1206), .B2(new_n970), .C1(new_n751), .C2(new_n895), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1189), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n1144), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1117), .A2(new_n1122), .A3(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n992), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1209), .B1(new_n1212), .B2(new_n1213), .ZN(G381));
  OR2_X1    g1014(.A1(G387), .A2(G390), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1010), .A2(new_n819), .A3(new_n1042), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(new_n1215), .A2(G384), .A3(G381), .A4(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1186), .B1(new_n1147), .B2(new_n1153), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1217), .A2(new_n1128), .A3(new_n1218), .ZN(G407));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1128), .ZN(new_n1220));
  OAI211_X1 g1020(.A(G407), .B(G213), .C1(G343), .C2(new_n1220), .ZN(G409));
  NAND2_X1  g1021(.A1(G393), .A2(G396), .ZN(new_n1222));
  AND2_X1   g1022(.A1(new_n1222), .A2(new_n1216), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(G387), .A2(G390), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1215), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1215), .A2(new_n1224), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1223), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT61), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT60), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n706), .B1(new_n1211), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(KEYINPUT60), .B2(new_n1212), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n857), .B1(new_n1233), .B2(new_n1208), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1212), .A2(KEYINPUT60), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n1231), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1236), .A2(G384), .A3(new_n1209), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1234), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(G343), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1239), .A2(G213), .A3(G2897), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1229), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(G213), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT124), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1150), .A2(KEYINPUT124), .A3(new_n1151), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n1245), .A3(new_n747), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1148), .A2(new_n1152), .A3(new_n992), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1246), .A2(new_n1247), .A3(new_n1128), .A4(new_n1185), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1242), .B(new_n1248), .C1(new_n1218), .C2(new_n1128), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT125), .ZN(new_n1250));
  AOI21_X1  g1050(.A(G384), .B1(new_n1236), .B2(new_n1209), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n857), .B(new_n1208), .C1(new_n1235), .C2(new_n1231), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1250), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1234), .A2(new_n1237), .A3(KEYINPUT125), .ZN(new_n1254));
  AND3_X1   g1054(.A1(new_n1253), .A2(new_n1254), .A3(new_n1240), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1241), .B1(new_n1249), .B2(new_n1255), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1257));
  OAI21_X1  g1057(.A(KEYINPUT62), .B1(new_n1249), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1256), .A2(new_n1258), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1249), .A2(new_n1257), .A3(KEYINPUT62), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1225), .B(new_n1228), .C1(new_n1259), .C2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT63), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n1249), .B2(new_n1257), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1256), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(G375), .A2(G378), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1248), .A2(new_n1242), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1265), .A2(new_n1266), .A3(KEYINPUT63), .A4(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1228), .A2(new_n1225), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT126), .B1(new_n1264), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1256), .A2(new_n1263), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT126), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1272), .A2(new_n1273), .A3(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1261), .B1(new_n1271), .B2(new_n1275), .ZN(G405));
  AOI21_X1  g1076(.A(new_n1238), .B1(new_n1265), .B2(new_n1220), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(KEYINPUT127), .B2(new_n1257), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1267), .A2(KEYINPUT127), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1279), .A2(new_n1220), .A3(new_n1265), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(new_n1269), .ZN(G402));
endmodule


