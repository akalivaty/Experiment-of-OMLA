//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 1 1 1 1 0 1 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 0 0 1 1 0 1 1 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1232, new_n1233, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1321, new_n1322;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OR2_X1    g0009(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n211));
  NAND3_X1  g0011(.A1(new_n210), .A2(G50), .A3(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT65), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n225));
  INV_X1    g0025(.A(G87), .ZN(new_n226));
  INV_X1    g0026(.A(G250), .ZN(new_n227));
  INV_X1    g0027(.A(G97), .ZN(new_n228));
  INV_X1    g0028(.A(G257), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n225), .B1(new_n226), .B2(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT66), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n206), .B1(new_n224), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n209), .B(new_n217), .C1(new_n232), .C2(KEYINPUT1), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(G226), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT68), .ZN(new_n245));
  XOR2_X1   g0045(.A(G58), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT81), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT81), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n254), .B1(new_n257), .B2(KEYINPUT3), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n258), .A2(KEYINPUT22), .A3(new_n215), .A4(G87), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT22), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n253), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n215), .A2(G87), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n260), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G116), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n257), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(new_n215), .ZN(new_n268));
  INV_X1    g0068(.A(G107), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G20), .ZN(new_n270));
  OR2_X1    g0070(.A1(new_n270), .A2(KEYINPUT23), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n270), .A2(KEYINPUT23), .B1(KEYINPUT87), .B2(KEYINPUT24), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n259), .A2(new_n265), .A3(new_n268), .A4(new_n273), .ZN(new_n274));
  OR2_X1    g0074(.A1(KEYINPUT87), .A2(KEYINPUT24), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n274), .B(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n214), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(new_n278), .B(KEYINPUT70), .ZN(new_n280));
  INV_X1    g0080(.A(G13), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(G1), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G20), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n280), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n285), .B1(G1), .B2(new_n261), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(new_n269), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n284), .A2(new_n269), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n288), .B(KEYINPUT25), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n291));
  INV_X1    g0091(.A(G45), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(G1), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT5), .B(G41), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n291), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G264), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT88), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT88), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n295), .A2(new_n298), .A3(G264), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G274), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n291), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n302), .A2(KEYINPUT85), .A3(new_n293), .A4(new_n294), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT85), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n294), .A2(new_n293), .ZN(new_n305));
  INV_X1    g0105(.A(G41), .ZN(new_n306));
  OAI211_X1 g0106(.A(G1), .B(G13), .C1(new_n261), .C2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G274), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n304), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  OR2_X1    g0110(.A1(KEYINPUT81), .A2(G33), .ZN(new_n311));
  NAND2_X1  g0111(.A1(KEYINPUT81), .A2(G33), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(KEYINPUT3), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n253), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n229), .A2(G1698), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(G250), .B2(G1698), .ZN(new_n316));
  INV_X1    g0116(.A(G294), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n314), .A2(new_n316), .B1(new_n317), .B2(new_n257), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n291), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n300), .A2(new_n310), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G179), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n319), .A2(new_n310), .A3(new_n296), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G169), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n279), .A2(new_n290), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n279), .A2(new_n290), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  OR3_X1    g0127(.A1(new_n323), .A2(KEYINPUT89), .A3(G190), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT89), .B1(new_n323), .B2(G190), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n328), .B(new_n329), .C1(G200), .C2(new_n321), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n325), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(G20), .A2(G33), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n332), .ZN(new_n333));
  XNOR2_X1  g0133(.A(KEYINPUT8), .B(G58), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT71), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT71), .ZN(new_n336));
  INV_X1    g0136(.A(G58), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT8), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n215), .A2(G33), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n333), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n341), .A2(new_n280), .B1(new_n202), .B2(new_n284), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT70), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n278), .B(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n283), .ZN(new_n345));
  INV_X1    g0145(.A(G1), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G20), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G50), .ZN(new_n348));
  XOR2_X1   g0148(.A(new_n348), .B(KEYINPUT72), .Z(new_n349));
  OAI21_X1  g0149(.A(new_n342), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT9), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n350), .A2(new_n351), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n253), .A2(new_n262), .ZN(new_n354));
  NOR2_X1   g0154(.A1(G222), .A2(G1698), .ZN(new_n355));
  INV_X1    g0155(.A(G1698), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n356), .A2(G223), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n354), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n358), .B(new_n291), .C1(G77), .C2(new_n354), .ZN(new_n359));
  AOI21_X1  g0159(.A(G1), .B1(new_n306), .B2(new_n292), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n302), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G226), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n291), .A2(new_n360), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n359), .B(new_n361), .C1(new_n362), .C2(new_n364), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n365), .B(KEYINPUT69), .ZN(new_n366));
  INV_X1    g0166(.A(G200), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI211_X1 g0168(.A(new_n352), .B(new_n353), .C1(new_n368), .C2(KEYINPUT76), .ZN(new_n369));
  XOR2_X1   g0169(.A(new_n365), .B(KEYINPUT69), .Z(new_n370));
  INV_X1    g0170(.A(G190), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT76), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(new_n367), .B2(new_n366), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT10), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT10), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n369), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G169), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n370), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G179), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n366), .A2(new_n381), .ZN(new_n382));
  AND3_X1   g0182(.A1(new_n380), .A2(new_n382), .A3(new_n350), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n378), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT80), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n332), .A2(G50), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n387), .B(KEYINPUT79), .ZN(new_n388));
  OAI22_X1  g0188(.A1(new_n340), .A2(new_n221), .B1(new_n215), .B2(G68), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n280), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT11), .ZN(new_n391));
  OR2_X1    g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n390), .A2(new_n391), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT12), .B1(new_n283), .B2(G68), .ZN(new_n394));
  OR3_X1    g0194(.A1(new_n283), .A2(KEYINPUT12), .A3(G68), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n284), .A2(new_n278), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n219), .B1(new_n346), .B2(G20), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n394), .A2(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n392), .A2(new_n393), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(G232), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G1698), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n354), .B(new_n402), .C1(G226), .C2(G1698), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G97), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n307), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n361), .B1(new_n364), .B2(new_n220), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT13), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n406), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT13), .B1(new_n405), .B2(new_n407), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(G169), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT14), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n379), .B1(new_n410), .B2(new_n411), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT14), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT78), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n410), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n406), .A2(new_n408), .A3(KEYINPUT78), .A4(new_n409), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(new_n421), .A3(new_n411), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n422), .A2(new_n381), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n400), .B1(new_n418), .B2(new_n423), .ZN(new_n424));
  AND3_X1   g0224(.A1(new_n412), .A2(KEYINPUT77), .A3(G200), .ZN(new_n425));
  AOI21_X1  g0225(.A(KEYINPUT77), .B1(new_n412), .B2(G200), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n400), .B1(new_n422), .B2(new_n371), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n386), .B1(new_n424), .B2(new_n429), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n427), .A2(new_n428), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n414), .B(new_n417), .C1(new_n381), .C2(new_n422), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n399), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n431), .A2(new_n433), .A3(KEYINPUT80), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n283), .A2(KEYINPUT75), .A3(G77), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT75), .B1(new_n283), .B2(G77), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n221), .B1(new_n346), .B2(G20), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n436), .A2(new_n437), .B1(new_n396), .B2(new_n438), .ZN(new_n439));
  XNOR2_X1  g0239(.A(KEYINPUT15), .B(G87), .ZN(new_n440));
  OAI22_X1  g0240(.A1(new_n440), .A2(new_n340), .B1(new_n215), .B2(new_n221), .ZN(new_n441));
  XOR2_X1   g0241(.A(new_n334), .B(KEYINPUT74), .Z(new_n442));
  AOI21_X1  g0242(.A(new_n441), .B1(new_n442), .B2(new_n332), .ZN(new_n443));
  INV_X1    g0243(.A(new_n278), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n439), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n354), .A2(G232), .A3(new_n356), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n269), .B2(new_n354), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n263), .A2(new_n220), .A3(new_n356), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n291), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT73), .ZN(new_n450));
  AOI22_X1  g0250(.A1(G244), .A2(new_n363), .B1(new_n302), .B2(new_n360), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n450), .B1(new_n449), .B2(new_n451), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n445), .B1(new_n454), .B2(G200), .ZN(new_n455));
  OAI21_X1  g0255(.A(G190), .B1(new_n452), .B2(new_n453), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n454), .A2(new_n379), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n381), .B1(new_n452), .B2(new_n453), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(new_n445), .A3(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n430), .A2(new_n434), .A3(new_n457), .A4(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT16), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT7), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(G20), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT3), .B1(new_n311), .B2(new_n312), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT83), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n466), .B1(new_n252), .B2(G33), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n261), .A2(KEYINPUT83), .A3(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n464), .B1(new_n465), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n463), .B1(new_n354), .B2(G20), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n219), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g0272(.A1(G58), .A2(G68), .ZN(new_n473));
  OAI21_X1  g0273(.A(G20), .B1(new_n473), .B2(new_n201), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n332), .A2(G159), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n462), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT82), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n474), .A2(new_n478), .A3(new_n475), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n478), .B1(new_n474), .B2(new_n475), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR3_X1   g0281(.A1(new_n255), .A2(new_n256), .A3(new_n252), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n463), .B(new_n215), .C1(new_n482), .C2(new_n254), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G68), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n463), .B1(new_n314), .B2(new_n215), .ZN(new_n485));
  OAI211_X1 g0285(.A(KEYINPUT16), .B(new_n481), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n477), .A2(new_n486), .A3(new_n278), .ZN(new_n487));
  INV_X1    g0287(.A(new_n339), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n347), .ZN(new_n489));
  OAI22_X1  g0289(.A1(new_n489), .A2(new_n345), .B1(new_n283), .B2(new_n488), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n361), .B1(new_n364), .B2(new_n401), .ZN(new_n493));
  NOR2_X1   g0293(.A1(G223), .A2(G1698), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n494), .B1(new_n362), .B2(G1698), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(new_n313), .A3(new_n253), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G87), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n307), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(G169), .B1(new_n493), .B2(new_n498), .ZN(new_n499));
  AOI22_X1  g0299(.A1(G232), .A2(new_n363), .B1(new_n302), .B2(new_n360), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n496), .A2(new_n497), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n500), .B(G179), .C1(new_n501), .C2(new_n307), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n492), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT18), .ZN(new_n505));
  XNOR2_X1  g0305(.A(new_n504), .B(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n367), .B1(new_n493), .B2(new_n498), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n500), .B(new_n371), .C1(new_n501), .C2(new_n307), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n487), .A2(new_n491), .A3(new_n509), .ZN(new_n510));
  XNOR2_X1  g0310(.A(new_n510), .B(KEYINPUT17), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n385), .A2(new_n461), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT21), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n266), .B1(new_n346), .B2(G33), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n396), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n282), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n215), .A2(G116), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n516), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G283), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n521), .B(new_n215), .C1(G33), .C2(new_n228), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n522), .A2(new_n519), .A3(new_n278), .ZN(new_n523));
  XNOR2_X1  g0323(.A(new_n523), .B(KEYINPUT20), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G169), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n295), .A2(G270), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n310), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n229), .A2(new_n356), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n258), .B(new_n530), .C1(G264), .C2(new_n356), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n263), .A2(G303), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n307), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n514), .B1(new_n527), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(G190), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n536), .B(new_n525), .C1(new_n367), .C2(new_n534), .ZN(new_n537));
  INV_X1    g0337(.A(new_n534), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n538), .A2(KEYINPUT21), .A3(G169), .A4(new_n526), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n529), .A2(new_n533), .A3(new_n381), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n526), .ZN(new_n541));
  AND4_X1   g0341(.A1(new_n535), .A2(new_n537), .A3(new_n539), .A4(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT7), .B1(new_n263), .B2(new_n215), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n467), .B(new_n468), .C1(new_n257), .C2(KEYINPUT3), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n543), .B1(new_n544), .B2(new_n464), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n545), .A2(new_n269), .ZN(new_n546));
  XNOR2_X1  g0346(.A(G97), .B(G107), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT6), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR3_X1   g0349(.A1(new_n548), .A2(new_n228), .A3(G107), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n332), .ZN(new_n552));
  OAI22_X1  g0352(.A1(new_n551), .A2(new_n215), .B1(new_n221), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n278), .B1(new_n546), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n345), .B1(new_n346), .B2(G33), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G97), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n284), .A2(new_n228), .ZN(new_n557));
  XNOR2_X1  g0357(.A(new_n557), .B(KEYINPUT84), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n554), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n354), .A2(KEYINPUT4), .A3(G244), .A4(new_n356), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n354), .A2(G250), .A3(G1698), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n560), .A2(new_n521), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n258), .A2(G244), .A3(new_n356), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT4), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n307), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n295), .A2(G257), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n310), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n379), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n560), .A2(new_n521), .A3(new_n561), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n570), .B1(new_n564), .B2(new_n563), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n310), .B(new_n567), .C1(new_n571), .C2(new_n307), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n559), .B(new_n569), .C1(G179), .C2(new_n572), .ZN(new_n573));
  OR2_X1    g0373(.A1(new_n545), .A2(new_n269), .ZN(new_n574));
  OR2_X1    g0374(.A1(new_n549), .A2(new_n550), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n575), .A2(G20), .B1(G77), .B2(new_n332), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n444), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n558), .B1(new_n286), .B2(new_n228), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n566), .A2(new_n568), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(G190), .ZN(new_n581));
  OAI21_X1  g0381(.A(G200), .B1(new_n566), .B2(new_n568), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n579), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n258), .A2(new_n215), .A3(G68), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n340), .A2(new_n228), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n584), .B1(KEYINPUT19), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n587));
  NOR2_X1   g0387(.A1(G97), .A2(G107), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n215), .A2(new_n587), .B1(new_n588), .B2(new_n226), .ZN(new_n589));
  XNOR2_X1  g0389(.A(new_n589), .B(KEYINPUT86), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n278), .B1(new_n586), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n284), .A2(new_n440), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n591), .B(new_n592), .C1(new_n286), .C2(new_n440), .ZN(new_n593));
  NOR2_X1   g0393(.A1(G238), .A2(G1698), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n594), .B1(new_n222), .B2(G1698), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n267), .B1(new_n258), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n596), .A2(new_n307), .ZN(new_n597));
  INV_X1    g0397(.A(new_n293), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n307), .A2(new_n598), .A3(G250), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n308), .B2(new_n598), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n379), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n381), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n593), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n602), .A2(G200), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n591), .A2(new_n592), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n555), .A2(G87), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n601), .A2(G190), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n606), .A2(new_n607), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  AND4_X1   g0410(.A1(new_n573), .A2(new_n583), .A3(new_n605), .A4(new_n610), .ZN(new_n611));
  AND4_X1   g0411(.A1(new_n331), .A2(new_n513), .A3(new_n542), .A4(new_n611), .ZN(G372));
  NAND2_X1  g0412(.A1(new_n327), .A2(new_n330), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n539), .A2(new_n541), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n535), .ZN(new_n616));
  OAI21_X1  g0416(.A(KEYINPUT90), .B1(new_n616), .B2(new_n325), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n322), .A2(new_n324), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n326), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT90), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n619), .A2(new_n615), .A3(new_n620), .A4(new_n535), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n614), .A2(new_n617), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n605), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n610), .A2(new_n605), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n573), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(KEYINPUT26), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT26), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n628), .B1(new_n624), .B2(new_n573), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n623), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n622), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n513), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n632), .B(KEYINPUT91), .ZN(new_n633));
  INV_X1    g0433(.A(new_n460), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n424), .B1(new_n431), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n511), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n506), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n383), .B1(new_n637), .B2(new_n378), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n633), .A2(new_n638), .ZN(G369));
  OR3_X1    g0439(.A1(new_n517), .A2(KEYINPUT27), .A3(G20), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT27), .B1(new_n517), .B2(G20), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(G213), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(G343), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n525), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n616), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n542), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n647), .B1(new_n648), .B2(new_n646), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(G330), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n331), .B1(new_n327), .B2(new_n645), .ZN(new_n653));
  OAI21_X1  g0453(.A(KEYINPUT92), .B1(new_n619), .B2(new_n645), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT92), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n325), .A2(new_n655), .A3(new_n644), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n652), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n616), .A2(new_n645), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n660), .B1(new_n653), .B2(new_n657), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n619), .A2(new_n644), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n659), .A2(new_n663), .ZN(G399));
  INV_X1    g0464(.A(new_n207), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(G41), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n588), .A2(new_n226), .A3(new_n266), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n667), .A2(G1), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n212), .B2(new_n667), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT93), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT28), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n300), .A2(new_n319), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n674), .A2(new_n601), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n675), .A2(KEYINPUT30), .A3(new_n540), .A4(new_n580), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n540), .A2(new_n580), .A3(new_n601), .A4(new_n674), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT30), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n534), .A2(G179), .A3(new_n601), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT94), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n321), .B2(new_n580), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n572), .A2(new_n320), .A3(KEYINPUT94), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n682), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n644), .B1(new_n680), .B2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT31), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT95), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n331), .A2(new_n611), .A3(new_n542), .A4(new_n645), .ZN(new_n691));
  OAI211_X1 g0491(.A(KEYINPUT31), .B(new_n644), .C1(new_n680), .C2(new_n686), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n651), .B1(new_n690), .B2(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n644), .B1(new_n622), .B2(new_n630), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n695), .A2(KEYINPUT29), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n614), .B1(new_n325), .B2(new_n616), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n644), .B1(new_n697), .B2(new_n630), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(KEYINPUT29), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n694), .B1(new_n696), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n673), .B1(new_n700), .B2(G1), .ZN(G364));
  NAND2_X1  g0501(.A1(new_n650), .A2(new_n651), .ZN(new_n702));
  INV_X1    g0502(.A(new_n652), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n281), .A2(G20), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G45), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n705), .A2(KEYINPUT96), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(KEYINPUT96), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(G1), .A3(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(new_n666), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n702), .A2(new_n703), .A3(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(G13), .A2(G33), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G20), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n214), .B1(G20), .B2(new_n379), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT98), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n247), .A2(new_n292), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n258), .A2(new_n665), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n720), .B1(new_n292), .B2(new_n213), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n718), .B1(KEYINPUT97), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(KEYINPUT97), .B2(new_n721), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n354), .A2(new_n207), .ZN(new_n724));
  INV_X1    g0524(.A(G355), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n726), .B1(new_n266), .B2(new_n665), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n717), .B1(new_n723), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n215), .A2(new_n381), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n730), .A2(KEYINPUT99), .ZN(new_n731));
  AOI21_X1  g0531(.A(G200), .B1(new_n730), .B2(KEYINPUT99), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n731), .A2(new_n371), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n381), .A2(new_n367), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT100), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G190), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  AOI22_X1  g0538(.A1(new_n734), .A2(G77), .B1(new_n738), .B2(G97), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n731), .A2(G190), .A3(new_n732), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n739), .B1(new_n337), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n215), .A2(G179), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(new_n371), .A3(G200), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n269), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n729), .A2(G200), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G190), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n371), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n746), .A2(G68), .B1(new_n747), .B2(G50), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n742), .A2(G190), .A3(G200), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n748), .B1(new_n226), .B2(new_n749), .ZN(new_n750));
  NOR4_X1   g0550(.A1(new_n741), .A2(new_n263), .A3(new_n744), .A4(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n736), .A2(G20), .A3(new_n371), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n752), .A2(KEYINPUT101), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(KEYINPUT101), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AND3_X1   g0556(.A1(new_n756), .A2(KEYINPUT32), .A3(G159), .ZN(new_n757));
  AOI21_X1  g0557(.A(KEYINPUT32), .B1(new_n756), .B2(G159), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n751), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT102), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n756), .A2(G329), .ZN(new_n762));
  INV_X1    g0562(.A(new_n749), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n354), .B1(new_n763), .B2(G303), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(KEYINPUT103), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n765), .B1(G311), .B2(new_n734), .ZN(new_n766));
  INV_X1    g0566(.A(new_n740), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n767), .A2(G322), .B1(new_n738), .B2(G294), .ZN(new_n768));
  NOR2_X1   g0568(.A1(KEYINPUT33), .A2(G317), .ZN(new_n769));
  AND2_X1   g0569(.A1(KEYINPUT33), .A2(G317), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n746), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n747), .A2(G326), .ZN(new_n772));
  INV_X1    g0572(.A(G283), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n771), .B(new_n772), .C1(new_n773), .C2(new_n743), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n774), .B1(KEYINPUT103), .B2(new_n764), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n762), .A2(new_n766), .A3(new_n768), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n759), .A2(new_n760), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n761), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n710), .B(new_n728), .C1(new_n778), .C2(new_n715), .ZN(new_n779));
  INV_X1    g0579(.A(new_n714), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n779), .B1(new_n649), .B2(new_n780), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n711), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(G396));
  NAND2_X1  g0583(.A1(new_n634), .A2(new_n645), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n455), .A2(new_n456), .B1(new_n445), .B2(new_n644), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n784), .B1(new_n785), .B2(new_n634), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n695), .B(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n694), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n709), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(new_n789), .B2(new_n788), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n715), .A2(new_n712), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n709), .B1(G77), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n756), .A2(G311), .ZN(new_n795));
  INV_X1    g0595(.A(new_n747), .ZN(new_n796));
  INV_X1    g0596(.A(G303), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n263), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n746), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n799), .A2(new_n773), .B1(new_n226), .B2(new_n743), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n798), .B(new_n800), .C1(G107), .C2(new_n763), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n767), .A2(G294), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n734), .A2(G116), .B1(new_n738), .B2(G97), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n795), .A2(new_n801), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n746), .A2(G150), .B1(new_n747), .B2(G137), .ZN(new_n805));
  INV_X1    g0605(.A(G143), .ZN(new_n806));
  INV_X1    g0606(.A(G159), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n805), .B1(new_n740), .B2(new_n806), .C1(new_n807), .C2(new_n733), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT34), .Z(new_n809));
  NOR2_X1   g0609(.A1(new_n743), .A2(new_n219), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n314), .B(new_n810), .C1(G50), .C2(new_n763), .ZN(new_n811));
  INV_X1    g0611(.A(new_n738), .ZN(new_n812));
  INV_X1    g0612(.A(G132), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n811), .B1(new_n337), .B2(new_n812), .C1(new_n755), .C2(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n804), .B1(new_n809), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n794), .B1(new_n815), .B2(new_n715), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n787), .B2(new_n713), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n791), .A2(new_n817), .ZN(G384));
  OR2_X1    g0618(.A1(new_n575), .A2(KEYINPUT35), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n575), .A2(KEYINPUT35), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n819), .A2(G116), .A3(new_n216), .A4(new_n820), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n821), .B(KEYINPUT36), .Z(new_n822));
  OR3_X1    g0622(.A1(new_n212), .A2(new_n221), .A3(new_n473), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n202), .A2(G68), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n346), .B(G13), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n433), .A2(new_n644), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT37), .ZN(new_n828));
  INV_X1    g0628(.A(new_n476), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n545), .B2(new_n219), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n444), .B1(new_n830), .B2(new_n462), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n490), .B1(new_n831), .B2(new_n486), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n828), .B(new_n510), .C1(new_n832), .C2(new_n642), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT106), .ZN(new_n834));
  AOI221_X4 g0634(.A(new_n834), .B1(new_n499), .B2(new_n502), .C1(new_n487), .C2(new_n491), .ZN(new_n835));
  AOI21_X1  g0635(.A(KEYINPUT106), .B1(new_n492), .B2(new_n503), .ZN(new_n836));
  OR3_X1    g0636(.A1(new_n833), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT105), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n484), .A2(new_n485), .ZN(new_n839));
  INV_X1    g0639(.A(new_n481), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n462), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(KEYINPUT7), .B1(new_n258), .B2(G20), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n842), .A2(G68), .A3(new_n483), .ZN(new_n843));
  NOR3_X1   g0643(.A1(new_n479), .A2(new_n480), .A3(new_n462), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n344), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n490), .B1(new_n841), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n510), .B1(new_n846), .B2(new_n642), .ZN(new_n847));
  INV_X1    g0647(.A(new_n503), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n838), .B(KEYINPUT37), .C1(new_n847), .C2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n486), .A2(new_n280), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT16), .B1(new_n843), .B2(new_n481), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n491), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n503), .ZN(new_n855));
  INV_X1    g0655(.A(new_n642), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n855), .A2(new_n857), .A3(new_n510), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n838), .B1(new_n858), .B2(KEYINPUT37), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n837), .B1(new_n851), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT107), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n857), .B1(new_n506), .B2(new_n511), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n837), .B(KEYINPUT107), .C1(new_n851), .C2(new_n859), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n862), .A2(KEYINPUT38), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT39), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT38), .ZN(new_n868));
  NOR3_X1   g0668(.A1(new_n833), .A2(new_n835), .A3(new_n836), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n492), .A2(new_n856), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n504), .A2(new_n870), .A3(new_n510), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n869), .B1(KEYINPUT37), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n870), .B1(new_n506), .B2(new_n511), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n868), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n866), .A2(new_n867), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n865), .A2(new_n864), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT37), .B1(new_n847), .B2(new_n849), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT105), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n850), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT107), .B1(new_n879), .B2(new_n837), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n868), .B1(new_n876), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n867), .B1(new_n881), .B2(new_n866), .ZN(new_n882));
  NOR3_X1   g0682(.A1(new_n875), .A2(new_n882), .A3(KEYINPUT108), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT108), .ZN(new_n884));
  NOR3_X1   g0684(.A1(new_n876), .A2(new_n880), .A3(new_n868), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n869), .B1(new_n878), .B2(new_n850), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n863), .B1(new_n886), .B2(KEYINPUT107), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT38), .B1(new_n887), .B2(new_n862), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT39), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n866), .A2(new_n867), .A3(new_n874), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n884), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n827), .B1(new_n883), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n506), .A2(new_n856), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n399), .A2(new_n644), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n894), .B(KEYINPUT104), .Z(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n424), .B2(new_n429), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n431), .A2(new_n433), .A3(new_n895), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n631), .A2(new_n787), .A3(new_n645), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n900), .B1(new_n901), .B2(new_n784), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n881), .A2(new_n866), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n893), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n892), .A2(KEYINPUT109), .A3(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT109), .ZN(new_n906));
  INV_X1    g0706(.A(new_n827), .ZN(new_n907));
  OAI21_X1  g0707(.A(KEYINPUT108), .B1(new_n875), .B2(new_n882), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n889), .A2(new_n884), .A3(new_n890), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n904), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n906), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n905), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n696), .A2(new_n513), .A3(new_n699), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n914), .A2(new_n638), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n913), .B(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT110), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n692), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n684), .A2(new_n685), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n681), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n920), .A2(new_n679), .A3(new_n676), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n921), .A2(KEYINPUT110), .A3(KEYINPUT31), .A4(new_n644), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n918), .A2(new_n922), .A3(new_n691), .A4(new_n689), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n786), .B1(new_n897), .B2(new_n898), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT40), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n903), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n923), .A2(new_n924), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n866), .B2(new_n874), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n928), .B1(new_n925), .B2(new_n930), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n513), .A2(new_n923), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n651), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n932), .B2(new_n931), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n916), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n346), .B2(new_n704), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n916), .A2(new_n934), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n826), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n938), .B(KEYINPUT111), .Z(G367));
  OAI211_X1 g0739(.A(new_n583), .B(new_n573), .C1(new_n579), .C2(new_n645), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n940), .A2(KEYINPUT113), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(KEYINPUT113), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n941), .B(new_n942), .C1(new_n573), .C2(new_n645), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n661), .A2(KEYINPUT42), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n661), .A2(new_n943), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT42), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n619), .B1(new_n941), .B2(new_n942), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n948), .A2(new_n626), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n944), .A2(new_n947), .B1(new_n645), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n607), .A2(new_n608), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n644), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n625), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n623), .A2(new_n951), .A3(new_n644), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT112), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n950), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n959), .B1(KEYINPUT43), .B2(new_n955), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n960), .B1(new_n950), .B2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n943), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n963), .B1(new_n659), .B2(new_n964), .ZN(new_n965));
  OR3_X1    g0765(.A1(new_n963), .A2(new_n659), .A3(new_n964), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n666), .B(KEYINPUT41), .Z(new_n967));
  INV_X1    g0767(.A(new_n661), .ZN(new_n968));
  INV_X1    g0768(.A(new_n662), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n968), .A2(new_n969), .A3(new_n943), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT45), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n663), .A2(KEYINPUT45), .A3(new_n943), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT44), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n663), .B2(new_n943), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n964), .B(KEYINPUT44), .C1(new_n661), .C2(new_n662), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n974), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n659), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n658), .B1(new_n616), .B2(new_n645), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n703), .B1(new_n982), .B2(new_n661), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NOR3_X1   g0784(.A1(new_n703), .A2(new_n982), .A3(new_n661), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n974), .A2(new_n978), .A3(new_n659), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n981), .A2(new_n700), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n967), .B1(new_n988), .B2(new_n700), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n965), .B(new_n966), .C1(new_n989), .C2(new_n708), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n743), .A2(new_n228), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G311), .B2(new_n747), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n992), .B(new_n314), .C1(new_n317), .C2(new_n799), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n749), .A2(new_n266), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT46), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n993), .B(new_n995), .C1(new_n756), .C2(G317), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n767), .A2(G303), .B1(new_n738), .B2(G107), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n996), .B(new_n997), .C1(new_n773), .C2(new_n733), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n756), .A2(G137), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n354), .B1(new_n796), .B2(new_n806), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n799), .A2(new_n807), .B1(new_n221), .B2(new_n743), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n1000), .B(new_n1001), .C1(G58), .C2(new_n763), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n734), .A2(G50), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n767), .A2(G150), .B1(new_n738), .B2(G68), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n999), .A2(new_n1002), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n998), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT47), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n715), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n242), .A2(new_n719), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n440), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n715), .B(new_n714), .C1(new_n665), .C2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n710), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1008), .B(new_n1012), .C1(new_n780), .C2(new_n955), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n990), .A2(new_n1013), .ZN(G387));
  OAI22_X1  g0814(.A1(new_n724), .A2(new_n669), .B1(G107), .B2(new_n207), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n239), .A2(new_n292), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n442), .A2(new_n202), .ZN(new_n1018));
  XOR2_X1   g0818(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n1019));
  XNOR2_X1  g0819(.A(new_n1018), .B(new_n1019), .ZN(new_n1020));
  AOI211_X1 g0820(.A(G45), .B(new_n668), .C1(G68), .C2(G77), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1017), .A2(KEYINPUT114), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT114), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n720), .B1(new_n1016), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1015), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n709), .B1(new_n1025), .B2(new_n717), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n314), .B(new_n991), .C1(G77), .C2(new_n763), .ZN(new_n1027));
  INV_X1    g0827(.A(G150), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1027), .B1(new_n755), .B2(new_n1028), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT116), .Z(new_n1030));
  NOR2_X1   g0830(.A1(new_n812), .A2(new_n440), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n488), .A2(new_n746), .B1(G159), .B2(new_n747), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G50), .A2(new_n767), .B1(new_n734), .B2(G68), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1030), .A2(new_n1032), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT117), .Z(new_n1036));
  AOI22_X1  g0836(.A1(new_n746), .A2(G311), .B1(new_n747), .B2(G322), .ZN(new_n1037));
  INV_X1    g0837(.A(G317), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1037), .B1(new_n740), .B2(new_n1038), .C1(new_n797), .C2(new_n733), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT48), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n738), .A2(G283), .B1(G294), .B2(new_n763), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT49), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n314), .B1(new_n266), .B2(new_n743), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n756), .B2(G326), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1046), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1036), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1026), .B1(new_n1051), .B2(new_n715), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n658), .B2(new_n780), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT118), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n708), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n986), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n700), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n666), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n986), .A2(new_n700), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1054), .B1(new_n1055), .B2(new_n1056), .C1(new_n1058), .C2(new_n1059), .ZN(G393));
  INV_X1    g0860(.A(new_n987), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n659), .B1(new_n974), .B2(new_n978), .ZN(new_n1062));
  NOR3_X1   g0862(.A1(new_n1061), .A2(new_n1055), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n964), .A2(new_n714), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n716), .B1(new_n228), .B2(new_n207), .C1(new_n720), .C2(new_n250), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n709), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n740), .A2(new_n807), .B1(new_n1028), .B2(new_n796), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT51), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n756), .A2(G143), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n812), .A2(new_n221), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n258), .B1(new_n226), .B2(new_n743), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n799), .A2(new_n202), .B1(new_n219), .B2(new_n749), .ZN(new_n1072));
  NOR3_X1   g0872(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n734), .A2(new_n442), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1068), .A2(new_n1069), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n767), .A2(G311), .B1(G317), .B2(new_n747), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT52), .Z(new_n1077));
  AOI22_X1  g0877(.A1(new_n738), .A2(G116), .B1(G303), .B2(new_n746), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1077), .B(new_n1078), .C1(new_n317), .C2(new_n733), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n354), .B(new_n744), .C1(G283), .C2(new_n763), .ZN(new_n1080));
  INV_X1    g0880(.A(G322), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1080), .B1(new_n755), .B2(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT119), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1075), .B1(new_n1079), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1066), .B1(new_n1084), .B2(new_n715), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1063), .B1(new_n1064), .B2(new_n1085), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n1061), .A2(new_n1062), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1087), .A2(new_n988), .A3(new_n666), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1086), .A2(new_n1088), .ZN(G390));
  INV_X1    g0889(.A(new_n784), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n695), .B2(new_n787), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n907), .B1(new_n1091), .B2(new_n900), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n908), .A2(new_n909), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n866), .A2(new_n874), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n785), .A2(new_n634), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1090), .B1(new_n698), .B2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n907), .B(new_n1094), .C1(new_n1096), .C2(new_n900), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n694), .A2(new_n787), .A3(new_n899), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1093), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n923), .A2(G330), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n924), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n908), .A2(new_n909), .A3(new_n712), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n709), .B1(new_n488), .B2(new_n793), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n810), .B1(G107), .B2(new_n746), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n773), .B2(new_n796), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n354), .B(new_n1108), .C1(G87), .C2(new_n763), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n317), .B2(new_n755), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1070), .B1(G97), .B2(new_n734), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n266), .B2(new_n740), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n756), .A2(G125), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n738), .A2(G159), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n263), .B1(new_n747), .B2(G128), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n743), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n746), .A2(G137), .B1(new_n1116), .B2(G50), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .A4(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n749), .A2(new_n1028), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT53), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(KEYINPUT54), .B(G143), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1120), .B1(new_n813), .B2(new_n740), .C1(new_n733), .C2(new_n1121), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1110), .A2(new_n1112), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1106), .B1(new_n1123), .B2(new_n715), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1104), .A2(new_n708), .B1(new_n1105), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n513), .A2(new_n1101), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n914), .A2(new_n638), .A3(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n923), .A2(new_n787), .A3(G330), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n900), .ZN(new_n1129));
  OR2_X1    g0929(.A1(new_n1129), .A2(KEYINPUT120), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(KEYINPUT120), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1130), .A2(new_n1096), .A3(new_n1098), .A4(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1091), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n899), .B1(new_n694), .B2(new_n787), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1102), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1133), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1127), .B1(new_n1132), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1093), .A2(new_n1097), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n1135), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1141), .A2(new_n1099), .A3(new_n1137), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1139), .A2(new_n666), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1125), .A2(new_n1143), .ZN(G378));
  NAND2_X1  g0944(.A1(new_n350), .A2(new_n856), .ZN(new_n1145));
  XOR2_X1   g0945(.A(new_n1145), .B(KEYINPUT55), .Z(new_n1146));
  NAND2_X1  g0946(.A1(new_n385), .A2(new_n1146), .ZN(new_n1147));
  XOR2_X1   g0947(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n1148));
  AOI21_X1  g0948(.A(new_n383), .B1(new_n375), .B2(new_n377), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1146), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1147), .A2(new_n1148), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1148), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n383), .B(new_n1146), .C1(new_n375), .C2(new_n377), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1153), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1152), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n929), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n925), .B1(new_n1094), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n926), .B1(new_n866), .B2(new_n881), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1157), .B(G330), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1157), .B1(new_n931), .B2(G330), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n1164), .A2(new_n905), .A3(new_n912), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1164), .B1(new_n912), .B2(new_n905), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n708), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1157), .A2(new_n712), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n793), .A2(G50), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n756), .A2(G283), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n734), .A2(new_n1010), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n767), .A2(G107), .B1(new_n738), .B2(G68), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n799), .A2(new_n228), .B1(new_n221), .B2(new_n749), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n796), .A2(new_n266), .B1(new_n337), .B2(new_n743), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n314), .A2(new_n306), .ZN(new_n1175));
  NOR3_X1   g0975(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .A4(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT58), .ZN(new_n1178));
  AOI21_X1  g0978(.A(G50), .B1(new_n261), .B2(new_n306), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1177), .A2(new_n1178), .B1(new_n1175), .B2(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n746), .A2(G132), .B1(new_n747), .B2(G125), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n749), .B2(new_n1121), .ZN(new_n1182));
  INV_X1    g0982(.A(G128), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n812), .A2(new_n1028), .B1(new_n1183), .B2(new_n740), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1182), .B(new_n1184), .C1(G137), .C2(new_n734), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT59), .Z(new_n1186));
  AOI211_X1 g0986(.A(G33), .B(G41), .C1(new_n1116), .C2(G159), .ZN(new_n1187));
  INV_X1    g0987(.A(G124), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1187), .B1(new_n755), .B2(new_n1188), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n1189), .B(KEYINPUT121), .Z(new_n1190));
  OAI221_X1 g0990(.A(new_n1180), .B1(new_n1178), .B2(new_n1177), .C1(new_n1186), .C2(new_n1190), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n710), .B(new_n1169), .C1(new_n1191), .C2(new_n715), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1168), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1167), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1163), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n1161), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT109), .B1(new_n892), .B2(new_n904), .ZN(new_n1197));
  NOR3_X1   g0997(.A1(new_n910), .A2(new_n906), .A3(new_n911), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1196), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1164), .A2(new_n905), .A3(new_n912), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1127), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1199), .A2(new_n1200), .B1(new_n1142), .B2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n667), .B1(new_n1202), .B2(KEYINPUT57), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT57), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1132), .A2(new_n1136), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1127), .B1(new_n1104), .B2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1204), .B1(new_n1205), .B2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1194), .B1(new_n1203), .B2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(G375));
  NAND2_X1  g1010(.A1(new_n747), .A2(G132), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1211), .B1(new_n807), .B2(new_n749), .C1(new_n799), .C2(new_n1121), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n314), .B(new_n1212), .C1(G58), .C2(new_n1116), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n1183), .B2(new_n755), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n767), .A2(G137), .B1(new_n738), .B2(G50), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1028), .B2(new_n733), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1032), .B1(new_n269), .B2(new_n733), .C1(new_n773), .C2(new_n740), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n796), .A2(new_n317), .B1(new_n228), .B2(new_n749), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G116), .B2(new_n746), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n354), .B1(new_n1116), .B2(G77), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1219), .B(new_n1220), .C1(new_n755), .C2(new_n797), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n1214), .A2(new_n1216), .B1(new_n1217), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n715), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n710), .B1(new_n219), .B2(new_n792), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(new_n899), .C2(new_n713), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n1206), .B2(new_n708), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n967), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1138), .A2(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1206), .A2(new_n1201), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1227), .B1(new_n1229), .B2(new_n1230), .ZN(G381));
  OR2_X1    g1031(.A1(G393), .A2(G396), .ZN(new_n1232));
  OR4_X1    g1032(.A1(G384), .A2(new_n1232), .A3(G381), .A4(G390), .ZN(new_n1233));
  OR4_X1    g1033(.A1(G387), .A2(G375), .A3(G378), .A4(new_n1233), .ZN(G407));
  INV_X1    g1034(.A(G378), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n643), .A2(G213), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1209), .A2(new_n1235), .A3(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(G407), .A2(G213), .A3(new_n1238), .ZN(G409));
  XNOR2_X1  g1039(.A(G393), .B(new_n782), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n990), .A2(new_n1013), .A3(G390), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(G390), .B1(new_n990), .B2(new_n1013), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1241), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(G390), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(G387), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1247), .A2(new_n1240), .A3(new_n1242), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1245), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT125), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1202), .A2(new_n1228), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1252), .A2(new_n708), .B1(new_n1168), .B2(new_n1192), .ZN(new_n1253));
  AOI21_X1  g1053(.A(G378), .B1(new_n1251), .B2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n1209), .B2(G378), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1250), .B1(new_n1255), .B2(new_n1237), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1142), .A2(new_n1201), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1252), .A2(KEYINPUT57), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n666), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1202), .A2(KEYINPUT57), .ZN(new_n1260));
  OAI211_X1 g1060(.A(G378), .B(new_n1253), .C1(new_n1259), .C2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1235), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(KEYINPUT125), .A3(new_n1236), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1227), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1138), .A2(KEYINPUT60), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1230), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n666), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1266), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  OR2_X1    g1072(.A1(G384), .A2(KEYINPUT123), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G384), .A2(KEYINPUT123), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  OR2_X1    g1075(.A1(new_n1272), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1271), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1227), .B(new_n1273), .C1(new_n1277), .C2(new_n1269), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1276), .A2(KEYINPUT62), .A3(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1256), .A2(new_n1265), .A3(new_n1280), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(new_n1236), .A3(new_n1264), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT62), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1281), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1237), .A2(G2897), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1278), .B(new_n1287), .C1(new_n1272), .C2(new_n1275), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT125), .B1(new_n1264), .B2(new_n1236), .ZN(new_n1292));
  AOI211_X1 g1092(.A(new_n1250), .B(new_n1237), .C1(new_n1261), .C2(new_n1263), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1291), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  XNOR2_X1  g1094(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1294), .A2(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1249), .B1(new_n1286), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT127), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT61), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1245), .A2(new_n1300), .A3(new_n1248), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(KEYINPUT124), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT124), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1245), .A2(new_n1248), .A3(new_n1303), .A4(new_n1300), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1302), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1264), .A2(new_n1236), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1305), .B1(new_n1306), .B2(new_n1291), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1256), .A2(KEYINPUT63), .A3(new_n1265), .A4(new_n1282), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT63), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1283), .A2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1307), .A2(new_n1308), .A3(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1298), .A2(new_n1299), .A3(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1249), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1256), .A2(new_n1265), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1295), .B1(new_n1314), .B2(new_n1291), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1281), .A2(new_n1285), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1313), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1307), .A2(new_n1308), .A3(new_n1310), .ZN(new_n1318));
  OAI21_X1  g1118(.A(KEYINPUT127), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1312), .A2(new_n1319), .ZN(G405));
  XNOR2_X1  g1120(.A(new_n1209), .B(G378), .ZN(new_n1321));
  XNOR2_X1  g1121(.A(new_n1321), .B(new_n1282), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(new_n1322), .B(new_n1249), .ZN(G402));
endmodule


