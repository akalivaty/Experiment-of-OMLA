//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 1 1 0 1 1 1 0 1 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n631,
    new_n632, new_n633, new_n634, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n806, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928;
  INV_X1    g000(.A(KEYINPUT79), .ZN(new_n202));
  XNOR2_X1  g001(.A(G155gat), .B(G162gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G141gat), .B(G148gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT2), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n207), .B1(G155gat), .B2(G162gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n206), .B1(KEYINPUT77), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G155gat), .ZN(new_n210));
  INV_X1    g009(.A(G162gat), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT2), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT77), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n204), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n208), .A2(KEYINPUT78), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n208), .A2(KEYINPUT78), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n216), .A2(new_n203), .A3(new_n206), .A4(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n202), .B1(new_n219), .B2(KEYINPUT3), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n215), .A2(KEYINPUT79), .A3(new_n221), .A4(new_n218), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT29), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(G211gat), .B(G218gat), .Z(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT71), .ZN(new_n226));
  XNOR2_X1  g025(.A(G197gat), .B(G204gat), .ZN(new_n227));
  INV_X1    g026(.A(G211gat), .ZN(new_n228));
  INV_X1    g027(.A(G218gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n227), .B1(KEYINPUT22), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n226), .B(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n224), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n231), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n234), .A2(new_n225), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT29), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(new_n234), .B2(new_n225), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n221), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n219), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n233), .A2(new_n239), .B1(G228gat), .B2(G233gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(G228gat), .ZN(new_n242));
  INV_X1    g041(.A(G233gat), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n221), .B1(new_n232), .B2(KEYINPUT29), .ZN(new_n244));
  AOI211_X1 g043(.A(new_n242), .B(new_n243), .C1(new_n244), .C2(new_n219), .ZN(new_n245));
  INV_X1    g044(.A(new_n232), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT81), .B1(new_n223), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NOR3_X1   g047(.A1(new_n223), .A2(KEYINPUT81), .A3(new_n246), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n245), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n250), .A2(KEYINPUT82), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n252));
  OR3_X1    g051(.A1(new_n223), .A2(KEYINPUT81), .A3(new_n246), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n247), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n252), .B1(new_n254), .B2(new_n245), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n241), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G78gat), .B(G106gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT31), .B(G50gat), .ZN(new_n258));
  XOR2_X1   g057(.A(new_n257), .B(new_n258), .Z(new_n259));
  NAND2_X1  g058(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT83), .B(G22gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n250), .A2(KEYINPUT82), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n254), .A2(new_n252), .A3(new_n245), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n259), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(new_n241), .A3(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n260), .A2(new_n261), .A3(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n261), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n265), .B1(new_n264), .B2(new_n241), .ZN(new_n269));
  AOI211_X1 g068(.A(new_n240), .B(new_n259), .C1(new_n262), .C2(new_n263), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(KEYINPUT23), .ZN(new_n273));
  NAND2_X1  g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT65), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT64), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(G183gat), .A2(G190gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT24), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OR2_X1    g079(.A1(G183gat), .A2(G190gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT64), .A4(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT25), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT27), .B(G183gat), .ZN(new_n287));
  INV_X1    g086(.A(G190gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(new_n289), .B(KEYINPUT28), .Z(new_n290));
  XOR2_X1   g089(.A(new_n272), .B(KEYINPUT26), .Z(new_n291));
  OAI211_X1 g090(.A(new_n290), .B(new_n278), .C1(new_n276), .C2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n286), .A2(new_n292), .ZN(new_n293));
  AND2_X1   g092(.A1(G226gat), .A2(G233gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT29), .B1(new_n286), .B2(new_n292), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n295), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(new_n232), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n295), .B(new_n246), .C1(new_n294), .C2(new_n296), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT37), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT38), .ZN(new_n302));
  XOR2_X1   g101(.A(G8gat), .B(G36gat), .Z(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(KEYINPUT72), .ZN(new_n304));
  XOR2_X1   g103(.A(new_n304), .B(KEYINPUT73), .Z(new_n305));
  XNOR2_X1  g104(.A(G64gat), .B(G92gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT37), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n298), .A2(new_n309), .A3(new_n299), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n301), .A2(new_n302), .A3(new_n308), .A4(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n311), .B(KEYINPUT85), .ZN(new_n312));
  XNOR2_X1  g111(.A(G113gat), .B(G120gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT67), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT1), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n315), .B1(new_n314), .B2(new_n313), .ZN(new_n316));
  INV_X1    g115(.A(G127gat), .ZN(new_n317));
  NOR3_X1   g116(.A1(new_n317), .A2(KEYINPUT66), .A3(G134gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(G127gat), .B(G134gat), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n318), .B1(new_n319), .B2(KEYINPUT66), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  OR2_X1    g122(.A1(new_n323), .A2(new_n313), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n325), .A2(new_n219), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(KEYINPUT4), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n220), .A2(new_n222), .ZN(new_n328));
  INV_X1    g127(.A(new_n325), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n329), .B1(KEYINPUT3), .B2(new_n219), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n327), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(G225gat), .A2(G233gat), .ZN(new_n332));
  XOR2_X1   g131(.A(new_n332), .B(KEYINPUT80), .Z(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n331), .A2(KEYINPUT5), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n327), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n330), .A2(new_n328), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(new_n334), .A3(new_n337), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n325), .B(new_n219), .Z(new_n339));
  OAI21_X1  g138(.A(KEYINPUT5), .B1(new_n339), .B2(new_n334), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n335), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G1gat), .B(G29gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n343), .B(KEYINPUT0), .ZN(new_n344));
  XNOR2_X1  g143(.A(G57gat), .B(G85gat), .ZN(new_n345));
  XOR2_X1   g144(.A(new_n344), .B(new_n345), .Z(new_n346));
  NAND2_X1  g145(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT6), .ZN(new_n348));
  INV_X1    g147(.A(new_n346), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n335), .A2(new_n341), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n347), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n301), .A2(new_n308), .A3(new_n310), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT38), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n335), .A2(new_n341), .A3(KEYINPUT6), .A4(new_n349), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n298), .A2(new_n307), .A3(new_n299), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT75), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT75), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n298), .A2(new_n357), .A3(new_n307), .A4(new_n299), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n351), .A2(new_n353), .A3(new_n354), .A4(new_n360), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n267), .B(new_n271), .C1(new_n312), .C2(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n331), .A2(new_n334), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT39), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n349), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n364), .B1(new_n339), .B2(new_n334), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n366), .B(KEYINPUT84), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n365), .B1(new_n363), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT40), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n365), .B(KEYINPUT40), .C1(new_n363), .C2(new_n367), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n370), .A2(new_n350), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT76), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n373), .B1(new_n359), .B2(KEYINPUT30), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT30), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n356), .A2(KEYINPUT76), .A3(new_n375), .A4(new_n358), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  OR3_X1    g176(.A1(new_n355), .A2(KEYINPUT74), .A3(new_n375), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT74), .B1(new_n355), .B2(new_n375), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n378), .A2(new_n379), .B1(new_n308), .B2(new_n300), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n372), .B1(new_n377), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n351), .A2(new_n354), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n377), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  NOR3_X1   g182(.A1(new_n269), .A2(new_n270), .A3(new_n268), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n261), .B1(new_n260), .B2(new_n266), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI22_X1  g185(.A1(new_n362), .A2(new_n381), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n293), .A2(new_n329), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n286), .A2(new_n325), .A3(new_n292), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(G227gat), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n390), .B1(new_n391), .B2(new_n243), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n392), .A2(KEYINPUT70), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT34), .ZN(new_n395));
  XNOR2_X1  g194(.A(G15gat), .B(G43gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(G71gat), .B(G99gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n396), .B(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n391), .A2(new_n243), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n388), .A2(new_n399), .A3(new_n389), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n398), .B1(new_n400), .B2(KEYINPUT32), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT33), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT69), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT69), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n401), .A2(new_n406), .A3(new_n403), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n400), .B(KEYINPUT32), .C1(new_n402), .C2(new_n398), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n395), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n401), .A2(new_n406), .A3(new_n403), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n406), .B1(new_n401), .B2(new_n403), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n395), .B(new_n409), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n394), .B1(new_n410), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT34), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n417), .A2(new_n393), .A3(new_n413), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT36), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n415), .A2(KEYINPUT36), .A3(new_n418), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n387), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT86), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n417), .A2(new_n393), .A3(new_n413), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n393), .B1(new_n417), .B2(new_n413), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n415), .A2(KEYINPUT86), .A3(new_n418), .ZN(new_n429));
  XOR2_X1   g228(.A(KEYINPUT87), .B(KEYINPUT35), .Z(new_n430));
  AND3_X1   g229(.A1(new_n271), .A2(new_n267), .A3(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n428), .A2(new_n429), .A3(new_n383), .A4(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT88), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n383), .A2(new_n419), .A3(new_n386), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n432), .A2(new_n433), .B1(new_n434), .B2(KEYINPUT35), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n271), .A2(new_n267), .A3(new_n430), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n377), .A2(new_n380), .ZN(new_n437));
  INV_X1    g236(.A(new_n382), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n439), .A2(KEYINPUT88), .A3(new_n428), .A4(new_n429), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n424), .B1(new_n435), .B2(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(KEYINPUT91), .B(G29gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(KEYINPUT92), .B(G36gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AND2_X1   g243(.A1(G43gat), .A2(G50gat), .ZN(new_n445));
  NOR2_X1   g244(.A1(G43gat), .A2(G50gat), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT15), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OR3_X1    g246(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n444), .A2(new_n447), .A3(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT93), .B(G43gat), .ZN(new_n452));
  INV_X1    g251(.A(G50gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n445), .A2(KEYINPUT15), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT94), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT94), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n454), .A2(new_n458), .A3(new_n455), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n451), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n448), .A2(KEYINPUT90), .ZN(new_n461));
  OR4_X1    g260(.A1(KEYINPUT90), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n462), .A3(new_n449), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n447), .B1(new_n463), .B2(new_n444), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  OR3_X1    g264(.A1(new_n465), .A2(KEYINPUT95), .A3(KEYINPUT17), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT95), .B1(new_n465), .B2(KEYINPUT17), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G15gat), .B(G22gat), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT96), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT16), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n471), .B1(new_n472), .B2(G1gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n469), .B(KEYINPUT96), .ZN(new_n474));
  INV_X1    g273(.A(G1gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(G8gat), .ZN(new_n478));
  INV_X1    g277(.A(G8gat), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n473), .A2(new_n479), .A3(new_n476), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n481), .B1(KEYINPUT17), .B2(new_n465), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n468), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(G229gat), .A2(G233gat), .ZN(new_n484));
  INV_X1    g283(.A(new_n465), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n483), .A2(KEYINPUT18), .A3(new_n484), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT97), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n468), .A2(new_n482), .B1(new_n485), .B2(new_n481), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT97), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n489), .A2(new_n490), .A3(KEYINPUT18), .A4(new_n484), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n489), .A2(new_n484), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT18), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n481), .B(new_n485), .ZN(new_n495));
  XOR2_X1   g294(.A(new_n484), .B(KEYINPUT13), .Z(new_n496));
  AOI22_X1  g295(.A1(new_n493), .A2(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(G113gat), .B(G141gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(G169gat), .B(G197gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  XOR2_X1   g302(.A(new_n503), .B(KEYINPUT12), .Z(new_n504));
  NAND2_X1  g303(.A1(new_n498), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n504), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n492), .A2(new_n497), .A3(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n465), .A2(KEYINPUT17), .ZN(new_n509));
  NAND2_X1  g308(.A1(G85gat), .A2(G92gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT7), .ZN(new_n511));
  NOR2_X1   g310(.A1(G85gat), .A2(G92gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(G99gat), .A2(G106gat), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n512), .B1(KEYINPUT8), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G99gat), .B(G106gat), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n511), .A2(new_n516), .A3(new_n514), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(KEYINPUT102), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n468), .A2(new_n509), .A3(new_n521), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n511), .A2(new_n516), .A3(new_n514), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n516), .B1(new_n511), .B2(new_n514), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AND2_X1   g324(.A1(G232gat), .A2(G233gat), .ZN(new_n526));
  AOI22_X1  g325(.A1(new_n485), .A2(new_n525), .B1(KEYINPUT41), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G190gat), .B(G218gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n526), .A2(KEYINPUT41), .ZN(new_n531));
  XNOR2_X1  g330(.A(G134gat), .B(G162gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n530), .A2(new_n533), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(G57gat), .B(G64gat), .Z(new_n538));
  NAND2_X1  g337(.A1(G71gat), .A2(G78gat), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT9), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n539), .A2(KEYINPUT98), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT98), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n544), .A2(G71gat), .A3(G78gat), .ZN(new_n545));
  AND2_X1   g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT99), .ZN(new_n547));
  INV_X1    g346(.A(G71gat), .ZN(new_n548));
  INV_X1    g347(.A(G78gat), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT99), .B1(G71gat), .B2(G78gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT100), .B1(new_n546), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n543), .A2(new_n545), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT100), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n554), .A2(new_n555), .A3(new_n551), .A4(new_n550), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n542), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n538), .A2(new_n541), .ZN(new_n558));
  INV_X1    g357(.A(new_n539), .ZN(new_n559));
  NOR2_X1   g358(.A1(G71gat), .A2(G78gat), .ZN(new_n560));
  NOR3_X1   g359(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT21), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G127gat), .B(G155gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n478), .B(new_n480), .C1(new_n563), .C2(new_n562), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT101), .ZN(new_n570));
  XOR2_X1   g369(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G183gat), .B(G211gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n568), .B(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT103), .B1(new_n537), .B2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT103), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n536), .A2(new_n578), .A3(new_n575), .ZN(new_n579));
  NAND2_X1  g378(.A1(G230gat), .A2(G233gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n556), .ZN(new_n582));
  AND2_X1   g381(.A1(new_n550), .A2(new_n551), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n555), .B1(new_n583), .B2(new_n554), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n558), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n561), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n585), .A2(new_n586), .A3(new_n520), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n525), .B1(new_n557), .B2(new_n561), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n587), .A2(new_n588), .A3(KEYINPUT104), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT104), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n562), .A2(new_n590), .A3(new_n520), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT10), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT105), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT105), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n592), .A2(new_n596), .A3(new_n593), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n588), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT10), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n581), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n592), .A2(new_n580), .ZN(new_n602));
  XNOR2_X1  g401(.A(G120gat), .B(G148gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(G176gat), .B(G204gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NOR3_X1   g404(.A1(new_n601), .A2(new_n602), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n605), .B1(new_n601), .B2(new_n602), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n577), .A2(new_n579), .A3(new_n610), .ZN(new_n611));
  NOR3_X1   g410(.A1(new_n441), .A2(new_n508), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(new_n438), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(G1gat), .ZN(G1324gat));
  INV_X1    g413(.A(new_n612), .ZN(new_n615));
  INV_X1    g414(.A(new_n437), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(KEYINPUT16), .B(G8gat), .Z(new_n618));
  AND2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n617), .A2(new_n479), .ZN(new_n620));
  OAI21_X1  g419(.A(KEYINPUT42), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n617), .A2(new_n618), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT42), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n621), .A2(new_n624), .ZN(G1325gat));
  INV_X1    g424(.A(new_n423), .ZN(new_n626));
  OAI21_X1  g425(.A(G15gat), .B1(new_n615), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n428), .A2(new_n429), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n628), .A2(G15gat), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n627), .B1(new_n615), .B2(new_n629), .ZN(G1326gat));
  NOR3_X1   g429(.A1(new_n441), .A2(new_n508), .A3(new_n386), .ZN(new_n631));
  INV_X1    g430(.A(new_n611), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT43), .B(G22gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(G1327gat));
  NAND2_X1  g434(.A1(new_n432), .A2(new_n433), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n434), .A2(KEYINPUT35), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n636), .A2(new_n440), .A3(new_n637), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n387), .A2(new_n423), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n536), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NOR3_X1   g439(.A1(new_n508), .A2(new_n575), .A3(new_n609), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n642), .A2(new_n382), .A3(new_n442), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n643), .B(KEYINPUT45), .Z(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(KEYINPUT44), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT44), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(new_n441), .B2(new_n536), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n641), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n442), .B1(new_n649), .B2(new_n382), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n644), .A2(new_n650), .ZN(G1328gat));
  INV_X1    g450(.A(new_n642), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n616), .A2(new_n443), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(KEYINPUT106), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT106), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n652), .A2(new_n656), .A3(new_n653), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT46), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n443), .B1(new_n649), .B2(new_n616), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n655), .A2(KEYINPUT46), .A3(new_n657), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(G1329gat));
  OAI21_X1  g462(.A(new_n452), .B1(new_n642), .B2(new_n628), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n626), .A2(new_n452), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n664), .B1(new_n649), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(KEYINPUT47), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT47), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n669), .B(new_n664), .C1(new_n649), .C2(new_n666), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(G1330gat));
  INV_X1    g470(.A(new_n386), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n645), .A2(new_n647), .A3(new_n672), .A4(new_n641), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(G50gat), .ZN(new_n674));
  NOR4_X1   g473(.A1(new_n536), .A2(new_n609), .A3(G50gat), .A4(new_n575), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n631), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT48), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1331gat));
  NAND3_X1  g478(.A1(new_n577), .A2(new_n508), .A3(new_n579), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n441), .A2(new_n610), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n438), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g482(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n437), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n685), .B(KEYINPUT107), .Z(new_n686));
  NAND2_X1  g485(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n687), .A2(KEYINPUT108), .ZN(new_n688));
  NOR2_X1   g487(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(KEYINPUT108), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n689), .B1(new_n688), .B2(new_n690), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(G1333gat));
  INV_X1    g492(.A(new_n628), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n681), .A2(new_n548), .A3(new_n694), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n681), .A2(new_n423), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n695), .B1(new_n696), .B2(new_n548), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT50), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1334gat));
  NAND2_X1  g498(.A1(new_n681), .A2(new_n672), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(G78gat), .ZN(G1335gat));
  INV_X1    g500(.A(new_n508), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n702), .A2(new_n575), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(new_n610), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n648), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(G85gat), .B1(new_n706), .B2(new_n382), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n610), .A2(new_n382), .A3(G85gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT110), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT109), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n704), .B1(new_n640), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(KEYINPUT109), .B1(new_n441), .B2(new_n536), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n711), .A2(KEYINPUT51), .A3(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT51), .B1(new_n711), .B2(new_n712), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n709), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n707), .A2(new_n716), .ZN(G1336gat));
  NOR3_X1   g516(.A1(new_n616), .A2(G92gat), .A3(new_n610), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT111), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n638), .A2(new_n639), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n720), .A2(new_n710), .A3(new_n537), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n712), .A2(new_n721), .A3(new_n703), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT51), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n719), .B1(new_n724), .B2(new_n713), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n645), .A2(new_n647), .A3(new_n437), .A4(new_n705), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n726), .A2(G92gat), .ZN(new_n727));
  OAI21_X1  g526(.A(KEYINPUT52), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n718), .B1(new_n714), .B2(new_n715), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT52), .B1(new_n726), .B2(G92gat), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n731), .ZN(G1337gat));
  OAI21_X1  g531(.A(G99gat), .B1(new_n706), .B2(new_n626), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n628), .A2(G99gat), .A3(new_n610), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n734), .B1(new_n714), .B2(new_n715), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(G1338gat));
  NOR3_X1   g535(.A1(new_n386), .A2(G106gat), .A3(new_n610), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n737), .B(KEYINPUT112), .Z(new_n738));
  AOI21_X1  g537(.A(new_n738), .B1(new_n724), .B2(new_n713), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n645), .A2(new_n647), .A3(new_n672), .A4(new_n705), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n740), .A2(G106gat), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT53), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n737), .B1(new_n714), .B2(new_n715), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT53), .B1(new_n740), .B2(G106gat), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n742), .A2(new_n745), .ZN(G1339gat));
  AOI21_X1  g545(.A(new_n596), .B1(new_n592), .B2(new_n593), .ZN(new_n747));
  AOI211_X1 g546(.A(KEYINPUT105), .B(KEYINPUT10), .C1(new_n589), .C2(new_n591), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n600), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT54), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n749), .A2(new_n750), .A3(new_n580), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n580), .B1(new_n599), .B2(KEYINPUT10), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(new_n747), .B2(new_n748), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT54), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n605), .B(new_n751), .C1(new_n601), .C2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT55), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n606), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(KEYINPUT55), .B1(new_n601), .B2(new_n754), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n751), .A2(new_n605), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n758), .A2(KEYINPUT113), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n750), .B1(new_n598), .B2(new_n752), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n749), .A2(new_n580), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n756), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n751), .A2(new_n605), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n761), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n757), .B1(new_n760), .B2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT114), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(KEYINPUT113), .B1(new_n758), .B2(new_n759), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n764), .A2(new_n765), .A3(new_n761), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n772), .A2(KEYINPUT114), .A3(new_n757), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n769), .A2(new_n702), .A3(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT115), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n775), .B1(new_n489), .B2(new_n484), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n495), .B2(new_n496), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n489), .A2(new_n775), .A3(new_n484), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n503), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n609), .A2(new_n507), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n537), .B1(new_n774), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n779), .A2(new_n782), .A3(new_n507), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n779), .B2(new_n507), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n783), .A2(new_n536), .A3(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n785), .A2(new_n769), .A3(new_n773), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n576), .B1(new_n781), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n611), .A2(new_n702), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n438), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n419), .A2(new_n386), .A3(new_n616), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(G113gat), .B1(new_n794), .B2(new_n702), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n672), .B1(new_n788), .B2(new_n790), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n437), .A2(new_n382), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n796), .A2(new_n694), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(G113gat), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n798), .A2(new_n799), .A3(new_n508), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n795), .A2(new_n800), .ZN(G1340gat));
  AOI21_X1  g600(.A(G120gat), .B1(new_n794), .B2(new_n609), .ZN(new_n802));
  INV_X1    g601(.A(G120gat), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n798), .A2(new_n803), .A3(new_n610), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n802), .A2(new_n804), .ZN(G1341gat));
  NAND3_X1  g604(.A1(new_n794), .A2(new_n317), .A3(new_n575), .ZN(new_n806));
  OAI21_X1  g605(.A(G127gat), .B1(new_n798), .B2(new_n576), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(G1342gat));
  NOR2_X1   g607(.A1(new_n536), .A2(G134gat), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT56), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT56), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n794), .A2(new_n812), .A3(new_n809), .ZN(new_n813));
  OAI21_X1  g612(.A(G134gat), .B1(new_n798), .B2(new_n536), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n811), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT117), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n811), .A2(new_n817), .A3(new_n813), .A4(new_n814), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(G1343gat));
  AOI21_X1  g618(.A(KEYINPUT57), .B1(new_n791), .B2(new_n672), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n672), .A2(KEYINPUT57), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n780), .B1(new_n767), .B2(new_n508), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n536), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n786), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n576), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n821), .B1(new_n790), .B2(new_n825), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n626), .B(new_n797), .C1(new_n820), .C2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(G141gat), .B1(new_n827), .B2(new_n508), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n626), .A2(new_n672), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT119), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n626), .A2(KEYINPUT119), .A3(new_n672), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n437), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n508), .A2(G141gat), .ZN(new_n834));
  XOR2_X1   g633(.A(new_n834), .B(KEYINPUT120), .Z(new_n835));
  AND2_X1   g634(.A1(new_n792), .A2(KEYINPUT118), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n792), .A2(KEYINPUT118), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n833), .B(new_n835), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n828), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(KEYINPUT58), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT58), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n828), .A2(new_n841), .A3(new_n838), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(G1344gat));
  OAI21_X1  g642(.A(new_n833), .B1(new_n836), .B2(new_n837), .ZN(new_n844));
  OR3_X1    g643(.A1(new_n844), .A2(G148gat), .A3(new_n610), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n785), .A2(new_n772), .A3(new_n757), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n575), .B1(new_n847), .B2(new_n823), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n672), .B1(new_n848), .B2(new_n789), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n821), .B1(new_n788), .B2(new_n790), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n851), .B1(new_n852), .B2(KEYINPUT121), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n854));
  AOI211_X1 g653(.A(new_n854), .B(new_n821), .C1(new_n788), .C2(new_n790), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NOR4_X1   g655(.A1(new_n423), .A2(new_n382), .A3(new_n437), .A4(new_n610), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n846), .B1(new_n858), .B2(G148gat), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n827), .A2(new_n610), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n846), .A2(G148gat), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n845), .B1(new_n859), .B2(new_n862), .ZN(G1345gat));
  OAI21_X1  g662(.A(G155gat), .B1(new_n827), .B2(new_n576), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n575), .A2(new_n210), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(new_n844), .B2(new_n865), .ZN(G1346gat));
  NOR3_X1   g665(.A1(new_n827), .A2(new_n211), .A3(new_n536), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n844), .A2(new_n536), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n867), .B1(new_n868), .B2(new_n211), .ZN(G1347gat));
  AOI21_X1  g668(.A(new_n438), .B1(new_n788), .B2(new_n790), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n419), .A2(new_n386), .A3(new_n437), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OR3_X1    g671(.A1(new_n872), .A2(G169gat), .A3(new_n508), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n616), .A2(new_n438), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n796), .A2(new_n694), .A3(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n702), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n877), .A2(new_n878), .A3(G169gat), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(new_n877), .B2(G169gat), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n873), .B1(new_n879), .B2(new_n880), .ZN(G1348gat));
  OAI21_X1  g680(.A(G176gat), .B1(new_n875), .B2(new_n610), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n610), .A2(G176gat), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n882), .B1(new_n872), .B2(new_n883), .ZN(G1349gat));
  OAI21_X1  g683(.A(G183gat), .B1(new_n875), .B2(new_n576), .ZN(new_n885));
  INV_X1    g684(.A(new_n872), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n575), .A2(new_n287), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n886), .A2(KEYINPUT123), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT123), .B1(new_n886), .B2(new_n887), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n885), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(KEYINPUT60), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT60), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n892), .B(new_n885), .C1(new_n888), .C2(new_n889), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n893), .ZN(G1350gat));
  NAND3_X1  g693(.A1(new_n886), .A2(new_n288), .A3(new_n537), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT61), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n876), .A2(new_n537), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(G190gat), .ZN(new_n898));
  AOI211_X1 g697(.A(KEYINPUT61), .B(new_n288), .C1(new_n876), .C2(new_n537), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n895), .B1(new_n898), .B2(new_n899), .ZN(G1351gat));
  NOR2_X1   g699(.A1(new_n829), .A2(new_n616), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n870), .A2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  XOR2_X1   g702(.A(KEYINPUT124), .B(G197gat), .Z(new_n904));
  NAND3_X1  g703(.A1(new_n903), .A2(new_n702), .A3(new_n904), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n423), .A2(new_n438), .A3(new_n616), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n856), .A2(new_n702), .A3(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n905), .B1(new_n908), .B2(new_n904), .ZN(G1352gat));
  XNOR2_X1  g708(.A(KEYINPUT125), .B(G204gat), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n902), .A2(new_n610), .A3(new_n910), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT62), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n609), .B(new_n906), .C1(new_n853), .C2(new_n855), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n913), .A2(KEYINPUT126), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n910), .B1(new_n913), .B2(KEYINPUT126), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(G1353gat));
  NAND3_X1  g715(.A1(new_n903), .A2(new_n228), .A3(new_n575), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n575), .B(new_n906), .C1(new_n853), .C2(new_n855), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n918), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n919));
  AOI21_X1  g718(.A(KEYINPUT63), .B1(new_n918), .B2(G211gat), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(G1354gat));
  OAI211_X1 g720(.A(new_n537), .B(new_n906), .C1(new_n853), .C2(new_n855), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(G218gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n903), .A2(new_n229), .A3(new_n537), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT127), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT127), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n923), .A2(new_n927), .A3(new_n924), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(G1355gat));
endmodule


