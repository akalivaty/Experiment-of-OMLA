

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U551 ( .A1(G2104), .A2(n522), .ZN(n883) );
  NOR2_X2 U552 ( .A1(n569), .A2(n568), .ZN(n570) );
  OR2_X1 U553 ( .A1(n751), .A2(KEYINPUT33), .ZN(n757) );
  BUF_X1 U554 ( .A(n685), .Z(n684) );
  NAND2_X2 U555 ( .A1(n683), .A2(n770), .ZN(n718) );
  NOR2_X4 U556 ( .A1(n522), .A2(n525), .ZN(n882) );
  INV_X1 U557 ( .A(KEYINPUT17), .ZN(n517) );
  NAND2_X1 U558 ( .A1(G8), .A2(n732), .ZN(n516) );
  AND2_X1 U559 ( .A1(G2067), .A2(n711), .ZN(n693) );
  OR2_X1 U560 ( .A1(n993), .A2(n698), .ZN(n699) );
  NOR2_X1 U561 ( .A1(n717), .A2(n716), .ZN(n728) );
  INV_X1 U562 ( .A(G286), .ZN(n735) );
  INV_X1 U563 ( .A(KEYINPUT105), .ZN(n730) );
  INV_X1 U564 ( .A(n1010), .ZN(n754) );
  NOR2_X1 U565 ( .A1(n755), .A2(n754), .ZN(n756) );
  INV_X1 U566 ( .A(KEYINPUT70), .ZN(n565) );
  XNOR2_X1 U567 ( .A(n565), .B(KEYINPUT13), .ZN(n566) );
  XNOR2_X1 U568 ( .A(n567), .B(n566), .ZN(n568) );
  INV_X1 U569 ( .A(G2104), .ZN(n525) );
  NOR2_X1 U570 ( .A1(G543), .A2(n534), .ZN(n535) );
  NOR2_X1 U571 ( .A1(n640), .A2(n534), .ZN(n649) );
  NOR2_X1 U572 ( .A1(G651), .A2(G543), .ZN(n648) );
  NOR2_X1 U573 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U574 ( .A(n529), .B(KEYINPUT66), .ZN(n682) );
  BUF_X1 U575 ( .A(n682), .Z(G160) );
  INV_X1 U576 ( .A(G2105), .ZN(n522) );
  NAND2_X1 U577 ( .A1(G113), .A2(n882), .ZN(n520) );
  NOR2_X1 U578 ( .A1(G2105), .A2(G2104), .ZN(n518) );
  XNOR2_X1 U579 ( .A(n518), .B(n517), .ZN(n545) );
  NAND2_X1 U580 ( .A1(n545), .A2(G137), .ZN(n519) );
  NAND2_X1 U581 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U582 ( .A(n521), .B(KEYINPUT67), .ZN(n524) );
  NAND2_X1 U583 ( .A1(G125), .A2(n883), .ZN(n523) );
  NAND2_X1 U584 ( .A1(n524), .A2(n523), .ZN(n528) );
  NOR2_X2 U585 ( .A1(G2105), .A2(n525), .ZN(n887) );
  NAND2_X1 U586 ( .A1(G101), .A2(n887), .ZN(n526) );
  XNOR2_X1 U587 ( .A(KEYINPUT23), .B(n526), .ZN(n527) );
  NAND2_X1 U588 ( .A1(n648), .A2(G89), .ZN(n530) );
  XNOR2_X1 U589 ( .A(n530), .B(KEYINPUT4), .ZN(n532) );
  XOR2_X1 U590 ( .A(KEYINPUT0), .B(G543), .Z(n640) );
  INV_X1 U591 ( .A(G651), .ZN(n534) );
  NAND2_X1 U592 ( .A1(G76), .A2(n649), .ZN(n531) );
  NAND2_X1 U593 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U594 ( .A(KEYINPUT5), .B(n533), .ZN(n541) );
  XOR2_X1 U595 ( .A(KEYINPUT1), .B(n535), .Z(n644) );
  NAND2_X1 U596 ( .A1(G63), .A2(n644), .ZN(n537) );
  NOR2_X2 U597 ( .A1(G651), .A2(n640), .ZN(n645) );
  NAND2_X1 U598 ( .A1(G51), .A2(n645), .ZN(n536) );
  NAND2_X1 U599 ( .A1(n537), .A2(n536), .ZN(n539) );
  XOR2_X1 U600 ( .A(KEYINPUT74), .B(KEYINPUT6), .Z(n538) );
  XNOR2_X1 U601 ( .A(n539), .B(n538), .ZN(n540) );
  NAND2_X1 U602 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U603 ( .A(KEYINPUT7), .B(n542), .ZN(G168) );
  XOR2_X1 U604 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U605 ( .A1(G114), .A2(n882), .ZN(n544) );
  NAND2_X1 U606 ( .A1(G126), .A2(n883), .ZN(n543) );
  NAND2_X1 U607 ( .A1(n544), .A2(n543), .ZN(n550) );
  NAND2_X1 U608 ( .A1(G102), .A2(n887), .ZN(n547) );
  NAND2_X1 U609 ( .A1(G138), .A2(n545), .ZN(n546) );
  NAND2_X1 U610 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U611 ( .A(KEYINPUT93), .B(n548), .Z(n549) );
  NOR2_X1 U612 ( .A1(n550), .A2(n549), .ZN(G164) );
  NAND2_X1 U613 ( .A1(G60), .A2(n644), .ZN(n552) );
  NAND2_X1 U614 ( .A1(G47), .A2(n645), .ZN(n551) );
  NAND2_X1 U615 ( .A1(n552), .A2(n551), .ZN(n556) );
  NAND2_X1 U616 ( .A1(G85), .A2(n648), .ZN(n554) );
  NAND2_X1 U617 ( .A1(G72), .A2(n649), .ZN(n553) );
  NAND2_X1 U618 ( .A1(n554), .A2(n553), .ZN(n555) );
  OR2_X1 U619 ( .A1(n556), .A2(n555), .ZN(G290) );
  AND2_X1 U620 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U621 ( .A(G132), .ZN(G219) );
  INV_X1 U622 ( .A(G69), .ZN(G235) );
  NAND2_X1 U623 ( .A1(G7), .A2(G661), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U625 ( .A(G223), .ZN(n833) );
  NAND2_X1 U626 ( .A1(n833), .A2(G567), .ZN(n558) );
  XOR2_X1 U627 ( .A(KEYINPUT11), .B(n558), .Z(G234) );
  NAND2_X1 U628 ( .A1(n644), .A2(G56), .ZN(n559) );
  XNOR2_X1 U629 ( .A(n559), .B(KEYINPUT14), .ZN(n561) );
  NAND2_X1 U630 ( .A1(G43), .A2(n645), .ZN(n560) );
  NAND2_X1 U631 ( .A1(n561), .A2(n560), .ZN(n569) );
  NAND2_X1 U632 ( .A1(n648), .A2(G81), .ZN(n562) );
  XNOR2_X1 U633 ( .A(n562), .B(KEYINPUT12), .ZN(n564) );
  NAND2_X1 U634 ( .A1(G68), .A2(n649), .ZN(n563) );
  NAND2_X1 U635 ( .A1(n564), .A2(n563), .ZN(n567) );
  XNOR2_X2 U636 ( .A(KEYINPUT71), .B(n570), .ZN(n1005) );
  INV_X1 U637 ( .A(n1005), .ZN(n571) );
  NAND2_X1 U638 ( .A1(n571), .A2(G860), .ZN(G153) );
  NAND2_X1 U639 ( .A1(G90), .A2(n648), .ZN(n573) );
  NAND2_X1 U640 ( .A1(G77), .A2(n649), .ZN(n572) );
  NAND2_X1 U641 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U642 ( .A(KEYINPUT9), .B(n574), .ZN(n578) );
  NAND2_X1 U643 ( .A1(G64), .A2(n644), .ZN(n576) );
  NAND2_X1 U644 ( .A1(G52), .A2(n645), .ZN(n575) );
  AND2_X1 U645 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U646 ( .A1(n578), .A2(n577), .ZN(G301) );
  NAND2_X1 U647 ( .A1(G79), .A2(n649), .ZN(n585) );
  NAND2_X1 U648 ( .A1(G66), .A2(n644), .ZN(n580) );
  NAND2_X1 U649 ( .A1(G92), .A2(n648), .ZN(n579) );
  NAND2_X1 U650 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U651 ( .A1(n645), .A2(G54), .ZN(n581) );
  XOR2_X1 U652 ( .A(KEYINPUT72), .B(n581), .Z(n582) );
  NOR2_X1 U653 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U655 ( .A(n586), .B(KEYINPUT15), .ZN(n993) );
  NOR2_X1 U656 ( .A1(n993), .A2(G868), .ZN(n587) );
  XNOR2_X1 U657 ( .A(n587), .B(KEYINPUT73), .ZN(n589) );
  NAND2_X1 U658 ( .A1(G868), .A2(G301), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n589), .A2(n588), .ZN(G284) );
  NAND2_X1 U660 ( .A1(G65), .A2(n644), .ZN(n591) );
  NAND2_X1 U661 ( .A1(G53), .A2(n645), .ZN(n590) );
  NAND2_X1 U662 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U663 ( .A1(G91), .A2(n648), .ZN(n593) );
  NAND2_X1 U664 ( .A1(G78), .A2(n649), .ZN(n592) );
  NAND2_X1 U665 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U666 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U667 ( .A(KEYINPUT68), .B(n596), .Z(G299) );
  XNOR2_X1 U668 ( .A(KEYINPUT75), .B(G868), .ZN(n597) );
  NOR2_X1 U669 ( .A1(G286), .A2(n597), .ZN(n599) );
  NOR2_X1 U670 ( .A1(G299), .A2(G868), .ZN(n598) );
  NOR2_X1 U671 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U672 ( .A(KEYINPUT76), .B(n600), .ZN(G297) );
  INV_X1 U673 ( .A(G559), .ZN(n604) );
  NOR2_X1 U674 ( .A1(G860), .A2(n604), .ZN(n601) );
  XNOR2_X1 U675 ( .A(KEYINPUT77), .B(n601), .ZN(n602) );
  NAND2_X1 U676 ( .A1(n602), .A2(n993), .ZN(n603) );
  XNOR2_X1 U677 ( .A(n603), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U678 ( .A1(n604), .A2(n993), .ZN(n605) );
  NAND2_X1 U679 ( .A1(n605), .A2(G868), .ZN(n607) );
  INV_X1 U680 ( .A(G868), .ZN(n662) );
  NAND2_X1 U681 ( .A1(n1005), .A2(n662), .ZN(n606) );
  NAND2_X1 U682 ( .A1(n607), .A2(n606), .ZN(G282) );
  XNOR2_X1 U683 ( .A(G2100), .B(KEYINPUT83), .ZN(n621) );
  XOR2_X1 U684 ( .A(KEYINPUT18), .B(KEYINPUT78), .Z(n609) );
  NAND2_X1 U685 ( .A1(G123), .A2(n883), .ZN(n608) );
  XNOR2_X1 U686 ( .A(n609), .B(n608), .ZN(n612) );
  BUF_X1 U687 ( .A(n545), .Z(n890) );
  NAND2_X1 U688 ( .A1(n890), .A2(G135), .ZN(n610) );
  XNOR2_X1 U689 ( .A(KEYINPUT79), .B(n610), .ZN(n611) );
  NOR2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U691 ( .A(KEYINPUT80), .B(n613), .ZN(n618) );
  NAND2_X1 U692 ( .A1(G99), .A2(n887), .ZN(n615) );
  NAND2_X1 U693 ( .A1(G111), .A2(n882), .ZN(n614) );
  NAND2_X1 U694 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U695 ( .A(KEYINPUT81), .B(n616), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n618), .A2(n617), .ZN(n962) );
  XOR2_X1 U697 ( .A(G2096), .B(KEYINPUT82), .Z(n619) );
  XNOR2_X1 U698 ( .A(n962), .B(n619), .ZN(n620) );
  NAND2_X1 U699 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U700 ( .A(n622), .B(KEYINPUT84), .ZN(G156) );
  NAND2_X1 U701 ( .A1(G88), .A2(n648), .ZN(n623) );
  XNOR2_X1 U702 ( .A(n623), .B(KEYINPUT86), .ZN(n625) );
  NAND2_X1 U703 ( .A1(n644), .A2(G62), .ZN(n624) );
  NAND2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U705 ( .A1(G50), .A2(n645), .ZN(n627) );
  NAND2_X1 U706 ( .A1(G75), .A2(n649), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U708 ( .A1(n629), .A2(n628), .ZN(G166) );
  NAND2_X1 U709 ( .A1(G61), .A2(n644), .ZN(n631) );
  NAND2_X1 U710 ( .A1(G48), .A2(n645), .ZN(n630) );
  NAND2_X1 U711 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U712 ( .A1(n649), .A2(G73), .ZN(n632) );
  XOR2_X1 U713 ( .A(KEYINPUT2), .B(n632), .Z(n633) );
  NOR2_X1 U714 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U715 ( .A1(n648), .A2(G86), .ZN(n635) );
  NAND2_X1 U716 ( .A1(n636), .A2(n635), .ZN(G305) );
  NAND2_X1 U717 ( .A1(G49), .A2(n645), .ZN(n638) );
  NAND2_X1 U718 ( .A1(G74), .A2(G651), .ZN(n637) );
  NAND2_X1 U719 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U720 ( .A1(n644), .A2(n639), .ZN(n642) );
  NAND2_X1 U721 ( .A1(n640), .A2(G87), .ZN(n641) );
  NAND2_X1 U722 ( .A1(n642), .A2(n641), .ZN(G288) );
  NAND2_X1 U723 ( .A1(G559), .A2(n993), .ZN(n643) );
  XNOR2_X1 U724 ( .A(n643), .B(n1005), .ZN(n839) );
  NAND2_X1 U725 ( .A1(G67), .A2(n644), .ZN(n647) );
  NAND2_X1 U726 ( .A1(G55), .A2(n645), .ZN(n646) );
  NAND2_X1 U727 ( .A1(n647), .A2(n646), .ZN(n653) );
  NAND2_X1 U728 ( .A1(G93), .A2(n648), .ZN(n651) );
  NAND2_X1 U729 ( .A1(G80), .A2(n649), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U731 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U732 ( .A(KEYINPUT85), .B(n654), .ZN(n840) );
  XNOR2_X1 U733 ( .A(G166), .B(KEYINPUT19), .ZN(n655) );
  XNOR2_X1 U734 ( .A(n655), .B(KEYINPUT87), .ZN(n656) );
  XOR2_X1 U735 ( .A(n840), .B(n656), .Z(n658) );
  XNOR2_X1 U736 ( .A(G305), .B(G299), .ZN(n657) );
  XNOR2_X1 U737 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U738 ( .A(n659), .B(G290), .ZN(n660) );
  XNOR2_X1 U739 ( .A(n660), .B(G288), .ZN(n903) );
  XNOR2_X1 U740 ( .A(n839), .B(n903), .ZN(n661) );
  NAND2_X1 U741 ( .A1(n661), .A2(G868), .ZN(n664) );
  NAND2_X1 U742 ( .A1(n662), .A2(n840), .ZN(n663) );
  NAND2_X1 U743 ( .A1(n664), .A2(n663), .ZN(G295) );
  NAND2_X1 U744 ( .A1(G2084), .A2(G2078), .ZN(n665) );
  XOR2_X1 U745 ( .A(KEYINPUT20), .B(n665), .Z(n666) );
  NAND2_X1 U746 ( .A1(n666), .A2(G2090), .ZN(n667) );
  XNOR2_X1 U747 ( .A(n667), .B(KEYINPUT21), .ZN(n668) );
  XNOR2_X1 U748 ( .A(KEYINPUT88), .B(n668), .ZN(n669) );
  NAND2_X1 U749 ( .A1(n669), .A2(G2072), .ZN(n670) );
  XOR2_X1 U750 ( .A(KEYINPUT89), .B(n670), .Z(G158) );
  XNOR2_X1 U751 ( .A(KEYINPUT90), .B(G44), .ZN(n671) );
  XNOR2_X1 U752 ( .A(n671), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U753 ( .A(KEYINPUT69), .B(G82), .ZN(G220) );
  NAND2_X1 U754 ( .A1(G120), .A2(G57), .ZN(n672) );
  NOR2_X1 U755 ( .A1(G235), .A2(n672), .ZN(n673) );
  XNOR2_X1 U756 ( .A(KEYINPUT92), .B(n673), .ZN(n674) );
  NAND2_X1 U757 ( .A1(n674), .A2(G108), .ZN(n837) );
  NAND2_X1 U758 ( .A1(n837), .A2(G567), .ZN(n680) );
  NOR2_X1 U759 ( .A1(G219), .A2(G220), .ZN(n676) );
  XNOR2_X1 U760 ( .A(KEYINPUT22), .B(KEYINPUT91), .ZN(n675) );
  XNOR2_X1 U761 ( .A(n676), .B(n675), .ZN(n677) );
  NOR2_X1 U762 ( .A1(G218), .A2(n677), .ZN(n678) );
  NAND2_X1 U763 ( .A1(G96), .A2(n678), .ZN(n838) );
  NAND2_X1 U764 ( .A1(n838), .A2(G2106), .ZN(n679) );
  NAND2_X1 U765 ( .A1(n680), .A2(n679), .ZN(n842) );
  NAND2_X1 U766 ( .A1(G661), .A2(G483), .ZN(n681) );
  NOR2_X1 U767 ( .A1(n842), .A2(n681), .ZN(n836) );
  NAND2_X1 U768 ( .A1(n836), .A2(G36), .ZN(G176) );
  INV_X1 U769 ( .A(G166), .ZN(G303) );
  INV_X1 U770 ( .A(G301), .ZN(G171) );
  NAND2_X1 U771 ( .A1(n682), .A2(G40), .ZN(n771) );
  INV_X1 U772 ( .A(n771), .ZN(n683) );
  NOR2_X1 U773 ( .A1(G164), .A2(G1384), .ZN(n770) );
  NAND2_X1 U774 ( .A1(G8), .A2(n718), .ZN(n685) );
  NOR2_X1 U775 ( .A1(G1966), .A2(n685), .ZN(n729) );
  AND2_X1 U776 ( .A1(n718), .A2(G1341), .ZN(n686) );
  NOR2_X1 U777 ( .A1(n686), .A2(n1005), .ZN(n690) );
  INV_X2 U778 ( .A(n718), .ZN(n711) );
  NAND2_X1 U779 ( .A1(n711), .A2(G1996), .ZN(n688) );
  XNOR2_X1 U780 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n687) );
  XNOR2_X1 U781 ( .A(n688), .B(n687), .ZN(n689) );
  AND2_X1 U782 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U783 ( .A(n691), .B(KEYINPUT65), .ZN(n697) );
  INV_X1 U784 ( .A(KEYINPUT103), .ZN(n692) );
  XNOR2_X1 U785 ( .A(n693), .B(n692), .ZN(n695) );
  INV_X1 U786 ( .A(G1348), .ZN(n994) );
  NOR2_X1 U787 ( .A1(n994), .A2(n711), .ZN(n694) );
  NOR2_X1 U788 ( .A1(n695), .A2(n694), .ZN(n698) );
  NAND2_X1 U789 ( .A1(n993), .A2(n698), .ZN(n696) );
  NAND2_X1 U790 ( .A1(n697), .A2(n696), .ZN(n700) );
  NAND2_X1 U791 ( .A1(n700), .A2(n699), .ZN(n705) );
  NAND2_X1 U792 ( .A1(n711), .A2(G2072), .ZN(n701) );
  XNOR2_X1 U793 ( .A(n701), .B(KEYINPUT27), .ZN(n703) );
  AND2_X1 U794 ( .A1(G1956), .A2(n718), .ZN(n702) );
  NOR2_X1 U795 ( .A1(n703), .A2(n702), .ZN(n706) );
  INV_X1 U796 ( .A(G299), .ZN(n1001) );
  NAND2_X1 U797 ( .A1(n706), .A2(n1001), .ZN(n704) );
  NAND2_X1 U798 ( .A1(n705), .A2(n704), .ZN(n709) );
  NOR2_X1 U799 ( .A1(n706), .A2(n1001), .ZN(n707) );
  XOR2_X1 U800 ( .A(n707), .B(KEYINPUT28), .Z(n708) );
  NAND2_X1 U801 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U802 ( .A(n710), .B(KEYINPUT29), .ZN(n717) );
  XOR2_X1 U803 ( .A(G2078), .B(KEYINPUT25), .Z(n944) );
  NOR2_X1 U804 ( .A1(n944), .A2(n718), .ZN(n713) );
  NOR2_X1 U805 ( .A1(n711), .A2(G1961), .ZN(n712) );
  NOR2_X1 U806 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U807 ( .A(KEYINPUT101), .B(n714), .ZN(n722) );
  AND2_X1 U808 ( .A1(n722), .A2(G171), .ZN(n715) );
  XNOR2_X1 U809 ( .A(n715), .B(KEYINPUT102), .ZN(n716) );
  NOR2_X1 U810 ( .A1(G2084), .A2(n718), .ZN(n732) );
  NOR2_X1 U811 ( .A1(n729), .A2(n732), .ZN(n719) );
  NAND2_X1 U812 ( .A1(G8), .A2(n719), .ZN(n720) );
  XNOR2_X1 U813 ( .A(KEYINPUT30), .B(n720), .ZN(n721) );
  NOR2_X1 U814 ( .A1(n721), .A2(G168), .ZN(n724) );
  NOR2_X1 U815 ( .A1(G171), .A2(n722), .ZN(n723) );
  NOR2_X1 U816 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U817 ( .A(n725), .B(KEYINPUT31), .ZN(n726) );
  XNOR2_X1 U818 ( .A(KEYINPUT104), .B(n726), .ZN(n727) );
  NOR2_X1 U819 ( .A1(n728), .A2(n727), .ZN(n736) );
  NOR2_X1 U820 ( .A1(n729), .A2(n736), .ZN(n731) );
  XNOR2_X1 U821 ( .A(n731), .B(n730), .ZN(n733) );
  NAND2_X1 U822 ( .A1(n733), .A2(n516), .ZN(n734) );
  XNOR2_X1 U823 ( .A(n734), .B(KEYINPUT106), .ZN(n746) );
  OR2_X1 U824 ( .A1(n736), .A2(n735), .ZN(n742) );
  NOR2_X1 U825 ( .A1(G1971), .A2(n684), .ZN(n738) );
  NOR2_X1 U826 ( .A1(G2090), .A2(n718), .ZN(n737) );
  NOR2_X1 U827 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U828 ( .A(KEYINPUT107), .B(n739), .Z(n740) );
  NAND2_X1 U829 ( .A1(n740), .A2(G303), .ZN(n741) );
  NAND2_X1 U830 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U831 ( .A1(G8), .A2(n743), .ZN(n744) );
  XNOR2_X1 U832 ( .A(n744), .B(KEYINPUT32), .ZN(n745) );
  NAND2_X1 U833 ( .A1(n746), .A2(n745), .ZN(n758) );
  NOR2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n752) );
  NOR2_X1 U835 ( .A1(G1971), .A2(G303), .ZN(n747) );
  NOR2_X1 U836 ( .A1(n752), .A2(n747), .ZN(n998) );
  NAND2_X1 U837 ( .A1(n758), .A2(n998), .ZN(n748) );
  NAND2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n992) );
  NAND2_X1 U839 ( .A1(n748), .A2(n992), .ZN(n749) );
  XNOR2_X1 U840 ( .A(n749), .B(KEYINPUT108), .ZN(n750) );
  NOR2_X1 U841 ( .A1(n684), .A2(n750), .ZN(n751) );
  NAND2_X1 U842 ( .A1(n752), .A2(KEYINPUT33), .ZN(n753) );
  NOR2_X1 U843 ( .A1(n753), .A2(n684), .ZN(n755) );
  XOR2_X1 U844 ( .A(G1981), .B(G305), .Z(n1010) );
  NAND2_X1 U845 ( .A1(n757), .A2(n756), .ZN(n768) );
  NOR2_X1 U846 ( .A1(G2090), .A2(G303), .ZN(n759) );
  NAND2_X1 U847 ( .A1(G8), .A2(n759), .ZN(n760) );
  NAND2_X1 U848 ( .A1(n758), .A2(n760), .ZN(n761) );
  NAND2_X1 U849 ( .A1(n684), .A2(n761), .ZN(n762) );
  XNOR2_X1 U850 ( .A(n762), .B(KEYINPUT109), .ZN(n766) );
  NOR2_X1 U851 ( .A1(G1981), .A2(G305), .ZN(n763) );
  XOR2_X1 U852 ( .A(n763), .B(KEYINPUT24), .Z(n764) );
  NOR2_X1 U853 ( .A1(n684), .A2(n764), .ZN(n765) );
  NOR2_X1 U854 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U856 ( .A(n769), .B(KEYINPUT110), .ZN(n807) );
  XNOR2_X1 U857 ( .A(G1986), .B(G290), .ZN(n1000) );
  NOR2_X1 U858 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U859 ( .A(n772), .B(KEYINPUT94), .ZN(n818) );
  NAND2_X1 U860 ( .A1(n1000), .A2(n818), .ZN(n805) );
  NAND2_X1 U861 ( .A1(G107), .A2(n882), .ZN(n774) );
  NAND2_X1 U862 ( .A1(G119), .A2(n883), .ZN(n773) );
  NAND2_X1 U863 ( .A1(n774), .A2(n773), .ZN(n779) );
  NAND2_X1 U864 ( .A1(G95), .A2(n887), .ZN(n776) );
  NAND2_X1 U865 ( .A1(G131), .A2(n890), .ZN(n775) );
  NAND2_X1 U866 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U867 ( .A(KEYINPUT95), .B(n777), .Z(n778) );
  NOR2_X1 U868 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U869 ( .A(KEYINPUT96), .B(n780), .Z(n878) );
  NAND2_X1 U870 ( .A1(G1991), .A2(n878), .ZN(n781) );
  XOR2_X1 U871 ( .A(KEYINPUT97), .B(n781), .Z(n792) );
  NAND2_X1 U872 ( .A1(G117), .A2(n882), .ZN(n782) );
  XOR2_X1 U873 ( .A(KEYINPUT98), .B(n782), .Z(n785) );
  NAND2_X1 U874 ( .A1(n887), .A2(G105), .ZN(n783) );
  XOR2_X1 U875 ( .A(KEYINPUT38), .B(n783), .Z(n784) );
  NOR2_X1 U876 ( .A1(n785), .A2(n784), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n883), .A2(G129), .ZN(n786) );
  NAND2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U879 ( .A(n788), .B(KEYINPUT99), .ZN(n790) );
  NAND2_X1 U880 ( .A1(G141), .A2(n890), .ZN(n789) );
  NAND2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n894) );
  NAND2_X1 U882 ( .A1(G1996), .A2(n894), .ZN(n791) );
  NAND2_X1 U883 ( .A1(n792), .A2(n791), .ZN(n984) );
  NAND2_X1 U884 ( .A1(n818), .A2(n984), .ZN(n793) );
  XOR2_X1 U885 ( .A(KEYINPUT100), .B(n793), .Z(n810) );
  NAND2_X1 U886 ( .A1(G104), .A2(n887), .ZN(n795) );
  NAND2_X1 U887 ( .A1(G140), .A2(n890), .ZN(n794) );
  NAND2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U889 ( .A(KEYINPUT34), .B(n796), .ZN(n801) );
  NAND2_X1 U890 ( .A1(G116), .A2(n882), .ZN(n798) );
  NAND2_X1 U891 ( .A1(G128), .A2(n883), .ZN(n797) );
  NAND2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U893 ( .A(KEYINPUT35), .B(n799), .Z(n800) );
  NOR2_X1 U894 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U895 ( .A(KEYINPUT36), .B(n802), .ZN(n877) );
  XNOR2_X1 U896 ( .A(G2067), .B(KEYINPUT37), .ZN(n815) );
  NOR2_X1 U897 ( .A1(n877), .A2(n815), .ZN(n971) );
  NAND2_X1 U898 ( .A1(n971), .A2(n818), .ZN(n813) );
  INV_X1 U899 ( .A(n813), .ZN(n803) );
  NOR2_X1 U900 ( .A1(n810), .A2(n803), .ZN(n804) );
  AND2_X1 U901 ( .A1(n805), .A2(n804), .ZN(n806) );
  NAND2_X1 U902 ( .A1(n807), .A2(n806), .ZN(n821) );
  NOR2_X1 U903 ( .A1(G1996), .A2(n894), .ZN(n967) );
  NOR2_X1 U904 ( .A1(G1991), .A2(n878), .ZN(n965) );
  NOR2_X1 U905 ( .A1(G1986), .A2(G290), .ZN(n808) );
  NOR2_X1 U906 ( .A1(n965), .A2(n808), .ZN(n809) );
  NOR2_X1 U907 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U908 ( .A1(n967), .A2(n811), .ZN(n812) );
  XNOR2_X1 U909 ( .A(n812), .B(KEYINPUT39), .ZN(n814) );
  NAND2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n816) );
  NAND2_X1 U911 ( .A1(n877), .A2(n815), .ZN(n972) );
  NAND2_X1 U912 ( .A1(n816), .A2(n972), .ZN(n817) );
  XOR2_X1 U913 ( .A(KEYINPUT111), .B(n817), .Z(n819) );
  NAND2_X1 U914 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U915 ( .A1(n821), .A2(n820), .ZN(n823) );
  XNOR2_X1 U916 ( .A(KEYINPUT112), .B(KEYINPUT40), .ZN(n822) );
  XNOR2_X1 U917 ( .A(n823), .B(n822), .ZN(G329) );
  XNOR2_X1 U918 ( .A(G1341), .B(G2454), .ZN(n824) );
  XNOR2_X1 U919 ( .A(n824), .B(G2430), .ZN(n825) );
  XNOR2_X1 U920 ( .A(n825), .B(G1348), .ZN(n831) );
  XOR2_X1 U921 ( .A(G2443), .B(G2427), .Z(n827) );
  XNOR2_X1 U922 ( .A(G2438), .B(G2446), .ZN(n826) );
  XNOR2_X1 U923 ( .A(n827), .B(n826), .ZN(n829) );
  XOR2_X1 U924 ( .A(G2451), .B(G2435), .Z(n828) );
  XNOR2_X1 U925 ( .A(n829), .B(n828), .ZN(n830) );
  XNOR2_X1 U926 ( .A(n831), .B(n830), .ZN(n832) );
  NAND2_X1 U927 ( .A1(n832), .A2(G14), .ZN(n908) );
  XNOR2_X1 U928 ( .A(KEYINPUT113), .B(n908), .ZN(G401) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U931 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U933 ( .A1(n836), .A2(n835), .ZN(G188) );
  XOR2_X1 U934 ( .A(G120), .B(KEYINPUT114), .Z(G236) );
  INV_X1 U936 ( .A(G108), .ZN(G238) );
  INV_X1 U937 ( .A(G96), .ZN(G221) );
  INV_X1 U938 ( .A(G57), .ZN(G237) );
  NOR2_X1 U939 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U940 ( .A(G325), .ZN(G261) );
  NOR2_X1 U941 ( .A1(n839), .A2(G860), .ZN(n841) );
  XOR2_X1 U942 ( .A(n841), .B(n840), .Z(G145) );
  INV_X1 U943 ( .A(n842), .ZN(G319) );
  XOR2_X1 U944 ( .A(KEYINPUT115), .B(G2072), .Z(n844) );
  XNOR2_X1 U945 ( .A(G2084), .B(G2078), .ZN(n843) );
  XNOR2_X1 U946 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U947 ( .A(n845), .B(G2096), .Z(n847) );
  XNOR2_X1 U948 ( .A(G2067), .B(G2090), .ZN(n846) );
  XNOR2_X1 U949 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U950 ( .A(G2100), .B(G2678), .Z(n849) );
  XNOR2_X1 U951 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n848) );
  XNOR2_X1 U952 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U953 ( .A(n851), .B(n850), .Z(G227) );
  XOR2_X1 U954 ( .A(G1961), .B(G1966), .Z(n853) );
  XNOR2_X1 U955 ( .A(G1981), .B(G1976), .ZN(n852) );
  XNOR2_X1 U956 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U957 ( .A(n854), .B(G2474), .Z(n856) );
  XNOR2_X1 U958 ( .A(G1996), .B(G1991), .ZN(n855) );
  XNOR2_X1 U959 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U960 ( .A(KEYINPUT41), .B(G1956), .Z(n858) );
  XNOR2_X1 U961 ( .A(G1986), .B(G1971), .ZN(n857) );
  XNOR2_X1 U962 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U963 ( .A(n860), .B(n859), .ZN(G229) );
  NAND2_X1 U964 ( .A1(G124), .A2(n883), .ZN(n861) );
  XNOR2_X1 U965 ( .A(n861), .B(KEYINPUT44), .ZN(n862) );
  XNOR2_X1 U966 ( .A(n862), .B(KEYINPUT116), .ZN(n864) );
  NAND2_X1 U967 ( .A1(G100), .A2(n887), .ZN(n863) );
  NAND2_X1 U968 ( .A1(n864), .A2(n863), .ZN(n868) );
  NAND2_X1 U969 ( .A1(G136), .A2(n890), .ZN(n866) );
  NAND2_X1 U970 ( .A1(G112), .A2(n882), .ZN(n865) );
  NAND2_X1 U971 ( .A1(n866), .A2(n865), .ZN(n867) );
  NOR2_X1 U972 ( .A1(n868), .A2(n867), .ZN(G162) );
  NAND2_X1 U973 ( .A1(G118), .A2(n882), .ZN(n870) );
  NAND2_X1 U974 ( .A1(G130), .A2(n883), .ZN(n869) );
  NAND2_X1 U975 ( .A1(n870), .A2(n869), .ZN(n876) );
  NAND2_X1 U976 ( .A1(G106), .A2(n887), .ZN(n872) );
  NAND2_X1 U977 ( .A1(G142), .A2(n890), .ZN(n871) );
  NAND2_X1 U978 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U979 ( .A(KEYINPUT45), .B(n873), .ZN(n874) );
  XNOR2_X1 U980 ( .A(KEYINPUT117), .B(n874), .ZN(n875) );
  NOR2_X1 U981 ( .A1(n876), .A2(n875), .ZN(n881) );
  XNOR2_X1 U982 ( .A(n878), .B(n877), .ZN(n879) );
  XNOR2_X1 U983 ( .A(n879), .B(n962), .ZN(n880) );
  XNOR2_X1 U984 ( .A(n881), .B(n880), .ZN(n896) );
  NAND2_X1 U985 ( .A1(G115), .A2(n882), .ZN(n885) );
  NAND2_X1 U986 ( .A1(G127), .A2(n883), .ZN(n884) );
  NAND2_X1 U987 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U988 ( .A(n886), .B(KEYINPUT47), .ZN(n889) );
  NAND2_X1 U989 ( .A1(G103), .A2(n887), .ZN(n888) );
  NAND2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n893) );
  NAND2_X1 U991 ( .A1(n890), .A2(G139), .ZN(n891) );
  XOR2_X1 U992 ( .A(KEYINPUT118), .B(n891), .Z(n892) );
  NOR2_X1 U993 ( .A1(n893), .A2(n892), .ZN(n974) );
  XNOR2_X1 U994 ( .A(n894), .B(n974), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n901) );
  XNOR2_X1 U996 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n898) );
  XNOR2_X1 U997 ( .A(G160), .B(G162), .ZN(n897) );
  XNOR2_X1 U998 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U999 ( .A(G164), .B(n899), .Z(n900) );
  XNOR2_X1 U1000 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n902), .ZN(G395) );
  XNOR2_X1 U1002 ( .A(n1005), .B(n903), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(G171), .B(n993), .ZN(n904) );
  XNOR2_X1 U1004 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1005 ( .A(G286), .B(n906), .Z(n907) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n907), .ZN(G397) );
  NAND2_X1 U1007 ( .A1(G319), .A2(n908), .ZN(n911) );
  NOR2_X1 U1008 ( .A1(G227), .A2(G229), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(n909), .B(KEYINPUT49), .ZN(n910) );
  NOR2_X1 U1010 ( .A1(n911), .A2(n910), .ZN(n912) );
  XOR2_X1 U1011 ( .A(KEYINPUT119), .B(n912), .Z(n914) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1015 ( .A(G4), .B(KEYINPUT127), .Z(n916) );
  XNOR2_X1 U1016 ( .A(G1348), .B(KEYINPUT59), .ZN(n915) );
  XNOR2_X1 U1017 ( .A(n916), .B(n915), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(G1981), .B(G6), .ZN(n918) );
  XNOR2_X1 U1019 ( .A(G1956), .B(G20), .ZN(n917) );
  NOR2_X1 U1020 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n923) );
  XNOR2_X1 U1022 ( .A(KEYINPUT126), .B(G1341), .ZN(n921) );
  XNOR2_X1 U1023 ( .A(G19), .B(n921), .ZN(n922) );
  NOR2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1025 ( .A(KEYINPUT60), .B(n924), .ZN(n928) );
  XNOR2_X1 U1026 ( .A(G1966), .B(G21), .ZN(n926) );
  XNOR2_X1 U1027 ( .A(G1961), .B(G5), .ZN(n925) );
  NOR2_X1 U1028 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n935) );
  XNOR2_X1 U1030 ( .A(G1976), .B(G23), .ZN(n930) );
  XNOR2_X1 U1031 ( .A(G1971), .B(G22), .ZN(n929) );
  NOR2_X1 U1032 ( .A1(n930), .A2(n929), .ZN(n932) );
  XOR2_X1 U1033 ( .A(G1986), .B(G24), .Z(n931) );
  NAND2_X1 U1034 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1035 ( .A(KEYINPUT58), .B(n933), .ZN(n934) );
  NOR2_X1 U1036 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1037 ( .A(KEYINPUT61), .B(n936), .Z(n937) );
  NOR2_X1 U1038 ( .A1(G16), .A2(n937), .ZN(n961) );
  INV_X1 U1039 ( .A(KEYINPUT55), .ZN(n986) );
  XNOR2_X1 U1040 ( .A(KEYINPUT54), .B(KEYINPUT123), .ZN(n938) );
  XNOR2_X1 U1041 ( .A(n938), .B(G34), .ZN(n939) );
  XNOR2_X1 U1042 ( .A(G2084), .B(n939), .ZN(n955) );
  XNOR2_X1 U1043 ( .A(G2090), .B(G35), .ZN(n953) );
  XOR2_X1 U1044 ( .A(G1991), .B(G25), .Z(n940) );
  NAND2_X1 U1045 ( .A1(n940), .A2(G28), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(G2067), .B(G26), .ZN(n942) );
  XNOR2_X1 U1047 ( .A(G2072), .B(G33), .ZN(n941) );
  NOR2_X1 U1048 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1049 ( .A(KEYINPUT122), .B(n943), .ZN(n948) );
  XNOR2_X1 U1050 ( .A(G1996), .B(G32), .ZN(n946) );
  XNOR2_X1 U1051 ( .A(n944), .B(G27), .ZN(n945) );
  NOR2_X1 U1052 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1053 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1054 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1055 ( .A(KEYINPUT53), .B(n951), .ZN(n952) );
  NOR2_X1 U1056 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1057 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1058 ( .A(n986), .B(n956), .ZN(n958) );
  INV_X1 U1059 ( .A(G29), .ZN(n957) );
  NAND2_X1 U1060 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1061 ( .A1(G11), .A2(n959), .ZN(n960) );
  NOR2_X1 U1062 ( .A1(n961), .A2(n960), .ZN(n990) );
  XNOR2_X1 U1063 ( .A(G160), .B(G2084), .ZN(n963) );
  NAND2_X1 U1064 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1065 ( .A1(n965), .A2(n964), .ZN(n982) );
  XOR2_X1 U1066 ( .A(G2090), .B(G162), .Z(n966) );
  NOR2_X1 U1067 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1068 ( .A(KEYINPUT51), .B(n968), .Z(n969) );
  XOR2_X1 U1069 ( .A(KEYINPUT120), .B(n969), .Z(n970) );
  NOR2_X1 U1070 ( .A1(n971), .A2(n970), .ZN(n973) );
  NAND2_X1 U1071 ( .A1(n973), .A2(n972), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(G2072), .B(n974), .ZN(n976) );
  XNOR2_X1 U1073 ( .A(G164), .B(G2078), .ZN(n975) );
  NAND2_X1 U1074 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1075 ( .A(KEYINPUT50), .B(n977), .Z(n978) );
  XNOR2_X1 U1076 ( .A(KEYINPUT121), .B(n978), .ZN(n979) );
  NOR2_X1 U1077 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1080 ( .A(KEYINPUT52), .B(n985), .ZN(n987) );
  NAND2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1082 ( .A1(n988), .A2(G29), .ZN(n989) );
  NAND2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n1019) );
  NAND2_X1 U1084 ( .A1(G1971), .A2(G303), .ZN(n991) );
  NAND2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(n994), .B(n993), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1009) );
  XNOR2_X1 U1090 ( .A(n1001), .B(G1956), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(G1961), .B(KEYINPUT125), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(n1002), .B(G301), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(G1341), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1015) );
  XNOR2_X1 U1097 ( .A(G168), .B(G1966), .ZN(n1011) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(n1012), .B(KEYINPUT57), .ZN(n1013) );
  XOR2_X1 U1100 ( .A(KEYINPUT124), .B(n1013), .Z(n1014) );
  NOR2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1017) );
  XOR2_X1 U1102 ( .A(G16), .B(KEYINPUT56), .Z(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(n1020), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
endmodule

