

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745;

  OR2_X1 U373 ( .A1(n510), .A2(n509), .ZN(n360) );
  NOR2_X1 U374 ( .A1(n660), .A2(n661), .ZN(n528) );
  NOR2_X1 U375 ( .A1(G902), .A2(n710), .ZN(n439) );
  NOR2_X1 U376 ( .A1(n362), .A2(G237), .ZN(n464) );
  XOR2_X1 U377 ( .A(G146), .B(G125), .Z(n430) );
  XNOR2_X1 U378 ( .A(n360), .B(KEYINPUT76), .ZN(n511) );
  BUF_X1 U379 ( .A(G953), .Z(n362) );
  XNOR2_X2 U380 ( .A(n379), .B(n393), .ZN(n378) );
  XNOR2_X2 U381 ( .A(n396), .B(n395), .ZN(n476) );
  XNOR2_X2 U382 ( .A(KEYINPUT78), .B(G143), .ZN(n396) );
  XNOR2_X2 U383 ( .A(n570), .B(n497), .ZN(n671) );
  INV_X2 U384 ( .A(n590), .ZN(n570) );
  INV_X2 U385 ( .A(G953), .ZN(n738) );
  AND2_X1 U386 ( .A1(n364), .A2(n601), .ZN(n361) );
  NOR2_X1 U387 ( .A1(n735), .A2(n354), .ZN(n367) );
  AND2_X1 U388 ( .A1(n358), .A2(n540), .ZN(n357) );
  XNOR2_X1 U389 ( .A(n703), .B(KEYINPUT119), .ZN(n704) );
  XNOR2_X1 U390 ( .A(n732), .B(n414), .ZN(n449) );
  NAND2_X1 U391 ( .A1(n738), .A2(G224), .ZN(n379) );
  XNOR2_X2 U392 ( .A(n409), .B(n408), .ZN(n506) );
  XNOR2_X1 U393 ( .A(KEYINPUT69), .B(KEYINPUT3), .ZN(n391) );
  INV_X1 U394 ( .A(G237), .ZN(n398) );
  INV_X1 U395 ( .A(KEYINPUT45), .ZN(n355) );
  INV_X1 U396 ( .A(G128), .ZN(n395) );
  NAND2_X1 U397 ( .A1(n400), .A2(G214), .ZN(n670) );
  INV_X1 U398 ( .A(KEYINPUT0), .ZN(n408) );
  OR2_X1 U399 ( .A1(n605), .A2(G902), .ZN(n451) );
  XNOR2_X1 U400 ( .A(G119), .B(G128), .ZN(n427) );
  AND2_X1 U401 ( .A1(n495), .A2(n671), .ZN(n386) );
  XNOR2_X1 U402 ( .A(KEYINPUT15), .B(G902), .ZN(n600) );
  XOR2_X1 U403 ( .A(G116), .B(G113), .Z(n392) );
  XNOR2_X1 U404 ( .A(n391), .B(n390), .ZN(n376) );
  INV_X1 U405 ( .A(G119), .ZN(n390) );
  XOR2_X1 U406 ( .A(G104), .B(G143), .Z(n466) );
  XNOR2_X1 U407 ( .A(KEYINPUT66), .B(G101), .ZN(n413) );
  INV_X1 U408 ( .A(KEYINPUT4), .ZN(n382) );
  NAND2_X1 U409 ( .A1(G234), .A2(G237), .ZN(n403) );
  NAND2_X1 U410 ( .A1(n663), .A2(n370), .ZN(n664) );
  INV_X1 U411 ( .A(G902), .ZN(n483) );
  XNOR2_X1 U412 ( .A(n442), .B(n372), .ZN(n715) );
  XNOR2_X1 U413 ( .A(n415), .B(n373), .ZN(n372) );
  XNOR2_X1 U414 ( .A(n374), .B(KEYINPUT16), .ZN(n373) );
  INV_X1 U415 ( .A(G122), .ZN(n374) );
  XOR2_X1 U416 ( .A(KEYINPUT7), .B(G107), .Z(n478) );
  XNOR2_X1 U417 ( .A(n375), .B(G110), .ZN(n415) );
  XNOR2_X1 U418 ( .A(G104), .B(G107), .ZN(n375) );
  INV_X1 U419 ( .A(n735), .ZN(n368) );
  INV_X1 U420 ( .A(KEYINPUT85), .ZN(n401) );
  NOR2_X1 U421 ( .A1(n656), .A2(n370), .ZN(n529) );
  AND2_X1 U422 ( .A1(n532), .A2(n547), .ZN(n495) );
  XNOR2_X1 U423 ( .A(n494), .B(n493), .ZN(n387) );
  XNOR2_X1 U424 ( .A(n371), .B(KEYINPUT99), .ZN(n551) );
  BUF_X1 U425 ( .A(n506), .Z(n534) );
  BUF_X1 U426 ( .A(n371), .Z(n370) );
  XNOR2_X1 U427 ( .A(n433), .B(n731), .ZN(n710) );
  XNOR2_X1 U428 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U429 ( .A(n614), .B(n613), .ZN(n615) );
  AND2_X1 U430 ( .A1(n609), .A2(n362), .ZN(n714) );
  AND2_X1 U431 ( .A1(n380), .A2(n527), .ZN(n629) );
  XNOR2_X1 U432 ( .A(n381), .B(n526), .ZN(n380) );
  XNOR2_X1 U433 ( .A(n376), .B(n392), .ZN(n442) );
  OR2_X1 U434 ( .A1(n645), .A2(n502), .ZN(n351) );
  XOR2_X1 U435 ( .A(KEYINPUT88), .B(KEYINPUT18), .Z(n352) );
  AND2_X1 U436 ( .A1(n645), .A2(n502), .ZN(n353) );
  AND2_X1 U437 ( .A1(n603), .A2(n654), .ZN(n354) );
  INV_X2 U438 ( .A(n720), .ZN(n369) );
  XNOR2_X2 U439 ( .A(n356), .B(n355), .ZN(n720) );
  NAND2_X1 U440 ( .A1(n357), .A2(n541), .ZN(n356) );
  NAND2_X1 U441 ( .A1(n544), .A2(KEYINPUT44), .ZN(n358) );
  XNOR2_X1 U442 ( .A(n366), .B(n715), .ZN(n623) );
  NAND2_X1 U443 ( .A1(n623), .A2(n600), .ZN(n365) );
  XNOR2_X2 U444 ( .A(n359), .B(n604), .ZN(n702) );
  NAND2_X1 U445 ( .A1(n361), .A2(n363), .ZN(n359) );
  XNOR2_X2 U446 ( .A(n499), .B(n498), .ZN(n592) );
  XNOR2_X1 U447 ( .A(n429), .B(n428), .ZN(n433) );
  NAND2_X1 U448 ( .A1(n528), .A2(n554), .ZN(n488) );
  XNOR2_X1 U449 ( .A(n377), .B(n394), .ZN(n397) );
  NAND2_X1 U450 ( .A1(n655), .A2(n599), .ZN(n363) );
  NAND2_X2 U451 ( .A1(n369), .A2(n368), .ZN(n655) );
  NAND2_X1 U452 ( .A1(n369), .A2(n367), .ZN(n364) );
  XNOR2_X2 U453 ( .A(n365), .B(n399), .ZN(n496) );
  XNOR2_X1 U454 ( .A(n397), .B(n412), .ZN(n366) );
  XNOR2_X2 U455 ( .A(n371), .B(KEYINPUT6), .ZN(n563) );
  AND2_X1 U456 ( .A1(n532), .A2(n370), .ZN(n533) );
  XNOR2_X2 U457 ( .A(n451), .B(n450), .ZN(n371) );
  XNOR2_X1 U458 ( .A(n378), .B(n352), .ZN(n377) );
  NOR2_X1 U459 ( .A1(n514), .A2(n563), .ZN(n381) );
  XNOR2_X2 U460 ( .A(n412), .B(n411), .ZN(n732) );
  XNOR2_X2 U461 ( .A(n476), .B(n382), .ZN(n412) );
  NAND2_X1 U462 ( .A1(n384), .A2(n383), .ZN(n558) );
  NAND2_X1 U463 ( .A1(n592), .A2(n502), .ZN(n383) );
  NOR2_X1 U464 ( .A1(n385), .A2(n353), .ZN(n384) );
  NOR2_X1 U465 ( .A1(n592), .A2(n351), .ZN(n385) );
  NAND2_X1 U466 ( .A1(n558), .A2(n745), .ZN(n560) );
  NAND2_X1 U467 ( .A1(n387), .A2(n495), .ZN(n572) );
  NAND2_X1 U468 ( .A1(n386), .A2(n387), .ZN(n499) );
  BUF_X1 U469 ( .A(n702), .Z(n708) );
  XOR2_X1 U470 ( .A(KEYINPUT19), .B(KEYINPUT73), .Z(n388) );
  AND2_X1 U471 ( .A1(n581), .A2(n580), .ZN(n389) );
  INV_X1 U472 ( .A(KEYINPUT46), .ZN(n559) );
  INV_X1 U473 ( .A(KEYINPUT17), .ZN(n393) );
  INV_X1 U474 ( .A(KEYINPUT77), .ZN(n508) );
  INV_X1 U475 ( .A(KEYINPUT24), .ZN(n426) );
  BUF_X1 U476 ( .A(n476), .Z(n480) );
  INV_X1 U477 ( .A(n431), .ZN(n432) );
  XNOR2_X1 U478 ( .A(n469), .B(n432), .ZN(n731) );
  INV_X1 U479 ( .A(KEYINPUT30), .ZN(n493) );
  INV_X1 U480 ( .A(KEYINPUT32), .ZN(n512) );
  XNOR2_X1 U481 ( .A(n413), .B(n430), .ZN(n394) );
  NAND2_X1 U482 ( .A1(n483), .A2(n398), .ZN(n400) );
  AND2_X1 U483 ( .A1(n400), .A2(G210), .ZN(n399) );
  NAND2_X2 U484 ( .A1(n496), .A2(n670), .ZN(n402) );
  XNOR2_X2 U485 ( .A(n402), .B(n401), .ZN(n564) );
  XNOR2_X1 U486 ( .A(n564), .B(n388), .ZN(n573) );
  XNOR2_X1 U487 ( .A(n403), .B(KEYINPUT14), .ZN(n404) );
  NAND2_X1 U488 ( .A1(G952), .A2(n404), .ZN(n684) );
  OR2_X1 U489 ( .A1(n684), .A2(n362), .ZN(n491) );
  NOR2_X1 U490 ( .A1(G898), .A2(n738), .ZN(n718) );
  NAND2_X1 U491 ( .A1(n404), .A2(G902), .ZN(n405) );
  XNOR2_X1 U492 ( .A(n405), .B(KEYINPUT89), .ZN(n489) );
  NAND2_X1 U493 ( .A1(n718), .A2(n489), .ZN(n406) );
  NAND2_X1 U494 ( .A1(n491), .A2(n406), .ZN(n407) );
  NAND2_X1 U495 ( .A1(n573), .A2(n407), .ZN(n409) );
  XNOR2_X1 U496 ( .A(G134), .B(G131), .ZN(n410) );
  XNOR2_X1 U497 ( .A(n410), .B(KEYINPUT67), .ZN(n411) );
  XNOR2_X1 U498 ( .A(n413), .B(G146), .ZN(n414) );
  XOR2_X1 U499 ( .A(G137), .B(G140), .Z(n431) );
  XOR2_X1 U500 ( .A(n415), .B(n431), .Z(n419) );
  NAND2_X1 U501 ( .A1(G227), .A2(n738), .ZN(n416) );
  XNOR2_X1 U502 ( .A(KEYINPUT74), .B(n416), .ZN(n417) );
  XNOR2_X1 U503 ( .A(n417), .B(KEYINPUT90), .ZN(n418) );
  XNOR2_X1 U504 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U505 ( .A(n449), .B(n420), .ZN(n697) );
  OR2_X1 U506 ( .A1(n697), .A2(G902), .ZN(n421) );
  XNOR2_X2 U507 ( .A(n421), .B(G469), .ZN(n554) );
  XNOR2_X2 U508 ( .A(n554), .B(KEYINPUT1), .ZN(n567) );
  XOR2_X1 U509 ( .A(G110), .B(KEYINPUT23), .Z(n425) );
  XOR2_X1 U510 ( .A(KEYINPUT80), .B(KEYINPUT8), .Z(n423) );
  NAND2_X1 U511 ( .A1(G234), .A2(n738), .ZN(n422) );
  XNOR2_X1 U512 ( .A(n423), .B(n422), .ZN(n473) );
  NAND2_X1 U513 ( .A1(n473), .A2(G221), .ZN(n424) );
  XNOR2_X1 U514 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U515 ( .A(n430), .B(KEYINPUT10), .Z(n469) );
  XOR2_X1 U516 ( .A(KEYINPUT91), .B(KEYINPUT25), .Z(n437) );
  NAND2_X1 U517 ( .A1(n600), .A2(G234), .ZN(n434) );
  XNOR2_X1 U518 ( .A(n434), .B(KEYINPUT92), .ZN(n435) );
  XNOR2_X1 U519 ( .A(KEYINPUT20), .B(n435), .ZN(n440) );
  NAND2_X1 U520 ( .A1(G217), .A2(n440), .ZN(n436) );
  XOR2_X1 U521 ( .A(n437), .B(n436), .Z(n438) );
  XNOR2_X2 U522 ( .A(n439), .B(n438), .ZN(n660) );
  NAND2_X1 U523 ( .A1(n440), .A2(G221), .ZN(n441) );
  XNOR2_X1 U524 ( .A(n441), .B(KEYINPUT21), .ZN(n661) );
  AND2_X1 U525 ( .A1(n567), .A2(n528), .ZN(n452) );
  NAND2_X1 U526 ( .A1(n464), .A2(G210), .ZN(n444) );
  XNOR2_X1 U527 ( .A(KEYINPUT5), .B(G137), .ZN(n443) );
  XNOR2_X1 U528 ( .A(n444), .B(n443), .ZN(n446) );
  XNOR2_X1 U529 ( .A(KEYINPUT72), .B(KEYINPUT94), .ZN(n445) );
  XNOR2_X1 U530 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U531 ( .A(n442), .B(n447), .ZN(n448) );
  XNOR2_X1 U532 ( .A(n449), .B(n448), .ZN(n605) );
  XNOR2_X1 U533 ( .A(KEYINPUT95), .B(G472), .ZN(n450) );
  NAND2_X1 U534 ( .A1(n452), .A2(n563), .ZN(n455) );
  XNOR2_X1 U535 ( .A(KEYINPUT100), .B(KEYINPUT33), .ZN(n453) );
  XNOR2_X1 U536 ( .A(n453), .B(KEYINPUT70), .ZN(n454) );
  XNOR2_X2 U537 ( .A(n455), .B(n454), .ZN(n686) );
  NAND2_X1 U538 ( .A1(n534), .A2(n686), .ZN(n457) );
  INV_X1 U539 ( .A(KEYINPUT34), .ZN(n456) );
  XNOR2_X1 U540 ( .A(n457), .B(n456), .ZN(n485) );
  XOR2_X1 U541 ( .A(KEYINPUT96), .B(KEYINPUT12), .Z(n459) );
  XNOR2_X1 U542 ( .A(G113), .B(G122), .ZN(n458) );
  XNOR2_X1 U543 ( .A(n459), .B(n458), .ZN(n463) );
  XOR2_X1 U544 ( .A(KEYINPUT97), .B(KEYINPUT11), .Z(n461) );
  XNOR2_X1 U545 ( .A(G131), .B(G140), .ZN(n460) );
  XNOR2_X1 U546 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U547 ( .A(n463), .B(n462), .ZN(n468) );
  NAND2_X1 U548 ( .A1(G214), .A2(n464), .ZN(n465) );
  XNOR2_X1 U549 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U550 ( .A(n468), .B(n467), .ZN(n470) );
  XNOR2_X1 U551 ( .A(n470), .B(n469), .ZN(n614) );
  NAND2_X1 U552 ( .A1(n614), .A2(n483), .ZN(n472) );
  XOR2_X1 U553 ( .A(KEYINPUT13), .B(G475), .Z(n471) );
  XNOR2_X1 U554 ( .A(n472), .B(n471), .ZN(n535) );
  XOR2_X1 U555 ( .A(G134), .B(KEYINPUT9), .Z(n475) );
  NAND2_X1 U556 ( .A1(G217), .A2(n473), .ZN(n474) );
  XNOR2_X1 U557 ( .A(n475), .B(n474), .ZN(n482) );
  XNOR2_X1 U558 ( .A(G116), .B(G122), .ZN(n477) );
  XNOR2_X1 U559 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U560 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U561 ( .A(n482), .B(n481), .ZN(n703) );
  NAND2_X1 U562 ( .A1(n703), .A2(n483), .ZN(n484) );
  XNOR2_X1 U563 ( .A(n484), .B(G478), .ZN(n503) );
  AND2_X1 U564 ( .A1(n535), .A2(n503), .ZN(n569) );
  NAND2_X1 U565 ( .A1(n485), .A2(n569), .ZN(n487) );
  XNOR2_X1 U566 ( .A(KEYINPUT75), .B(KEYINPUT35), .ZN(n486) );
  XNOR2_X2 U567 ( .A(n487), .B(n486), .ZN(n542) );
  XNOR2_X1 U568 ( .A(n542), .B(G122), .ZN(G24) );
  XNOR2_X1 U569 ( .A(n488), .B(KEYINPUT93), .ZN(n532) );
  NAND2_X1 U570 ( .A1(n362), .A2(n489), .ZN(n490) );
  OR2_X1 U571 ( .A1(n490), .A2(G900), .ZN(n492) );
  NAND2_X1 U572 ( .A1(n492), .A2(n491), .ZN(n547) );
  NAND2_X1 U573 ( .A1(n551), .A2(n670), .ZN(n494) );
  INV_X1 U574 ( .A(n496), .ZN(n590) );
  XNOR2_X1 U575 ( .A(KEYINPUT71), .B(KEYINPUT38), .ZN(n497) );
  INV_X1 U576 ( .A(KEYINPUT39), .ZN(n498) );
  INV_X1 U577 ( .A(n503), .ZN(n536) );
  NAND2_X1 U578 ( .A1(n535), .A2(n536), .ZN(n645) );
  XNOR2_X1 U579 ( .A(KEYINPUT105), .B(KEYINPUT40), .ZN(n501) );
  INV_X1 U580 ( .A(KEYINPUT104), .ZN(n500) );
  XNOR2_X1 U581 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U582 ( .A(n558), .B(G131), .ZN(G33) );
  NOR2_X1 U583 ( .A1(n503), .A2(n535), .ZN(n504) );
  XOR2_X1 U584 ( .A(n504), .B(KEYINPUT98), .Z(n673) );
  NOR2_X1 U585 ( .A1(n661), .A2(n673), .ZN(n505) );
  NAND2_X1 U586 ( .A1(n506), .A2(n505), .ZN(n507) );
  XNOR2_X2 U587 ( .A(n507), .B(KEYINPUT22), .ZN(n514) );
  NAND2_X1 U588 ( .A1(n567), .A2(n660), .ZN(n510) );
  XNOR2_X1 U589 ( .A(n563), .B(n508), .ZN(n509) );
  NOR2_X2 U590 ( .A1(n514), .A2(n511), .ZN(n513) );
  XNOR2_X1 U591 ( .A(n513), .B(n512), .ZN(n742) );
  INV_X1 U592 ( .A(n514), .ZN(n518) );
  INV_X1 U593 ( .A(n660), .ZN(n515) );
  OR2_X1 U594 ( .A1(n567), .A2(n515), .ZN(n516) );
  NOR2_X1 U595 ( .A1(n516), .A2(n551), .ZN(n517) );
  NAND2_X1 U596 ( .A1(n518), .A2(n517), .ZN(n636) );
  NAND2_X1 U597 ( .A1(n742), .A2(n636), .ZN(n522) );
  INV_X1 U598 ( .A(n522), .ZN(n543) );
  INV_X1 U599 ( .A(KEYINPUT44), .ZN(n519) );
  AND2_X1 U600 ( .A1(n519), .A2(KEYINPUT84), .ZN(n520) );
  NAND2_X1 U601 ( .A1(n543), .A2(n520), .ZN(n524) );
  INV_X1 U602 ( .A(KEYINPUT84), .ZN(n521) );
  NAND2_X1 U603 ( .A1(n522), .A2(n521), .ZN(n523) );
  NAND2_X1 U604 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U605 ( .A1(n525), .A2(n542), .ZN(n541) );
  INV_X1 U606 ( .A(KEYINPUT83), .ZN(n526) );
  NOR2_X1 U607 ( .A1(n567), .A2(n660), .ZN(n527) );
  INV_X1 U608 ( .A(n528), .ZN(n656) );
  AND2_X1 U609 ( .A1(n567), .A2(n529), .ZN(n666) );
  NAND2_X1 U610 ( .A1(n534), .A2(n666), .ZN(n531) );
  INV_X1 U611 ( .A(KEYINPUT31), .ZN(n530) );
  XNOR2_X1 U612 ( .A(n531), .B(n530), .ZN(n648) );
  NAND2_X1 U613 ( .A1(n534), .A2(n533), .ZN(n631) );
  NAND2_X1 U614 ( .A1(n648), .A2(n631), .ZN(n538) );
  OR2_X1 U615 ( .A1(n536), .A2(n535), .ZN(n649) );
  AND2_X1 U616 ( .A1(n645), .A2(n649), .ZN(n675) );
  XNOR2_X1 U617 ( .A(n675), .B(KEYINPUT79), .ZN(n537) );
  AND2_X1 U618 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U619 ( .A1(n629), .A2(n539), .ZN(n540) );
  NAND2_X1 U620 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U621 ( .A1(n670), .A2(n671), .ZN(n545) );
  XNOR2_X1 U622 ( .A(KEYINPUT106), .B(n545), .ZN(n674) );
  NOR2_X1 U623 ( .A1(n674), .A2(n673), .ZN(n546) );
  XNOR2_X1 U624 ( .A(n546), .B(KEYINPUT41), .ZN(n685) );
  INV_X1 U625 ( .A(n547), .ZN(n548) );
  NOR2_X1 U626 ( .A1(n548), .A2(n661), .ZN(n549) );
  XNOR2_X1 U627 ( .A(KEYINPUT68), .B(n549), .ZN(n550) );
  AND2_X1 U628 ( .A1(n660), .A2(n550), .ZN(n561) );
  NAND2_X1 U629 ( .A1(n551), .A2(n561), .ZN(n553) );
  XNOR2_X1 U630 ( .A(KEYINPUT103), .B(KEYINPUT28), .ZN(n552) );
  XNOR2_X1 U631 ( .A(n553), .B(n552), .ZN(n555) );
  NAND2_X1 U632 ( .A1(n555), .A2(n554), .ZN(n575) );
  NOR2_X1 U633 ( .A1(n685), .A2(n575), .ZN(n557) );
  XNOR2_X1 U634 ( .A(KEYINPUT107), .B(KEYINPUT42), .ZN(n556) );
  XNOR2_X1 U635 ( .A(n557), .B(n556), .ZN(n745) );
  XNOR2_X1 U636 ( .A(n560), .B(n559), .ZN(n582) );
  INV_X1 U637 ( .A(n645), .ZN(n642) );
  AND2_X1 U638 ( .A1(n561), .A2(n642), .ZN(n562) );
  AND2_X1 U639 ( .A1(n563), .A2(n562), .ZN(n585) );
  INV_X1 U640 ( .A(n585), .ZN(n565) );
  NOR2_X1 U641 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U642 ( .A(KEYINPUT36), .B(n566), .Z(n568) );
  INV_X1 U643 ( .A(n567), .ZN(n657) );
  NOR2_X1 U644 ( .A1(n568), .A2(n657), .ZN(n651) );
  NAND2_X1 U645 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U646 ( .A1(n572), .A2(n571), .ZN(n641) );
  NOR2_X1 U647 ( .A1(n651), .A2(n641), .ZN(n581) );
  INV_X1 U648 ( .A(n573), .ZN(n574) );
  NOR2_X1 U649 ( .A1(n575), .A2(n574), .ZN(n643) );
  OR2_X1 U650 ( .A1(n643), .A2(KEYINPUT47), .ZN(n579) );
  NOR2_X1 U651 ( .A1(KEYINPUT47), .A2(KEYINPUT79), .ZN(n576) );
  XNOR2_X1 U652 ( .A(n576), .B(n675), .ZN(n577) );
  NAND2_X1 U653 ( .A1(n643), .A2(n577), .ZN(n578) );
  NAND2_X1 U654 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U655 ( .A1(n582), .A2(n389), .ZN(n584) );
  INV_X1 U656 ( .A(KEYINPUT48), .ZN(n583) );
  XNOR2_X1 U657 ( .A(n584), .B(n583), .ZN(n597) );
  NAND2_X1 U658 ( .A1(n585), .A2(n670), .ZN(n586) );
  XNOR2_X1 U659 ( .A(KEYINPUT101), .B(n586), .ZN(n587) );
  NAND2_X1 U660 ( .A1(n587), .A2(n657), .ZN(n589) );
  XNOR2_X1 U661 ( .A(KEYINPUT102), .B(KEYINPUT43), .ZN(n588) );
  XNOR2_X1 U662 ( .A(n589), .B(n588), .ZN(n591) );
  NAND2_X1 U663 ( .A1(n591), .A2(n590), .ZN(n653) );
  OR2_X1 U664 ( .A1(n592), .A2(n649), .ZN(n594) );
  INV_X1 U665 ( .A(KEYINPUT108), .ZN(n593) );
  XNOR2_X1 U666 ( .A(n594), .B(n593), .ZN(n744) );
  INV_X1 U667 ( .A(n744), .ZN(n595) );
  AND2_X1 U668 ( .A1(n653), .A2(n595), .ZN(n596) );
  NAND2_X1 U669 ( .A1(n597), .A2(n596), .ZN(n735) );
  INV_X1 U670 ( .A(KEYINPUT2), .ZN(n654) );
  INV_X1 U671 ( .A(KEYINPUT81), .ZN(n598) );
  AND2_X1 U672 ( .A1(n654), .A2(n598), .ZN(n599) );
  INV_X1 U673 ( .A(n600), .ZN(n602) );
  OR2_X1 U674 ( .A1(KEYINPUT81), .A2(n602), .ZN(n601) );
  NAND2_X1 U675 ( .A1(n602), .A2(KEYINPUT81), .ZN(n603) );
  INV_X1 U676 ( .A(KEYINPUT64), .ZN(n604) );
  NAND2_X1 U677 ( .A1(n702), .A2(G472), .ZN(n608) );
  XOR2_X1 U678 ( .A(KEYINPUT109), .B(KEYINPUT62), .Z(n606) );
  XNOR2_X1 U679 ( .A(n605), .B(n606), .ZN(n607) );
  XNOR2_X1 U680 ( .A(n608), .B(n607), .ZN(n610) );
  INV_X1 U681 ( .A(G952), .ZN(n609) );
  NOR2_X2 U682 ( .A1(n610), .A2(n714), .ZN(n612) );
  XOR2_X1 U683 ( .A(KEYINPUT110), .B(KEYINPUT63), .Z(n611) );
  XNOR2_X1 U684 ( .A(n612), .B(n611), .ZN(G57) );
  NAND2_X1 U685 ( .A1(n702), .A2(G475), .ZN(n616) );
  XOR2_X1 U686 ( .A(KEYINPUT65), .B(KEYINPUT59), .Z(n613) );
  XNOR2_X1 U687 ( .A(n616), .B(n615), .ZN(n617) );
  NOR2_X2 U688 ( .A1(n617), .A2(n714), .ZN(n619) );
  XNOR2_X1 U689 ( .A(KEYINPUT118), .B(KEYINPUT60), .ZN(n618) );
  XNOR2_X1 U690 ( .A(n619), .B(n618), .ZN(G60) );
  NAND2_X1 U691 ( .A1(n702), .A2(G210), .ZN(n625) );
  XOR2_X1 U692 ( .A(KEYINPUT87), .B(KEYINPUT54), .Z(n621) );
  XNOR2_X1 U693 ( .A(KEYINPUT55), .B(KEYINPUT86), .ZN(n620) );
  XNOR2_X1 U694 ( .A(n621), .B(n620), .ZN(n622) );
  XNOR2_X1 U695 ( .A(n623), .B(n622), .ZN(n624) );
  XNOR2_X1 U696 ( .A(n625), .B(n624), .ZN(n626) );
  NOR2_X2 U697 ( .A1(n626), .A2(n714), .ZN(n628) );
  XNOR2_X1 U698 ( .A(KEYINPUT82), .B(KEYINPUT56), .ZN(n627) );
  XNOR2_X1 U699 ( .A(n628), .B(n627), .ZN(G51) );
  XOR2_X1 U700 ( .A(G101), .B(n629), .Z(G3) );
  NOR2_X1 U701 ( .A1(n645), .A2(n631), .ZN(n630) );
  XOR2_X1 U702 ( .A(G104), .B(n630), .Z(G6) );
  NOR2_X1 U703 ( .A1(n631), .A2(n649), .ZN(n635) );
  XOR2_X1 U704 ( .A(KEYINPUT111), .B(KEYINPUT26), .Z(n633) );
  XNOR2_X1 U705 ( .A(G107), .B(KEYINPUT27), .ZN(n632) );
  XNOR2_X1 U706 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U707 ( .A(n635), .B(n634), .ZN(G9) );
  XNOR2_X1 U708 ( .A(G110), .B(n636), .ZN(G12) );
  XOR2_X1 U709 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n639) );
  INV_X1 U710 ( .A(n649), .ZN(n637) );
  NAND2_X1 U711 ( .A1(n643), .A2(n637), .ZN(n638) );
  XNOR2_X1 U712 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U713 ( .A(G128), .B(n640), .ZN(G30) );
  XOR2_X1 U714 ( .A(G143), .B(n641), .Z(G45) );
  NAND2_X1 U715 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U716 ( .A(n644), .B(G146), .ZN(G48) );
  NOR2_X1 U717 ( .A1(n645), .A2(n648), .ZN(n647) );
  XNOR2_X1 U718 ( .A(G113), .B(KEYINPUT113), .ZN(n646) );
  XNOR2_X1 U719 ( .A(n647), .B(n646), .ZN(G15) );
  NOR2_X1 U720 ( .A1(n649), .A2(n648), .ZN(n650) );
  XOR2_X1 U721 ( .A(G116), .B(n650), .Z(G18) );
  XNOR2_X1 U722 ( .A(n651), .B(G125), .ZN(n652) );
  XNOR2_X1 U723 ( .A(n652), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U724 ( .A(G140), .B(n653), .ZN(G42) );
  XNOR2_X1 U725 ( .A(n655), .B(n654), .ZN(n692) );
  NAND2_X1 U726 ( .A1(n657), .A2(n656), .ZN(n659) );
  XOR2_X1 U727 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n658) );
  XNOR2_X1 U728 ( .A(n659), .B(n658), .ZN(n665) );
  NAND2_X1 U729 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U730 ( .A(KEYINPUT49), .B(n662), .Z(n663) );
  NOR2_X1 U731 ( .A1(n665), .A2(n664), .ZN(n667) );
  OR2_X1 U732 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U733 ( .A(KEYINPUT51), .B(n668), .ZN(n669) );
  NOR2_X1 U734 ( .A1(n685), .A2(n669), .ZN(n681) );
  NOR2_X1 U735 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U736 ( .A1(n673), .A2(n672), .ZN(n677) );
  NOR2_X1 U737 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U738 ( .A1(n677), .A2(n676), .ZN(n679) );
  INV_X1 U739 ( .A(n686), .ZN(n678) );
  NOR2_X1 U740 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U741 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U742 ( .A(n682), .B(KEYINPUT52), .ZN(n683) );
  NOR2_X1 U743 ( .A1(n684), .A2(n683), .ZN(n690) );
  INV_X1 U744 ( .A(n685), .ZN(n687) );
  NAND2_X1 U745 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U746 ( .A(n688), .B(KEYINPUT115), .ZN(n689) );
  NOR2_X1 U747 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U748 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U749 ( .A1(n693), .A2(n362), .ZN(n694) );
  XNOR2_X1 U750 ( .A(n694), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U751 ( .A1(n708), .A2(G469), .ZN(n700) );
  XOR2_X1 U752 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n696) );
  XNOR2_X1 U753 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n695) );
  XNOR2_X1 U754 ( .A(n696), .B(n695), .ZN(n698) );
  XOR2_X1 U755 ( .A(n698), .B(n697), .Z(n699) );
  XNOR2_X1 U756 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U757 ( .A1(n714), .A2(n701), .ZN(G54) );
  NAND2_X1 U758 ( .A1(n702), .A2(G478), .ZN(n705) );
  XNOR2_X1 U759 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X2 U760 ( .A1(n706), .A2(n714), .ZN(n707) );
  XNOR2_X1 U761 ( .A(n707), .B(KEYINPUT120), .ZN(G63) );
  NAND2_X1 U762 ( .A1(n708), .A2(G217), .ZN(n712) );
  INV_X1 U763 ( .A(KEYINPUT121), .ZN(n709) );
  XNOR2_X1 U764 ( .A(n710), .B(n709), .ZN(n711) );
  XNOR2_X1 U765 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U766 ( .A1(n714), .A2(n713), .ZN(G66) );
  XOR2_X1 U767 ( .A(KEYINPUT125), .B(KEYINPUT124), .Z(n717) );
  XNOR2_X1 U768 ( .A(G101), .B(n715), .ZN(n716) );
  XNOR2_X1 U769 ( .A(n717), .B(n716), .ZN(n719) );
  NOR2_X1 U770 ( .A1(n719), .A2(n718), .ZN(n730) );
  BUF_X1 U771 ( .A(n720), .Z(n721) );
  NOR2_X1 U772 ( .A1(n721), .A2(n362), .ZN(n722) );
  XOR2_X1 U773 ( .A(KEYINPUT123), .B(n722), .Z(n727) );
  NAND2_X1 U774 ( .A1(n362), .A2(G224), .ZN(n723) );
  XNOR2_X1 U775 ( .A(KEYINPUT61), .B(n723), .ZN(n724) );
  NAND2_X1 U776 ( .A1(n724), .A2(G898), .ZN(n725) );
  XOR2_X1 U777 ( .A(n725), .B(KEYINPUT122), .Z(n726) );
  NOR2_X1 U778 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U779 ( .A(KEYINPUT126), .B(n728), .Z(n729) );
  XNOR2_X1 U780 ( .A(n730), .B(n729), .ZN(G69) );
  XNOR2_X1 U781 ( .A(n732), .B(n731), .ZN(n736) );
  XNOR2_X1 U782 ( .A(n736), .B(G227), .ZN(n733) );
  NAND2_X1 U783 ( .A1(n733), .A2(G900), .ZN(n734) );
  NAND2_X1 U784 ( .A1(n734), .A2(n362), .ZN(n741) );
  XOR2_X1 U785 ( .A(n736), .B(KEYINPUT127), .Z(n737) );
  XNOR2_X1 U786 ( .A(n735), .B(n737), .ZN(n739) );
  NAND2_X1 U787 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U788 ( .A1(n741), .A2(n740), .ZN(G72) );
  BUF_X1 U789 ( .A(n742), .Z(n743) );
  XNOR2_X1 U790 ( .A(n743), .B(G119), .ZN(G21) );
  XOR2_X1 U791 ( .A(G134), .B(n744), .Z(G36) );
  XNOR2_X1 U792 ( .A(G137), .B(n745), .ZN(G39) );
endmodule

