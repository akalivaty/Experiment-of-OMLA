//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 1 0 1 0 0 1 1 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 0 1 1 1 1 1 1 0 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n876, new_n877,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n996, new_n997, new_n998;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(KEYINPUT92), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(KEYINPUT92), .ZN(new_n204));
  AND3_X1   g003(.A1(new_n203), .A2(KEYINPUT15), .A3(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT14), .ZN(new_n206));
  INV_X1    g005(.A(G36gat), .ZN(new_n207));
  NOR3_X1   g006(.A1(new_n206), .A2(new_n207), .A3(G29gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT14), .B(G29gat), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n208), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n205), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT93), .B(G50gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n213), .A2(G43gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT94), .ZN(new_n215));
  AOI21_X1  g014(.A(KEYINPUT15), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G50gat), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n215), .B1(G43gat), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(new_n213), .B2(G43gat), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n210), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n212), .B1(new_n220), .B2(new_n205), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT17), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n223), .B1(new_n224), .B2(G1gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G1gat), .B2(new_n223), .ZN(new_n226));
  XOR2_X1   g025(.A(new_n226), .B(G8gat), .Z(new_n227));
  INV_X1    g026(.A(KEYINPUT17), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n212), .B(new_n228), .C1(new_n205), .C2(new_n220), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n222), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G229gat), .A2(G233gat), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n221), .A2(new_n227), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT18), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n221), .B(new_n227), .ZN(new_n236));
  XOR2_X1   g035(.A(new_n231), .B(KEYINPUT13), .Z(new_n237));
  AOI22_X1  g036(.A1(new_n233), .A2(new_n234), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G113gat), .B(G141gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G169gat), .B(G197gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(KEYINPUT12), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n235), .A2(new_n238), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n244), .B1(new_n235), .B2(new_n238), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT6), .ZN(new_n250));
  INV_X1    g049(.A(G141gat), .ZN(new_n251));
  INV_X1    g050(.A(G148gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G141gat), .A2(G148gat), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OR2_X1    g054(.A1(G155gat), .A2(G162gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(G155gat), .A2(G162gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT77), .B(G155gat), .ZN(new_n259));
  INV_X1    g058(.A(G162gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT2), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n255), .B(new_n258), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n256), .A2(KEYINPUT75), .A3(new_n257), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT75), .ZN(new_n265));
  AND2_X1   g064(.A1(G155gat), .A2(G162gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(G155gat), .A2(G162gat), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT76), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n253), .B(new_n254), .C1(new_n266), .C2(new_n262), .ZN(new_n271));
  AND3_X1   g070(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n270), .B1(new_n269), .B2(new_n271), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n263), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT1), .ZN(new_n276));
  INV_X1    g075(.A(G113gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n277), .A2(G120gat), .ZN(new_n278));
  INV_X1    g077(.A(G120gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n279), .A2(G113gat), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n275), .B(new_n276), .C1(new_n278), .C2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G127gat), .B(G134gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(KEYINPUT68), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT68), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n284), .B(new_n276), .C1(new_n278), .C2(new_n280), .ZN(new_n285));
  INV_X1    g084(.A(new_n282), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n279), .A2(G113gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n277), .A2(G120gat), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT1), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n284), .B1(new_n290), .B2(new_n275), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n283), .B1(new_n287), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT4), .B1(new_n274), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n258), .A2(new_n253), .A3(new_n254), .ZN(new_n295));
  XOR2_X1   g094(.A(KEYINPUT77), .B(G155gat), .Z(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G162gat), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n295), .B1(new_n297), .B2(KEYINPUT2), .ZN(new_n298));
  NOR3_X1   g097(.A1(new_n266), .A2(new_n267), .A3(new_n265), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT75), .B1(new_n256), .B2(new_n257), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n271), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT76), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n298), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT4), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(new_n305), .A3(new_n292), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT79), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n294), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n274), .A2(KEYINPUT3), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT3), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n310), .B(new_n263), .C1(new_n272), .C2(new_n273), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n309), .A2(new_n293), .A3(new_n311), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n304), .A2(KEYINPUT79), .A3(new_n305), .A4(new_n292), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n308), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n316), .A2(KEYINPUT5), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n294), .A2(new_n306), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n320), .A2(new_n315), .A3(new_n312), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT5), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n304), .A2(new_n292), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n274), .A2(new_n293), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n322), .B1(new_n325), .B2(new_n316), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n321), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT78), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT78), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n321), .A2(new_n326), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n319), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G1gat), .B(G29gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(KEYINPUT0), .ZN(new_n333));
  XNOR2_X1  g132(.A(G57gat), .B(G85gat), .ZN(new_n334));
  XOR2_X1   g133(.A(new_n333), .B(new_n334), .Z(new_n335));
  OAI21_X1  g134(.A(new_n250), .B1(new_n331), .B2(new_n335), .ZN(new_n336));
  OR2_X1    g135(.A1(new_n314), .A2(new_n318), .ZN(new_n337));
  AND3_X1   g136(.A1(new_n321), .A2(new_n326), .A3(new_n329), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n329), .B1(new_n321), .B2(new_n326), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n337), .B(new_n335), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT80), .B1(new_n336), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n343));
  INV_X1    g142(.A(new_n335), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT80), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n345), .A2(new_n346), .A3(new_n250), .A4(new_n340), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n343), .A2(KEYINPUT6), .A3(new_n344), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n342), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G226gat), .A2(G233gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n350), .B(KEYINPUT72), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n351), .B(KEYINPUT73), .Z(new_n352));
  AOI21_X1  g151(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(G169gat), .A2(G176gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT23), .ZN(new_n359));
  NAND2_X1  g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(G169gat), .ZN(new_n362));
  INV_X1    g161(.A(G176gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT23), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n361), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n357), .A2(new_n359), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT25), .ZN(new_n368));
  NAND2_X1  g167(.A1(G183gat), .A2(G190gat), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT65), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT24), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT24), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n369), .A2(new_n370), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT66), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n375), .B1(G183gat), .B2(G190gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n354), .A2(KEYINPUT66), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n372), .A2(new_n374), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n365), .B1(G169gat), .B2(G176gat), .ZN(new_n379));
  AND4_X1   g178(.A1(KEYINPUT25), .A2(new_n359), .A3(new_n379), .A4(new_n360), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n367), .A2(new_n368), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(G183gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT27), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT27), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(G183gat), .ZN(new_n385));
  INV_X1    g184(.A(G190gat), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n383), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AND2_X1   g186(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n387), .A2(new_n388), .B1(G183gat), .B2(G190gat), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n383), .A2(new_n385), .A3(new_n386), .ZN(new_n390));
  NOR2_X1   g189(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n364), .B1(new_n361), .B2(KEYINPUT26), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT26), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n358), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n389), .A2(new_n393), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n352), .B1(new_n381), .B2(new_n398), .ZN(new_n399));
  AND2_X1   g198(.A1(G211gat), .A2(G218gat), .ZN(new_n400));
  NOR2_X1   g199(.A1(G211gat), .A2(G218gat), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AND2_X1   g201(.A1(G197gat), .A2(G204gat), .ZN(new_n403));
  NOR2_X1   g202(.A1(G197gat), .A2(G204gat), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n402), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G211gat), .B(G218gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(G197gat), .B(G204gat), .ZN(new_n409));
  INV_X1    g208(.A(new_n406), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n380), .A2(new_n378), .ZN(new_n413));
  INV_X1    g212(.A(new_n356), .ZN(new_n414));
  NOR3_X1   g213(.A1(new_n414), .A2(new_n353), .A3(new_n354), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n359), .A2(new_n360), .A3(new_n379), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n368), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n390), .A2(new_n392), .B1(new_n394), .B2(new_n396), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n389), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT29), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n399), .B(new_n412), .C1(new_n421), .C2(new_n351), .ZN(new_n422));
  XNOR2_X1  g221(.A(G8gat), .B(G36gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(G64gat), .B(G92gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  INV_X1    g224(.A(KEYINPUT29), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n426), .B1(new_n381), .B2(new_n398), .ZN(new_n427));
  INV_X1    g226(.A(new_n352), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n418), .A2(new_n420), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n427), .A2(new_n428), .B1(new_n351), .B2(new_n429), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n422), .B(new_n425), .C1(new_n430), .C2(new_n412), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n431), .B(KEYINPUT30), .ZN(new_n432));
  INV_X1    g231(.A(new_n422), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n413), .A2(new_n417), .B1(new_n419), .B2(new_n389), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n428), .B1(new_n434), .B2(KEYINPUT29), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n429), .A2(new_n351), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n412), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT74), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT74), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n439), .B(new_n422), .C1(new_n430), .C2(new_n412), .ZN(new_n440));
  INV_X1    g239(.A(new_n425), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n432), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n349), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT3), .B1(new_n412), .B2(new_n426), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n302), .A2(new_n303), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n446), .B1(new_n447), .B2(new_n263), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n311), .A2(new_n426), .ZN(new_n449));
  INV_X1    g248(.A(new_n412), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT82), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n452), .B1(new_n304), .B2(new_n446), .ZN(new_n453));
  NAND2_X1  g252(.A1(G228gat), .A2(G233gat), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n412), .B1(new_n311), .B2(new_n426), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n453), .B(new_n455), .C1(new_n458), .C2(new_n448), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n457), .A2(G22gat), .A3(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(KEYINPUT83), .B(G22gat), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n462), .B1(new_n457), .B2(new_n459), .ZN(new_n463));
  XNOR2_X1  g262(.A(G78gat), .B(G106gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n464), .B(new_n217), .ZN(new_n465));
  XOR2_X1   g264(.A(KEYINPUT81), .B(KEYINPUT31), .Z(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NOR3_X1   g267(.A1(new_n460), .A2(new_n463), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT84), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n457), .A2(new_n459), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n461), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n459), .A3(new_n462), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n471), .B1(new_n475), .B2(new_n468), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n457), .A2(new_n459), .A3(new_n462), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n471), .B(new_n468), .C1(new_n477), .C2(new_n463), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n470), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT85), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n468), .B1(new_n477), .B2(new_n463), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT84), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n478), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT85), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(new_n485), .A3(new_n470), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n481), .A2(KEYINPUT86), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT86), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n485), .B1(new_n484), .B2(new_n470), .ZN(new_n489));
  AOI211_X1 g288(.A(KEYINPUT85), .B(new_n469), .C1(new_n483), .C2(new_n478), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n445), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT36), .ZN(new_n493));
  INV_X1    g292(.A(G227gat), .ZN(new_n494));
  INV_X1    g293(.A(G233gat), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  XOR2_X1   g295(.A(new_n496), .B(KEYINPUT64), .Z(new_n497));
  AND3_X1   g296(.A1(new_n418), .A2(new_n292), .A3(new_n420), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n292), .B1(new_n418), .B2(new_n420), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT32), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT33), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  XOR2_X1   g302(.A(G15gat), .B(G43gat), .Z(new_n504));
  XNOR2_X1  g303(.A(G71gat), .B(G99gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n501), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n499), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n434), .A2(new_n292), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n508), .B(new_n509), .C1(new_n494), .C2(new_n495), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n498), .A2(new_n499), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n497), .A2(KEYINPUT34), .ZN(new_n512));
  AOI22_X1  g311(.A1(new_n510), .A2(KEYINPUT34), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n506), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n500), .B(KEYINPUT32), .C1(new_n502), .C2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n507), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT71), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT71), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n507), .A2(new_n513), .A3(new_n518), .A4(new_n515), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n507), .A2(new_n515), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT70), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n513), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n507), .A2(KEYINPUT70), .A3(new_n515), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n493), .B1(new_n520), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n513), .B1(new_n507), .B2(new_n515), .ZN(new_n528));
  AOI211_X1 g327(.A(KEYINPUT36), .B(new_n528), .C1(new_n517), .C2(new_n519), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n481), .A2(new_n486), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n438), .A2(KEYINPUT37), .A3(new_n440), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n441), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT90), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT90), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n532), .A2(new_n535), .A3(new_n441), .ZN(new_n536));
  OR3_X1    g335(.A1(new_n433), .A2(new_n437), .A3(KEYINPUT37), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT38), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n345), .A2(new_n250), .A3(new_n340), .ZN(new_n540));
  INV_X1    g339(.A(new_n431), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n425), .A2(KEYINPUT38), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n430), .A2(new_n412), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n544), .A2(KEYINPUT89), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n399), .B1(new_n421), .B2(new_n351), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n546), .A2(new_n450), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n544), .A2(KEYINPUT89), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n545), .B(KEYINPUT37), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n541), .B1(new_n543), .B2(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n539), .A2(new_n540), .A3(new_n348), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n345), .A2(new_n443), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT40), .ZN(new_n553));
  XOR2_X1   g352(.A(KEYINPUT87), .B(KEYINPUT39), .Z(new_n554));
  NAND3_X1  g353(.A1(new_n314), .A2(new_n316), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n335), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT39), .B1(new_n325), .B2(new_n316), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n557), .B1(new_n314), .B2(new_n316), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n553), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n314), .A2(new_n316), .ZN(new_n560));
  INV_X1    g359(.A(new_n557), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n562), .A2(KEYINPUT40), .A3(new_n335), .A4(new_n555), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT88), .B1(new_n552), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g364(.A1(new_n343), .A2(new_n344), .B1(new_n432), .B2(new_n442), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT88), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n566), .A2(new_n567), .A3(new_n559), .A4(new_n563), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n531), .A2(new_n551), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n492), .A2(new_n530), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n513), .B1(new_n521), .B2(new_n522), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n525), .A2(new_n572), .B1(new_n517), .B2(new_n519), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n573), .B1(new_n489), .B2(new_n490), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT35), .B1(new_n445), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n489), .A2(new_n490), .ZN(new_n576));
  INV_X1    g375(.A(new_n528), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n520), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n578), .A2(new_n443), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n540), .A2(new_n348), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT35), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n576), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n575), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n249), .B1(new_n571), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G134gat), .B(G162gat), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G99gat), .A2(G106gat), .ZN(new_n588));
  INV_X1    g387(.A(G85gat), .ZN(new_n589));
  INV_X1    g388(.A(G92gat), .ZN(new_n590));
  AOI22_X1  g389(.A1(KEYINPUT8), .A2(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT7), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n592), .B1(new_n589), .B2(new_n590), .ZN(new_n593));
  NAND3_X1  g392(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G99gat), .B(G106gat), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n596), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT99), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n600), .A2(new_n229), .A3(new_n222), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n221), .A2(new_n599), .ZN(new_n602));
  AND2_X1   g401(.A1(G232gat), .A2(G233gat), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n603), .A2(KEYINPUT41), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G190gat), .B(G218gat), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n607), .A2(KEYINPUT100), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n587), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  AOI211_X1 g409(.A(new_n586), .B(new_n608), .C1(new_n601), .C2(new_n605), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n603), .A2(KEYINPUT41), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT98), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n607), .A2(KEYINPUT100), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n614), .B(new_n615), .Z(new_n616));
  NAND2_X1  g415(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n616), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n618), .B1(new_n610), .B2(new_n611), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  OR2_X1    g419(.A1(G57gat), .A2(G64gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(G57gat), .A2(G64gat), .ZN(new_n622));
  AND2_X1   g421(.A1(G71gat), .A2(G78gat), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n621), .B(new_n622), .C1(new_n623), .C2(KEYINPUT9), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT95), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(G71gat), .A2(G78gat), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n624), .B(new_n626), .C1(new_n623), .C2(new_n628), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n632), .A2(KEYINPUT21), .ZN(new_n633));
  XNOR2_X1  g432(.A(G127gat), .B(G155gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT21), .ZN(new_n636));
  INV_X1    g435(.A(new_n632), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n227), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n635), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT97), .ZN(new_n641));
  NAND2_X1  g440(.A1(G231gat), .A2(G233gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT96), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n641), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G183gat), .B(G211gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n639), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G120gat), .B(G148gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(G176gat), .B(G204gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n632), .A2(new_n597), .A3(new_n598), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n651), .A2(KEYINPUT101), .A3(KEYINPUT10), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n599), .A2(new_n637), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(KEYINPUT10), .B1(new_n651), .B2(KEYINPUT101), .ZN(new_n655));
  NAND2_X1  g454(.A1(G230gat), .A2(G233gat), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n654), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n656), .B1(new_n653), .B2(new_n651), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n650), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n659), .A2(KEYINPUT102), .ZN(new_n661));
  INV_X1    g460(.A(new_n655), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n662), .A2(new_n656), .A3(new_n653), .A4(new_n652), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n650), .B1(new_n659), .B2(KEYINPUT102), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n661), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n620), .A2(new_n647), .A3(new_n666), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n349), .A2(KEYINPUT103), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n349), .A2(KEYINPUT103), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n585), .A2(new_n667), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT104), .B(G1gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(G1324gat));
  NAND2_X1  g473(.A1(new_n571), .A2(new_n584), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n248), .ZN(new_n676));
  INV_X1    g475(.A(new_n667), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n676), .A2(new_n444), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT16), .B(G8gat), .Z(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n681));
  INV_X1    g480(.A(new_n678), .ZN(new_n682));
  AOI22_X1  g481(.A1(new_n680), .A2(new_n681), .B1(new_n682), .B2(G8gat), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT106), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT42), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n684), .B1(new_n680), .B2(new_n685), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n678), .A2(KEYINPUT106), .A3(KEYINPUT42), .A4(new_n679), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n683), .A2(new_n686), .A3(new_n687), .ZN(G1325gat));
  NOR2_X1   g487(.A1(new_n676), .A2(new_n677), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT107), .B1(new_n527), .B2(new_n529), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n520), .A2(new_n493), .A3(new_n577), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT107), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n691), .B(new_n692), .C1(new_n573), .C2(new_n493), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(G15gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT108), .ZN(new_n696));
  INV_X1    g495(.A(new_n578), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n585), .A2(new_n697), .A3(new_n667), .ZN(new_n698));
  INV_X1    g497(.A(G15gat), .ZN(new_n699));
  AOI22_X1  g498(.A1(new_n689), .A2(new_n696), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT109), .ZN(G1326gat));
  NAND2_X1  g500(.A1(new_n491), .A2(new_n487), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n585), .A2(new_n703), .A3(new_n667), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT43), .B(G22gat), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1327gat));
  INV_X1    g505(.A(new_n647), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(new_n666), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n620), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n676), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n670), .A2(G29gat), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT45), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n445), .A2(new_n487), .A3(new_n491), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n690), .A2(new_n693), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n570), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n348), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n717), .B1(new_n540), .B2(KEYINPUT80), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n443), .B1(new_n718), .B2(new_n347), .ZN(new_n719));
  INV_X1    g518(.A(new_n573), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n720), .B1(new_n481), .B2(new_n486), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n581), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n576), .A2(new_n582), .ZN(new_n723));
  OAI22_X1  g522(.A1(new_n714), .A2(new_n716), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(KEYINPUT44), .B1(new_n724), .B2(new_n620), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n617), .A2(new_n619), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n729), .B1(new_n571), .B2(new_n584), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n248), .A2(new_n708), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n725), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G29gat), .B1(new_n733), .B2(new_n670), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n713), .A2(new_n734), .ZN(G1328gat));
  INV_X1    g534(.A(new_n709), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n585), .A2(new_n207), .A3(new_n443), .A4(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT46), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT110), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(new_n740));
  OR3_X1    g539(.A1(new_n737), .A2(KEYINPUT111), .A3(KEYINPUT46), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT111), .B1(new_n737), .B2(KEYINPUT46), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(G36gat), .B1(new_n733), .B2(new_n444), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n740), .A2(new_n743), .A3(new_n744), .ZN(G1329gat));
  INV_X1    g544(.A(KEYINPUT47), .ZN(new_n746));
  INV_X1    g545(.A(G43gat), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n747), .B1(new_n732), .B2(new_n694), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n578), .A2(G43gat), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n585), .A2(new_n736), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT112), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT112), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n585), .A2(new_n752), .A3(new_n736), .A4(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n746), .B1(new_n748), .B2(new_n754), .ZN(new_n755));
  AOI22_X1  g554(.A1(new_n481), .A2(new_n486), .B1(new_n565), .B2(new_n568), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n694), .B1(new_n756), .B2(new_n551), .ZN(new_n757));
  AOI22_X1  g556(.A1(new_n492), .A2(new_n757), .B1(new_n575), .B2(new_n583), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n727), .B1(new_n758), .B2(new_n726), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n675), .A2(new_n728), .ZN(new_n760));
  INV_X1    g559(.A(new_n731), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n759), .A2(new_n694), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G43gat), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n763), .A2(KEYINPUT47), .A3(new_n751), .A4(new_n753), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n755), .A2(new_n764), .ZN(G1330gat));
  NAND4_X1  g564(.A1(new_n759), .A2(new_n703), .A3(new_n760), .A4(new_n761), .ZN(new_n766));
  INV_X1    g565(.A(new_n213), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n702), .A2(new_n767), .ZN(new_n768));
  AOI22_X1  g567(.A1(new_n766), .A2(new_n767), .B1(new_n710), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n213), .B1(new_n732), .B2(new_n576), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n710), .A2(new_n768), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT48), .ZN(new_n772));
  OAI22_X1  g571(.A1(KEYINPUT48), .A2(new_n769), .B1(new_n770), .B2(new_n772), .ZN(G1331gat));
  INV_X1    g572(.A(new_n666), .ZN(new_n774));
  NOR4_X1   g573(.A1(new_n248), .A2(new_n620), .A3(new_n647), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n724), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n776), .A2(new_n670), .ZN(new_n777));
  XOR2_X1   g576(.A(new_n777), .B(G57gat), .Z(G1332gat));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n724), .A2(KEYINPUT113), .A3(new_n775), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n443), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n783), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n784));
  XNOR2_X1  g583(.A(KEYINPUT49), .B(G64gat), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n782), .A2(new_n443), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(G1333gat));
  XNOR2_X1  g586(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n780), .A2(new_n694), .A3(new_n781), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(G71gat), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n578), .A2(G71gat), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n788), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n788), .ZN(new_n795));
  AOI211_X1 g594(.A(new_n792), .B(new_n795), .C1(new_n789), .C2(G71gat), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n794), .A2(new_n796), .ZN(G1334gat));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n703), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g598(.A1(new_n248), .A2(new_n707), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n724), .A2(new_n620), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n724), .A2(KEYINPUT51), .A3(new_n620), .A4(new_n800), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n801), .A2(KEYINPUT115), .A3(new_n802), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n670), .A2(G85gat), .A3(new_n774), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n248), .A2(new_n707), .A3(new_n774), .ZN(new_n810));
  AND4_X1   g609(.A1(new_n671), .A2(new_n759), .A3(new_n760), .A4(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n809), .B1(new_n589), .B2(new_n811), .ZN(G1336gat));
  NOR3_X1   g611(.A1(new_n444), .A2(G92gat), .A3(new_n774), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n806), .A2(new_n807), .A3(new_n813), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n759), .A2(new_n443), .A3(new_n760), .A4(new_n810), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(G92gat), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n805), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n819), .A2(new_n813), .B1(new_n815), .B2(G92gat), .ZN(new_n820));
  OAI22_X1  g619(.A1(new_n814), .A2(new_n818), .B1(new_n820), .B2(new_n817), .ZN(G1337gat));
  INV_X1    g620(.A(G99gat), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n759), .A2(new_n694), .A3(new_n760), .A4(new_n810), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT116), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n825), .B1(new_n824), .B2(new_n823), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n578), .A2(G99gat), .A3(new_n774), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n806), .A2(new_n807), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(G1338gat));
  NOR3_X1   g628(.A1(new_n531), .A2(G106gat), .A3(new_n774), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n806), .A2(new_n807), .A3(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n759), .A2(new_n576), .A3(new_n760), .A4(new_n810), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(G106gat), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n759), .A2(new_n703), .A3(new_n760), .A4(new_n810), .ZN(new_n836));
  AOI22_X1  g635(.A1(new_n819), .A2(new_n830), .B1(new_n836), .B2(G106gat), .ZN(new_n837));
  OAI22_X1  g636(.A1(new_n831), .A2(new_n835), .B1(new_n837), .B2(new_n834), .ZN(G1339gat));
  OR2_X1    g637(.A1(new_n663), .A2(KEYINPUT54), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n657), .B1(new_n654), .B2(new_n655), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n840), .A2(new_n663), .A3(KEYINPUT54), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n839), .A2(new_n650), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n839), .A2(KEYINPUT55), .A3(new_n841), .A4(new_n650), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(new_n665), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n236), .A2(new_n237), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n231), .B1(new_n230), .B2(new_n232), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n243), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n245), .A2(new_n849), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n726), .A2(new_n846), .A3(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n665), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n852), .B1(new_n842), .B2(new_n843), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n853), .B(new_n845), .C1(new_n246), .C2(new_n247), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n245), .A2(new_n666), .A3(new_n849), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n620), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n647), .B1(new_n851), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n667), .A2(new_n249), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n860), .A2(new_n670), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n574), .A2(new_n443), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(G113gat), .B1(new_n864), .B2(new_n248), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n860), .A2(new_n703), .ZN(new_n866));
  AND3_X1   g665(.A1(new_n866), .A2(new_n579), .A3(new_n671), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n249), .A2(new_n277), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n865), .B1(new_n867), .B2(new_n868), .ZN(G1340gat));
  AOI21_X1  g668(.A(new_n279), .B1(new_n867), .B2(new_n666), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT117), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n870), .A2(new_n871), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n666), .A2(new_n279), .ZN(new_n874));
  OAI22_X1  g673(.A1(new_n872), .A2(new_n873), .B1(new_n863), .B2(new_n874), .ZN(G1341gat));
  NAND3_X1  g674(.A1(new_n867), .A2(G127gat), .A3(new_n707), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n876), .A2(KEYINPUT118), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(KEYINPUT118), .ZN(new_n878));
  AOI21_X1  g677(.A(G127gat), .B1(new_n864), .B2(new_n707), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(G1342gat));
  INV_X1    g679(.A(new_n867), .ZN(new_n881));
  OAI21_X1  g680(.A(G134gat), .B1(new_n881), .B2(new_n726), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT56), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n726), .A2(G134gat), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n863), .A2(new_n884), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n885), .A2(KEYINPUT119), .A3(new_n883), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT119), .B1(new_n885), .B2(new_n883), .ZN(new_n887));
  OAI221_X1 g686(.A(new_n882), .B1(new_n883), .B2(new_n885), .C1(new_n886), .C2(new_n887), .ZN(G1343gat));
  NAND2_X1  g687(.A1(new_n846), .A2(KEYINPUT120), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n853), .A2(new_n890), .A3(new_n845), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n889), .A2(new_n248), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n620), .B1(new_n892), .B2(new_n855), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n647), .B1(new_n893), .B2(new_n851), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n702), .B1(new_n894), .B2(new_n858), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(KEYINPUT57), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n859), .A2(new_n576), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT57), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT121), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n895), .A2(KEYINPUT121), .A3(KEYINPUT57), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n715), .A2(new_n444), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n670), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n900), .A2(new_n248), .A3(new_n901), .A4(new_n903), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n904), .A2(G141gat), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n694), .A2(new_n531), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n861), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n671), .A2(new_n859), .ZN(new_n909));
  INV_X1    g708(.A(new_n907), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT123), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n248), .A2(new_n251), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT122), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n908), .A2(new_n911), .A3(new_n444), .A4(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT58), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AND4_X1   g715(.A1(new_n444), .A2(new_n861), .A3(new_n907), .A4(new_n913), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n917), .B1(new_n904), .B2(G141gat), .ZN(new_n918));
  OAI22_X1  g717(.A1(new_n905), .A2(new_n916), .B1(new_n918), .B2(new_n915), .ZN(G1344gat));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n898), .B1(new_n859), .B2(new_n576), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n921), .B1(new_n895), .B2(new_n898), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n903), .A2(new_n666), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n252), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT59), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n920), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n894), .A2(new_n858), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n928), .A2(new_n898), .A3(new_n703), .ZN(new_n929));
  INV_X1    g728(.A(new_n921), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(G148gat), .B1(new_n931), .B2(new_n923), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n932), .A2(KEYINPUT124), .A3(KEYINPUT59), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n900), .A2(new_n666), .A3(new_n901), .A4(new_n903), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n252), .A2(KEYINPUT59), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n927), .A2(new_n933), .A3(new_n936), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n908), .A2(new_n911), .A3(new_n444), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n938), .A2(new_n252), .A3(new_n666), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(G1345gat));
  NAND3_X1  g739(.A1(new_n900), .A2(new_n901), .A3(new_n903), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n296), .B1(new_n941), .B2(new_n647), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n938), .A2(new_n259), .A3(new_n707), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1346gat));
  NOR3_X1   g743(.A1(new_n941), .A2(new_n260), .A3(new_n726), .ZN(new_n945));
  AOI21_X1  g744(.A(G162gat), .B1(new_n938), .B2(new_n620), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n945), .A2(new_n946), .ZN(G1347gat));
  NAND4_X1  g746(.A1(new_n866), .A2(new_n443), .A3(new_n697), .A4(new_n670), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n948), .A2(new_n362), .A3(new_n249), .ZN(new_n949));
  NOR4_X1   g748(.A1(new_n860), .A2(new_n671), .A3(new_n444), .A4(new_n574), .ZN(new_n950));
  AOI21_X1  g749(.A(G169gat), .B1(new_n950), .B2(new_n248), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n949), .A2(new_n951), .ZN(G1348gat));
  OAI21_X1  g751(.A(G176gat), .B1(new_n948), .B2(new_n774), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n950), .A2(new_n363), .A3(new_n666), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1349gat));
  OAI21_X1  g754(.A(G183gat), .B1(new_n948), .B2(new_n647), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n950), .A2(new_n383), .A3(new_n385), .A4(new_n707), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT60), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n959), .A2(KEYINPUT125), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n958), .B(new_n960), .ZN(G1350gat));
  NAND3_X1  g760(.A1(new_n950), .A2(new_n386), .A3(new_n620), .ZN(new_n962));
  OR2_X1    g761(.A1(new_n948), .A2(new_n726), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT61), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n963), .A2(new_n964), .A3(G190gat), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n964), .B1(new_n963), .B2(G190gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n962), .B1(new_n965), .B2(new_n966), .ZN(G1351gat));
  NOR3_X1   g766(.A1(new_n671), .A2(new_n444), .A3(new_n694), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n922), .A2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(G197gat), .ZN(new_n970));
  NOR3_X1   g769(.A1(new_n969), .A2(new_n970), .A3(new_n249), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n860), .A2(new_n671), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n910), .A2(new_n444), .ZN(new_n973));
  AND2_X1   g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g773(.A(G197gat), .B1(new_n974), .B2(new_n248), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n971), .A2(new_n975), .ZN(G1352gat));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n774), .A2(G204gat), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n977), .B1(new_n974), .B2(new_n978), .ZN(new_n979));
  AND4_X1   g778(.A1(new_n977), .A2(new_n972), .A3(new_n973), .A4(new_n978), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT62), .ZN(new_n981));
  OR3_X1    g780(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  OAI21_X1  g781(.A(G204gat), .B1(new_n969), .B2(new_n774), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n981), .B1(new_n979), .B2(new_n980), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(G1353gat));
  INV_X1    g784(.A(G211gat), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n974), .A2(new_n986), .A3(new_n707), .ZN(new_n987));
  NAND4_X1  g786(.A1(new_n929), .A2(new_n968), .A3(new_n930), .A4(new_n707), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n988), .A2(G211gat), .ZN(new_n989));
  NOR2_X1   g788(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g790(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n989), .A2(new_n990), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n987), .B1(new_n993), .B2(new_n994), .ZN(G1354gat));
  OAI21_X1  g794(.A(G218gat), .B1(new_n969), .B2(new_n726), .ZN(new_n996));
  INV_X1    g795(.A(G218gat), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n974), .A2(new_n997), .A3(new_n620), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n996), .A2(new_n998), .ZN(G1355gat));
endmodule


