//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 1 1 1 1 1 1 1 1 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 1 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n613, new_n614, new_n615, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n790, new_n791, new_n793,
    new_n794, new_n795, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930;
  AND2_X1   g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  AND2_X1   g002(.A1(G211gat), .A2(G218gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(KEYINPUT22), .B2(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(G211gat), .B(G218gat), .Z(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G155gat), .B(G162gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n208), .B(KEYINPUT82), .ZN(new_n209));
  AND2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n211));
  OR2_X1    g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XOR2_X1   g011(.A(G141gat), .B(G148gat), .Z(new_n213));
  AOI21_X1  g012(.A(new_n209), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(KEYINPUT83), .B(G155gat), .Z(new_n215));
  AOI21_X1  g014(.A(new_n211), .B1(new_n215), .B2(G162gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(new_n208), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT29), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n207), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT3), .B1(new_n207), .B2(new_n222), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n202), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n223), .A2(new_n202), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT86), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n205), .A2(new_n228), .A3(new_n206), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n222), .B(new_n229), .C1(new_n207), .C2(new_n228), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n219), .B1(new_n230), .B2(new_n220), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n226), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  XOR2_X1   g031(.A(KEYINPUT31), .B(G50gat), .Z(new_n233));
  XNOR2_X1  g032(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G78gat), .B(G106gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n235), .B(G22gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n234), .B(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(G226gat), .A2(G233gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT25), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT24), .ZN(new_n241));
  INV_X1    g040(.A(G183gat), .ZN(new_n242));
  INV_X1    g041(.A(G190gat), .ZN(new_n243));
  NOR3_X1   g042(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(G183gat), .A2(G190gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT64), .ZN(new_n248));
  OR2_X1    g047(.A1(new_n247), .A2(KEYINPUT64), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n246), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n250), .B(KEYINPUT65), .Z(new_n251));
  INV_X1    g050(.A(G169gat), .ZN(new_n252));
  INV_X1    g051(.A(G176gat), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT23), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(G169gat), .A2(G176gat), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n255), .A2(KEYINPUT66), .A3(KEYINPUT23), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT66), .B1(new_n255), .B2(KEYINPUT23), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n260), .B(KEYINPUT67), .Z(new_n261));
  OAI21_X1  g060(.A(new_n240), .B1(new_n251), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n240), .B1(new_n255), .B2(KEYINPUT23), .ZN(new_n263));
  NAND2_X1  g062(.A1(G183gat), .A2(G190gat), .ZN(new_n264));
  AND2_X1   g063(.A1(KEYINPUT68), .A2(KEYINPUT24), .ZN(new_n265));
  NOR2_X1   g064(.A1(KEYINPUT68), .A2(KEYINPUT24), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(KEYINPUT69), .ZN(new_n268));
  INV_X1    g067(.A(new_n246), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n257), .B(new_n263), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT70), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n262), .A2(new_n271), .ZN(new_n272));
  AND2_X1   g071(.A1(KEYINPUT72), .A2(KEYINPUT26), .ZN(new_n273));
  NOR2_X1   g072(.A1(KEYINPUT72), .A2(KEYINPUT26), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n255), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n275), .B(KEYINPUT73), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n277), .B1(new_n256), .B2(KEYINPUT26), .ZN(new_n278));
  AND3_X1   g077(.A1(new_n256), .A2(new_n277), .A3(KEYINPUT26), .ZN(new_n279));
  OAI221_X1 g078(.A(new_n276), .B1(new_n252), .B2(new_n253), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT27), .B(G183gat), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n282), .A2(G190gat), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  OR2_X1    g083(.A1(new_n284), .A2(KEYINPUT28), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(KEYINPUT28), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n280), .A2(new_n264), .A3(new_n285), .A4(new_n286), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n272), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n239), .B1(new_n288), .B2(KEYINPUT29), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n287), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n290), .A2(G226gat), .A3(G233gat), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n207), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n289), .A2(new_n207), .A3(new_n291), .ZN(new_n294));
  XOR2_X1   g093(.A(G8gat), .B(G36gat), .Z(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(KEYINPUT79), .ZN(new_n296));
  XNOR2_X1  g095(.A(G64gat), .B(G92gat), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n296), .B(new_n297), .Z(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n293), .A2(KEYINPUT30), .A3(new_n294), .A4(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n294), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(new_n292), .ZN(new_n302));
  XOR2_X1   g101(.A(new_n298), .B(KEYINPUT80), .Z(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n300), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT30), .B1(new_n302), .B2(new_n299), .ZN(new_n306));
  OR2_X1    g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT3), .B1(new_n214), .B2(new_n218), .ZN(new_n308));
  XNOR2_X1  g107(.A(G113gat), .B(G120gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n309), .A2(KEYINPUT1), .ZN(new_n310));
  XNOR2_X1  g109(.A(G127gat), .B(G134gat), .ZN(new_n311));
  OR2_X1    g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n309), .A2(KEYINPUT74), .ZN(new_n313));
  INV_X1    g112(.A(G120gat), .ZN(new_n314));
  OR3_X1    g113(.A1(new_n314), .A2(KEYINPUT74), .A3(G113gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT75), .B(KEYINPUT1), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n313), .A2(new_n311), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n221), .A2(new_n308), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT4), .ZN(new_n320));
  INV_X1    g119(.A(new_n318), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n219), .A2(KEYINPUT84), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n219), .A2(new_n321), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n324), .B(new_n320), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT84), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n323), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G225gat), .A2(G233gat), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n329), .A2(KEYINPUT5), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT85), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT85), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n327), .A2(new_n333), .A3(new_n330), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n325), .A2(new_n329), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(new_n319), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT5), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n219), .B(new_n321), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n338), .B1(new_n339), .B2(new_n329), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n335), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G1gat), .B(G29gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n343), .B(KEYINPUT0), .ZN(new_n344));
  XNOR2_X1  g143(.A(G57gat), .B(G85gat), .ZN(new_n345));
  XOR2_X1   g144(.A(new_n344), .B(new_n345), .Z(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n327), .A2(new_n328), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT39), .B1(new_n339), .B2(new_n329), .ZN(new_n350));
  OR2_X1    g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT39), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n347), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n351), .A2(KEYINPUT40), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n348), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT40), .B1(new_n351), .B2(new_n353), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n307), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT37), .B1(new_n301), .B2(new_n292), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT37), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n293), .A2(new_n360), .A3(new_n294), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n359), .A2(new_n361), .A3(new_n298), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT87), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(new_n363), .A3(KEYINPUT38), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n363), .B1(new_n362), .B2(KEYINPUT38), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n332), .A2(new_n334), .B1(new_n337), .B2(new_n340), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT6), .B1(new_n368), .B2(new_n346), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n348), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n304), .A2(KEYINPUT38), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n359), .A2(new_n361), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n342), .A2(KEYINPUT6), .A3(new_n347), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n302), .A2(new_n299), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n370), .A2(new_n372), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n238), .B(new_n358), .C1(new_n367), .C2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n288), .A2(new_n318), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n290), .A2(new_n321), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n377), .A2(G227gat), .A3(G233gat), .A4(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT76), .B(KEYINPUT33), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G15gat), .B(G43gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(KEYINPUT77), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n383), .B(G71gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n384), .B(G99gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  XOR2_X1   g185(.A(KEYINPUT78), .B(KEYINPUT34), .Z(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n387), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n381), .A2(new_n389), .A3(new_n385), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n379), .A2(KEYINPUT32), .ZN(new_n392));
  NAND2_X1  g191(.A1(G227gat), .A2(G233gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n393), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n396), .A2(KEYINPUT32), .A3(new_n379), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n391), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n388), .A2(new_n395), .A3(new_n397), .A4(new_n390), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(KEYINPUT36), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n400), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT36), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n370), .A2(new_n373), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n305), .A2(KEYINPUT81), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT81), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n300), .B(new_n407), .C1(new_n302), .C2(new_n304), .ZN(new_n408));
  INV_X1    g207(.A(new_n306), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n405), .A2(new_n406), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  AOI22_X1  g209(.A1(new_n401), .A2(new_n404), .B1(new_n410), .B2(new_n237), .ZN(new_n411));
  AOI211_X1 g210(.A(KEYINPUT35), .B(new_n237), .C1(new_n373), .C2(new_n370), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n305), .A2(new_n306), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n399), .A2(KEYINPUT88), .A3(new_n400), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT88), .B1(new_n399), .B2(new_n400), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n412), .B(new_n413), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n238), .A3(new_n400), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT35), .B1(new_n410), .B2(new_n417), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n376), .A2(new_n411), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G229gat), .A2(G233gat), .ZN(new_n420));
  NOR2_X1   g219(.A1(G29gat), .A2(G36gat), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT14), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT89), .B(G29gat), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(G36gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(G43gat), .B(G50gat), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n423), .A2(new_n425), .A3(KEYINPUT15), .A4(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n423), .A2(new_n425), .A3(KEYINPUT15), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n426), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT15), .B1(new_n423), .B2(new_n425), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n428), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT17), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n423), .A2(new_n425), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT15), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n436), .A2(new_n429), .A3(new_n426), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT17), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(new_n438), .A3(new_n428), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n433), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G15gat), .B(G22gat), .ZN(new_n441));
  INV_X1    g240(.A(G1gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT16), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n444), .B1(G1gat), .B2(new_n441), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(G8gat), .ZN(new_n446));
  INV_X1    g245(.A(G8gat), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n444), .B(new_n447), .C1(G1gat), .C2(new_n441), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT90), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n449), .B(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n440), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n432), .A2(new_n449), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT91), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n454), .A2(KEYINPUT18), .ZN(new_n455));
  AND4_X1   g254(.A1(new_n420), .A2(new_n452), .A3(new_n453), .A4(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n453), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n457), .B1(new_n440), .B2(new_n451), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n455), .B1(new_n458), .B2(new_n420), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT92), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n460), .B1(new_n432), .B2(new_n449), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n446), .A2(new_n448), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n462), .A2(new_n437), .A3(KEYINPUT92), .A4(new_n428), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n461), .A2(new_n463), .A3(new_n453), .ZN(new_n464));
  XOR2_X1   g263(.A(new_n420), .B(KEYINPUT13), .Z(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n466), .A2(KEYINPUT93), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT93), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n468), .B1(new_n464), .B2(new_n465), .ZN(new_n469));
  OAI22_X1  g268(.A1(new_n456), .A2(new_n459), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(G113gat), .B(G141gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n471), .B(G197gat), .ZN(new_n472));
  XOR2_X1   g271(.A(KEYINPUT11), .B(G169gat), .Z(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(KEYINPUT12), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n466), .B(KEYINPUT93), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n452), .A2(new_n420), .A3(new_n453), .ZN(new_n479));
  INV_X1    g278(.A(new_n455), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n458), .A2(new_n420), .A3(new_n455), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n478), .A2(new_n483), .A3(new_n475), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n477), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n419), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(G231gat), .A2(G233gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(KEYINPUT99), .ZN(new_n489));
  XOR2_X1   g288(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n490));
  XOR2_X1   g289(.A(new_n489), .B(new_n490), .Z(new_n491));
  INV_X1    g290(.A(G57gat), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n492), .A2(G64gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT97), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(G64gat), .ZN(new_n495));
  INV_X1    g294(.A(G64gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(G57gat), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT97), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n494), .A2(new_n495), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT98), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT98), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n494), .A2(new_n499), .A3(new_n502), .A4(new_n495), .ZN(new_n503));
  INV_X1    g302(.A(G71gat), .ZN(new_n504));
  INV_X1    g303(.A(G78gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT9), .ZN(new_n506));
  NAND2_X1  g305(.A1(G71gat), .A2(G78gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n501), .A2(new_n503), .A3(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT95), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n496), .A2(G57gat), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n510), .B1(new_n511), .B2(new_n493), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n495), .A2(new_n497), .A3(KEYINPUT95), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT9), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n507), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n512), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT96), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n507), .A2(KEYINPUT94), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n507), .A2(KEYINPUT94), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n518), .A2(new_n519), .B1(new_n504), .B2(new_n505), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n516), .A2(new_n517), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n517), .B1(new_n516), .B2(new_n520), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n509), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT21), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(new_n462), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT100), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n526), .A2(KEYINPUT100), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n491), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n529), .ZN(new_n531));
  INV_X1    g330(.A(new_n491), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(new_n527), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(G127gat), .B(G155gat), .ZN(new_n535));
  NOR3_X1   g334(.A1(new_n524), .A2(KEYINPUT21), .A3(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(G183gat), .B(G211gat), .Z(new_n537));
  INV_X1    g336(.A(new_n535), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT21), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n538), .B1(new_n523), .B2(new_n539), .ZN(new_n540));
  OR3_X1    g339(.A1(new_n536), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n537), .B1(new_n536), .B2(new_n540), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n534), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n530), .A2(new_n533), .A3(new_n542), .A4(new_n541), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G190gat), .B(G218gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT102), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(G85gat), .A2(G92gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(G99gat), .A2(G106gat), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n550), .B1(KEYINPUT8), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G85gat), .A2(G92gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT7), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT7), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n555), .A2(G85gat), .A3(G92gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G99gat), .B(G106gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT101), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n440), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G232gat), .A2(G233gat), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT41), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n566), .B1(new_n432), .B2(new_n560), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n549), .B1(new_n563), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n563), .A2(new_n549), .A3(new_n567), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n564), .A2(new_n565), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(G134gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(G162gat), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n574), .B1(new_n568), .B2(KEYINPUT103), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n571), .B(new_n575), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n546), .A2(KEYINPUT104), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT104), .B1(new_n546), .B2(new_n576), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G230gat), .A2(G233gat), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n560), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n523), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT10), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n560), .B(new_n509), .C1(new_n521), .C2(new_n522), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n586), .A2(new_n585), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n582), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n581), .B1(new_n584), .B2(new_n586), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G120gat), .B(G148gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(G176gat), .B(G204gat), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n592), .B(new_n593), .Z(new_n594));
  XNOR2_X1  g393(.A(new_n591), .B(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n580), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n487), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n597), .A2(new_n405), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(new_n442), .ZN(G1324gat));
  INV_X1    g398(.A(new_n597), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n447), .B1(new_n600), .B2(new_n307), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT16), .B(G8gat), .ZN(new_n602));
  NOR3_X1   g401(.A1(new_n597), .A2(new_n413), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(KEYINPUT42), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n604), .B1(KEYINPUT42), .B2(new_n603), .ZN(G1325gat));
  NAND2_X1  g404(.A1(new_n404), .A2(new_n401), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT105), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(G15gat), .B1(new_n597), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n414), .A2(new_n415), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n610), .A2(G15gat), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n609), .B1(new_n597), .B2(new_n611), .ZN(G1326gat));
  NOR3_X1   g411(.A1(new_n419), .A2(new_n238), .A3(new_n486), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n596), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT43), .B(G22gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(G1327gat));
  INV_X1    g415(.A(KEYINPUT45), .ZN(new_n617));
  INV_X1    g416(.A(new_n546), .ZN(new_n618));
  INV_X1    g417(.A(new_n595), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n620), .A2(new_n576), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n487), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT106), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n405), .A2(new_n424), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n624), .B1(new_n623), .B2(new_n625), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n617), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n628), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n630), .A2(KEYINPUT45), .A3(new_n626), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT44), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n632), .B1(new_n419), .B2(new_n576), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n410), .A2(new_n237), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n358), .A2(new_n238), .ZN(new_n635));
  INV_X1    g434(.A(new_n366), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n375), .B1(new_n636), .B2(new_n364), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n606), .B(new_n634), .C1(new_n635), .C2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n416), .A2(new_n418), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n576), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n640), .A2(KEYINPUT44), .A3(new_n641), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n633), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n405), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n620), .A2(new_n486), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT107), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n424), .B1(new_n646), .B2(new_n647), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n629), .B(new_n631), .C1(new_n648), .C2(new_n649), .ZN(G1328gat));
  NOR3_X1   g449(.A1(new_n622), .A2(G36gat), .A3(new_n413), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT46), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n643), .A2(new_n645), .ZN(new_n653));
  OAI21_X1  g452(.A(G36gat), .B1(new_n653), .B2(new_n413), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(G1329gat));
  OAI21_X1  g454(.A(G43gat), .B1(new_n653), .B2(new_n606), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n622), .A2(G43gat), .A3(new_n610), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT47), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n633), .A2(new_n642), .A3(new_n607), .A4(new_n645), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n661), .A2(KEYINPUT108), .A3(G43gat), .ZN(new_n662));
  AOI21_X1  g461(.A(KEYINPUT108), .B1(new_n661), .B2(G43gat), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n662), .A2(new_n663), .A3(new_n657), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n660), .B1(new_n664), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g464(.A1(new_n633), .A2(new_n642), .A3(new_n237), .A4(new_n645), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(G50gat), .ZN(new_n667));
  INV_X1    g466(.A(G50gat), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n613), .A2(new_n668), .A3(new_n621), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n670), .B(KEYINPUT48), .Z(G1331gat));
  NOR3_X1   g470(.A1(new_n580), .A2(new_n485), .A3(new_n619), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n640), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n405), .B(KEYINPUT109), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(new_n492), .ZN(G1332gat));
  INV_X1    g475(.A(new_n673), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT110), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n413), .B(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT49), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n677), .B(new_n679), .C1(new_n680), .C2(new_n496), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT111), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n681), .A2(KEYINPUT111), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n681), .A2(KEYINPUT111), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n684), .A2(new_n680), .A3(new_n496), .A4(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n683), .A2(new_n686), .ZN(G1333gat));
  OAI21_X1  g486(.A(new_n504), .B1(new_n673), .B2(new_n610), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT112), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n608), .A2(new_n504), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n689), .B1(new_n690), .B2(new_n677), .ZN(new_n691));
  NOR4_X1   g490(.A1(new_n673), .A2(new_n608), .A3(KEYINPUT112), .A4(new_n504), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n688), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g493(.A1(new_n673), .A2(new_n238), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(new_n505), .ZN(G1335gat));
  NOR3_X1   g495(.A1(new_n546), .A2(new_n485), .A3(new_n619), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n643), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(G85gat), .B1(new_n698), .B2(new_n405), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT113), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n700), .B1(new_n419), .B2(new_n576), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n640), .A2(KEYINPUT113), .A3(new_n641), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n546), .A2(new_n485), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT51), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT51), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n701), .A2(new_n702), .A3(new_n706), .A4(new_n703), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n405), .A2(G85gat), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n705), .A2(new_n595), .A3(new_n707), .A4(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n699), .A2(new_n709), .ZN(G1336gat));
  NAND3_X1  g509(.A1(new_n643), .A2(new_n307), .A3(new_n697), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G92gat), .ZN(new_n712));
  INV_X1    g511(.A(new_n679), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(G92gat), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n705), .A2(new_n595), .A3(new_n707), .A4(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(KEYINPUT52), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n643), .A2(new_n679), .A3(new_n697), .ZN(new_n718));
  AOI21_X1  g517(.A(KEYINPUT52), .B1(new_n718), .B2(G92gat), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n715), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n717), .A2(new_n720), .ZN(G1337gat));
  OAI21_X1  g520(.A(G99gat), .B1(new_n698), .B2(new_n608), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n610), .A2(G99gat), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n705), .A2(new_n595), .A3(new_n707), .A4(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(G1338gat));
  NAND3_X1  g524(.A1(new_n643), .A2(new_n237), .A3(new_n697), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(G106gat), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n238), .A2(G106gat), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n705), .A2(new_n595), .A3(new_n707), .A4(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(KEYINPUT53), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT53), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n727), .A2(new_n729), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(G1339gat));
  NAND2_X1  g533(.A1(new_n546), .A2(new_n576), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n546), .A2(KEYINPUT104), .A3(new_n576), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n737), .A2(new_n486), .A3(new_n738), .A4(new_n619), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n587), .A2(new_n588), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n581), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT54), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n582), .B1(new_n586), .B2(new_n585), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n743), .B1(new_n745), .B2(new_n587), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n594), .B1(new_n589), .B2(new_n743), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT55), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n594), .ZN(new_n750));
  OR3_X1    g549(.A1(new_n589), .A2(new_n590), .A3(new_n750), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n752));
  OAI21_X1  g551(.A(KEYINPUT54), .B1(new_n752), .B2(new_n744), .ZN(new_n753));
  OAI21_X1  g552(.A(KEYINPUT55), .B1(new_n753), .B2(new_n589), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n741), .A2(new_n743), .A3(new_n581), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n750), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n751), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n747), .A2(new_n748), .A3(KEYINPUT55), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n760), .A2(KEYINPUT114), .A3(new_n751), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n749), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n458), .A2(new_n420), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n464), .A2(new_n465), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n474), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n484), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n576), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n762), .A2(new_n767), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n595), .A2(new_n484), .A3(new_n765), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n769), .B1(new_n762), .B2(new_n485), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n768), .B1(new_n770), .B2(new_n641), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n546), .B1(new_n771), .B2(KEYINPUT115), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n773), .B(new_n768), .C1(new_n770), .C2(new_n641), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n740), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n775), .A2(new_n674), .ZN(new_n776));
  INV_X1    g575(.A(new_n417), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(new_n679), .ZN(new_n779));
  AOI21_X1  g578(.A(G113gat), .B1(new_n779), .B2(new_n485), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n775), .A2(new_n237), .A3(new_n610), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n679), .A2(new_n405), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT116), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n783), .A2(KEYINPUT116), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n485), .A2(G113gat), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n780), .B1(new_n787), .B2(new_n788), .ZN(G1340gat));
  AOI21_X1  g588(.A(G120gat), .B1(new_n779), .B2(new_n595), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n619), .A2(new_n314), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n790), .B1(new_n787), .B2(new_n791), .ZN(G1341gat));
  INV_X1    g591(.A(G127gat), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n779), .A2(new_n793), .A3(new_n546), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n785), .A2(new_n786), .A3(new_n618), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n795), .B2(new_n793), .ZN(G1342gat));
  NAND2_X1  g595(.A1(new_n413), .A2(new_n641), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n778), .A2(G134gat), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT56), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n798), .B1(KEYINPUT117), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n799), .A2(KEYINPUT117), .ZN(new_n801));
  XOR2_X1   g600(.A(new_n800), .B(new_n801), .Z(new_n802));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n641), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(G134gat), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(G1343gat));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n806), .B(new_n807), .C1(new_n775), .C2(new_n238), .ZN(new_n808));
  INV_X1    g607(.A(new_n749), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n589), .A2(new_n590), .A3(new_n750), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n742), .B2(new_n746), .ZN(new_n812));
  AOI211_X1 g611(.A(new_n758), .B(new_n810), .C1(new_n748), .C2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT114), .B1(new_n760), .B2(new_n751), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n485), .B(new_n809), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n595), .A2(new_n484), .A3(new_n765), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n641), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n762), .A2(new_n767), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT115), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n819), .A2(new_n774), .A3(new_n618), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n238), .B1(new_n820), .B2(new_n739), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT118), .B1(new_n821), .B2(KEYINPUT57), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n238), .A2(new_n807), .ZN(new_n823));
  INV_X1    g622(.A(new_n757), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n485), .A2(new_n824), .A3(new_n809), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n825), .A2(new_n816), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n768), .B1(new_n826), .B2(new_n641), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n827), .A2(new_n618), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n823), .B1(new_n828), .B2(new_n740), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n808), .A2(new_n822), .A3(new_n829), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n782), .A2(new_n606), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(G141gat), .B1(new_n832), .B2(new_n486), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n607), .A2(new_n238), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(new_n713), .A3(new_n776), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n486), .A2(G141gat), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n833), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g637(.A(KEYINPUT122), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n782), .A2(new_n606), .A3(new_n595), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n579), .A2(KEYINPUT120), .A3(new_n486), .A4(new_n619), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n739), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n827), .A2(new_n618), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n238), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n845), .A2(KEYINPUT121), .A3(new_n846), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT57), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n820), .A2(new_n739), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n823), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n841), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n840), .B1(new_n855), .B2(G148gat), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n830), .A2(new_n595), .A3(new_n831), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n840), .A2(G148gat), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT119), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n857), .A2(new_n861), .A3(new_n858), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n856), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n835), .A2(G148gat), .A3(new_n619), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n839), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n864), .ZN(new_n866));
  AND3_X1   g665(.A1(new_n857), .A2(new_n861), .A3(new_n858), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n861), .B1(new_n857), .B2(new_n858), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI211_X1 g668(.A(KEYINPUT122), .B(new_n866), .C1(new_n869), .C2(new_n856), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n865), .A2(new_n870), .ZN(G1345gat));
  OAI21_X1  g670(.A(new_n215), .B1(new_n832), .B2(new_n618), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n618), .A2(new_n215), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n835), .B2(new_n873), .ZN(G1346gat));
  OAI21_X1  g673(.A(G162gat), .B1(new_n832), .B2(new_n576), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n797), .A2(G162gat), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n834), .A2(new_n776), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n877), .ZN(G1347gat));
  NAND2_X1  g677(.A1(new_n852), .A2(new_n405), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT123), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n679), .A2(new_n777), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(G169gat), .B1(new_n883), .B2(new_n485), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n674), .A2(new_n307), .ZN(new_n885));
  XOR2_X1   g684(.A(new_n885), .B(KEYINPUT124), .Z(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n781), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n887), .A2(new_n252), .A3(new_n486), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n884), .A2(new_n888), .ZN(G1348gat));
  NAND3_X1  g688(.A1(new_n883), .A2(new_n253), .A3(new_n595), .ZN(new_n890));
  OAI21_X1  g689(.A(G176gat), .B1(new_n887), .B2(new_n619), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(G1349gat));
  NAND4_X1  g691(.A1(new_n880), .A2(new_n281), .A3(new_n546), .A4(new_n882), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT125), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n893), .A2(new_n894), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n886), .A2(new_n546), .A3(new_n781), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  OAI22_X1  g697(.A1(new_n895), .A2(new_n896), .B1(new_n242), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT60), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT60), .ZN(new_n901));
  OAI221_X1 g700(.A(new_n901), .B1(new_n242), .B2(new_n898), .C1(new_n895), .C2(new_n896), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(G1350gat));
  NAND3_X1  g702(.A1(new_n883), .A2(new_n243), .A3(new_n641), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT126), .ZN(new_n905));
  OAI21_X1  g704(.A(G190gat), .B1(new_n887), .B2(new_n576), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT61), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(new_n907), .ZN(G1351gat));
  NOR3_X1   g707(.A1(new_n607), .A2(new_n238), .A3(new_n713), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n880), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(G197gat), .B1(new_n911), .B2(new_n485), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n849), .A2(new_n850), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n853), .B1(new_n913), .B2(KEYINPUT57), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n914), .A2(new_n608), .A3(new_n886), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n485), .A2(G197gat), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n912), .B1(new_n915), .B2(new_n916), .ZN(G1352gat));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n595), .ZN(new_n918));
  OR3_X1    g717(.A1(new_n910), .A2(G204gat), .A3(new_n619), .ZN(new_n919));
  AOI22_X1  g718(.A1(new_n918), .A2(G204gat), .B1(new_n919), .B2(KEYINPUT62), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n920), .B1(KEYINPUT62), .B2(new_n919), .ZN(G1353gat));
  OR3_X1    g720(.A1(new_n910), .A2(G211gat), .A3(new_n618), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n914), .A2(new_n546), .A3(new_n608), .A4(new_n886), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n923), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT63), .B1(new_n923), .B2(G211gat), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(G1354gat));
  AOI21_X1  g725(.A(G218gat), .B1(new_n911), .B2(new_n641), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n927), .A2(KEYINPUT127), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(KEYINPUT127), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n641), .A2(G218gat), .ZN(new_n930));
  AOI22_X1  g729(.A1(new_n928), .A2(new_n929), .B1(new_n915), .B2(new_n930), .ZN(G1355gat));
endmodule


